-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 23 2024 16:31:47

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    A : in std_logic_vector(31 downto 1);
    TICK50 : out std_logic;
    nROMEN : out std_logic;
    nCIACS1 : out std_logic;
    TICK60 : out std_logic;
    CLKCIA : out std_logic;
    CLK6 : in std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    TSn : in std_logic;
    nBUFEN : out std_logic;
    nREGSPACE : out std_logic;
    nRAMSPACE : out std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    TACKn : inout std_logic;
    nCIACS0 : out std_logic;
    PORTSIZE : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__6073\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2655\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2586\ : std_logic;
signal \N__2583\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2526\ : std_logic;
signal \N__2523\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2458\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2394\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2388\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2385\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2364\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U409_CIA.g0Z0Z_11\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U409_ADDRESS_DECODE.HIROM_0_cascade_\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U409_ADDRESS_DECODE.HIROM_0\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEm_6\ : std_logic;
signal \A_c_25\ : std_logic;
signal \U409_CIA.g0Z0Z_2_cascade_\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_28\ : std_logic;
signal \A_c_29\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\ : std_logic;
signal \A_c_24\ : std_logic;
signal \A_c_26\ : std_logic;
signal \A_c_31\ : std_logic;
signal \A_c_27\ : std_logic;
signal \U409_CIA.g0Z0Z_10\ : std_logic;
signal \A_c_22\ : std_logic;
signal \A_c_21\ : std_logic;
signal \U409_CIA.g0Z0Z_8\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_nREGSPACEZ0_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nREGSPACE_i\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.i6_mux_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.m9_bm_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_4\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.m9_am\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_97\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\ : std_logic;
signal \U409_ADDRESS_DECODE.HIROMZ0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_ROMEN_0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_ROMEN_0_cascade_\ : std_logic;
signal \ROMENm_i\ : std_logic;
signal \U409_TICK.TICK603_11_cascade_\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.TICK603_8\ : std_logic;
signal \bfn_10_6_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \bfn_10_7_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.RESETn_c_i\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\ : std_logic;
signal \TSn_c\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nCIACS1_i\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nCIACS0_i\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_CIA.N_9_cascade_\ : std_logic;
signal \U409_CIA.CIA_HOLDZ0\ : std_logic;
signal \U409_CIA.g0Z0Z_14\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \U409_CIA.g0Z0Z_13\ : std_logic;
signal \CIA_ENABLEm\ : std_logic;
signal \U409_CIA.N_20_cascade_\ : std_logic;
signal \U409_CIA.CLKCIA8_0_a2_0\ : std_logic;
signal \U409_CIA.CLKCIA6_0_a2_1\ : std_logic;
signal \U409_CIA.CLKCIAZ0_cascade_\ : std_logic;
signal \CLKCIA_c\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_EN_iC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\ : std_logic;
signal \U409_ADDRESS_DECODE_Z2_SPACE\ : std_logic;
signal \OVL_c\ : std_logic;
signal \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \bfn_12_7_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a2_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \TACK_EN_i\ : std_logic;
signal \N_353_i\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \nBUFEN_c\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \CLKCIA_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \nCIACS0_wire\ : std_logic;
signal \nCIACS1_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \nRAMSPACE_wire\ : std_logic;
signal \nROMEN_wire\ : std_logic;
signal \nBUFEN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \nREGSPACE_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    CLKCIA <= \CLKCIA_wire\;
    \A_wire\ <= A;
    nCIACS0 <= \nCIACS0_wire\;
    nCIACS1 <= \nCIACS1_wire\;
    \TSn_wire\ <= TSn;
    PORTSIZE <= \PORTSIZE_wire\;
    nRAMSPACE <= \nRAMSPACE_wire\;
    nROMEN <= \nROMEN_wire\;
    nBUFEN <= \nBUFEN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    nREGSPACE <= \nREGSPACE_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TICK60 <= \TICK60_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__3654\,
            RESETB => \N__4362\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6071\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6073\,
            DIN => \N__6072\,
            DOUT => \N__6071\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6073\,
            PADOUT => \N__6072\,
            PADIN => \N__6071\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6061\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6063\,
            DIN => \N__6062\,
            DOUT => \N__6061\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6063\,
            PADOUT => \N__6062\,
            PADIN => \N__6061\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKCIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6052\,
            DIN => \N__6051\,
            DOUT => \N__6050\,
            PACKAGEPIN => \CLKCIA_wire\
        );

    \CLKCIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6052\,
            PADOUT => \N__6051\,
            PADIN => \N__6050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4323\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6043\,
            DIN => \N__6042\,
            DOUT => \N__6041\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6043\,
            PADOUT => \N__6042\,
            PADIN => \N__6041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6034\,
            DIN => \N__6033\,
            DOUT => \N__6032\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6034\,
            PADOUT => \N__6033\,
            PADIN => \N__6032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCIACS0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6025\,
            DIN => \N__6024\,
            DOUT => \N__6023\,
            PACKAGEPIN => \nCIACS0_wire\
        );

    \nCIACS0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6025\,
            PADOUT => \N__6024\,
            PADIN => \N__6023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3720\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCIACS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6016\,
            DIN => \N__6015\,
            DOUT => \N__6014\,
            PACKAGEPIN => \nCIACS1_wire\
        );

    \nCIACS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6016\,
            PADOUT => \N__6015\,
            PADIN => \N__6014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3762\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6007\,
            DIN => \N__6006\,
            DOUT => \N__6005\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6007\,
            PADOUT => \N__6006\,
            PADIN => \N__6005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5998\,
            DIN => \N__5997\,
            DOUT => \N__5996\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5998\,
            PADOUT => \N__5997\,
            PADIN => \N__5996\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5989\,
            DIN => \N__5988\,
            DOUT => \N__5987\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5989\,
            PADOUT => \N__5988\,
            PADIN => \N__5987\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5980\,
            DIN => \N__5979\,
            DOUT => \N__5978\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__5980\,
            PADOUT => \N__5979\,
            PADIN => \N__5978\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5547\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__3846\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5971\,
            DIN => \N__5970\,
            DOUT => \N__5969\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5971\,
            PADOUT => \N__5970\,
            PADIN => \N__5969\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5962\,
            DIN => \N__5961\,
            DOUT => \N__5960\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5962\,
            PADOUT => \N__5961\,
            PADIN => \N__5960\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5953\,
            DIN => \N__5952\,
            DOUT => \N__5951\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5953\,
            PADOUT => \N__5952\,
            PADIN => \N__5951\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2973\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nRAMSPACE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5944\,
            DIN => \N__5943\,
            DOUT => \N__5942\,
            PACKAGEPIN => \nRAMSPACE_wire\
        );

    \nRAMSPACE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5944\,
            PADOUT => \N__5943\,
            PADIN => \N__5942\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4383\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nROMEN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5935\,
            DIN => \N__5934\,
            DOUT => \N__5933\,
            PACKAGEPIN => \nROMEN_wire\
        );

    \nROMEN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5935\,
            PADOUT => \N__5934\,
            PADIN => \N__5933\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3141\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5926\,
            DIN => \N__5925\,
            DOUT => \N__5924\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5926\,
            PADOUT => \N__5925\,
            PADIN => \N__5924\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5917\,
            DIN => \N__5916\,
            DOUT => \N__5915\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5917\,
            PADOUT => \N__5916\,
            PADIN => \N__5915\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nBUFEN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5908\,
            DIN => \N__5907\,
            DOUT => \N__5906\,
            PACKAGEPIN => \nBUFEN_wire\
        );

    \nBUFEN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5908\,
            PADOUT => \N__5907\,
            PADIN => \N__5906\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5511\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5899\,
            DIN => \N__5898\,
            DOUT => \N__5897\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5899\,
            PADOUT => \N__5898\,
            PADIN => \N__5897\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5890\,
            DIN => \N__5889\,
            DOUT => \N__5888\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5890\,
            PADOUT => \N__5889\,
            PADIN => \N__5888\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5881\,
            DIN => \N__5880\,
            DOUT => \N__5879\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5881\,
            PADOUT => \N__5880\,
            PADIN => \N__5879\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5872\,
            DIN => \N__5871\,
            DOUT => \N__5870\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5872\,
            PADOUT => \N__5871\,
            PADIN => \N__5870\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5863\,
            DIN => \N__5862\,
            DOUT => \N__5861\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5863\,
            PADOUT => \N__5862\,
            PADIN => \N__5861\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5854\,
            DIN => \N__5853\,
            DOUT => \N__5852\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5854\,
            PADOUT => \N__5853\,
            PADIN => \N__5852\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5845\,
            DIN => \N__5844\,
            DOUT => \N__5843\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5845\,
            PADOUT => \N__5844\,
            PADIN => \N__5843\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nREGSPACE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5836\,
            DIN => \N__5835\,
            DOUT => \N__5834\,
            PACKAGEPIN => \nREGSPACE_wire\
        );

    \nREGSPACE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5836\,
            PADOUT => \N__5835\,
            PADIN => \N__5834\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2871\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5827\,
            DIN => \N__5826\,
            DOUT => \N__5825\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5827\,
            PADOUT => \N__5826\,
            PADIN => \N__5825\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4233\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5818\,
            DIN => \N__5817\,
            DOUT => \N__5816\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5818\,
            PADOUT => \N__5817\,
            PADIN => \N__5816\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5809\,
            DIN => \N__5808\,
            DOUT => \N__5807\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5809\,
            PADOUT => \N__5808\,
            PADIN => \N__5807\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5800\,
            DIN => \N__5799\,
            DOUT => \N__5798\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5800\,
            PADOUT => \N__5799\,
            PADIN => \N__5798\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5791\,
            DIN => \N__5790\,
            DOUT => \N__5789\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5791\,
            PADOUT => \N__5790\,
            PADIN => \N__5789\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5782\,
            DIN => \N__5781\,
            DOUT => \N__5780\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5782\,
            PADOUT => \N__5781\,
            PADIN => \N__5780\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5773\,
            DIN => \N__5772\,
            DOUT => \N__5771\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5773\,
            PADOUT => \N__5772\,
            PADIN => \N__5771\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3282\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5764\,
            DIN => \N__5763\,
            DOUT => \N__5762\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5764\,
            PADOUT => \N__5763\,
            PADIN => \N__5762\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1332\ : CascadeMux
    port map (
            O => \N__5745\,
            I => \N__5742\
        );

    \I__1331\ : InMux
    port map (
            O => \N__5742\,
            I => \N__5736\
        );

    \I__1330\ : InMux
    port map (
            O => \N__5741\,
            I => \N__5731\
        );

    \I__1329\ : InMux
    port map (
            O => \N__5740\,
            I => \N__5731\
        );

    \I__1328\ : InMux
    port map (
            O => \N__5739\,
            I => \N__5728\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__5736\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__5731\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__5728\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1324\ : InMux
    port map (
            O => \N__5721\,
            I => \N__5713\
        );

    \I__1323\ : InMux
    port map (
            O => \N__5720\,
            I => \N__5713\
        );

    \I__1322\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5708\
        );

    \I__1321\ : InMux
    port map (
            O => \N__5718\,
            I => \N__5708\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__5713\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__5708\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__5703\,
            I => \N__5700\
        );

    \I__1317\ : InMux
    port map (
            O => \N__5700\,
            I => \N__5692\
        );

    \I__1316\ : InMux
    port map (
            O => \N__5699\,
            I => \N__5692\
        );

    \I__1315\ : InMux
    port map (
            O => \N__5698\,
            I => \N__5687\
        );

    \I__1314\ : InMux
    port map (
            O => \N__5697\,
            I => \N__5687\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5692\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__5687\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1311\ : InMux
    port map (
            O => \N__5682\,
            I => \N__5674\
        );

    \I__1310\ : InMux
    port map (
            O => \N__5681\,
            I => \N__5667\
        );

    \I__1309\ : InMux
    port map (
            O => \N__5680\,
            I => \N__5667\
        );

    \I__1308\ : InMux
    port map (
            O => \N__5679\,
            I => \N__5667\
        );

    \I__1307\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5662\
        );

    \I__1306\ : InMux
    port map (
            O => \N__5677\,
            I => \N__5662\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__5674\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__5667\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__5662\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5655\,
            I => \N__5652\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__5652\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\
        );

    \I__1300\ : CascadeMux
    port map (
            O => \N__5649\,
            I => \N__5639\
        );

    \I__1299\ : InMux
    port map (
            O => \N__5648\,
            I => \N__5636\
        );

    \I__1298\ : InMux
    port map (
            O => \N__5647\,
            I => \N__5627\
        );

    \I__1297\ : InMux
    port map (
            O => \N__5646\,
            I => \N__5627\
        );

    \I__1296\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5627\
        );

    \I__1295\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5627\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5620\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5642\,
            I => \N__5620\
        );

    \I__1292\ : InMux
    port map (
            O => \N__5639\,
            I => \N__5620\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5636\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__5627\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5620\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__5613\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_\
        );

    \I__1287\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5607\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__5607\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\
        );

    \I__1285\ : InMux
    port map (
            O => \N__5604\,
            I => \N__5593\
        );

    \I__1284\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5593\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5602\,
            I => \N__5588\
        );

    \I__1282\ : InMux
    port map (
            O => \N__5601\,
            I => \N__5588\
        );

    \I__1281\ : InMux
    port map (
            O => \N__5600\,
            I => \N__5581\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5599\,
            I => \N__5581\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5598\,
            I => \N__5581\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5593\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5588\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__5581\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1275\ : ClkMux
    port map (
            O => \N__5574\,
            I => \N__5565\
        );

    \I__1274\ : ClkMux
    port map (
            O => \N__5573\,
            I => \N__5565\
        );

    \I__1273\ : ClkMux
    port map (
            O => \N__5572\,
            I => \N__5565\
        );

    \I__1272\ : GlobalMux
    port map (
            O => \N__5565\,
            I => \N__5562\
        );

    \I__1271\ : gio2CtrlBuf
    port map (
            O => \N__5562\,
            I => \CLK28_IN_c_g\
        );

    \I__1270\ : InMux
    port map (
            O => \N__5559\,
            I => \N__5556\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__5556\,
            I => \N__5553\
        );

    \I__1268\ : Span4Mux_v
    port map (
            O => \N__5553\,
            I => \N__5550\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__5550\,
            I => \TACK_EN_i\
        );

    \I__1266\ : IoInMux
    port map (
            O => \N__5547\,
            I => \N__5544\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__5544\,
            I => \N__5541\
        );

    \I__1264\ : Span12Mux_s2_v
    port map (
            O => \N__5541\,
            I => \N__5538\
        );

    \I__1263\ : Span12Mux_v
    port map (
            O => \N__5538\,
            I => \N__5535\
        );

    \I__1262\ : Odrv12
    port map (
            O => \N__5535\,
            I => \N_353_i\
        );

    \I__1261\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5529\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__5529\,
            I => \N__5526\
        );

    \I__1259\ : Span4Mux_v
    port map (
            O => \N__5526\,
            I => \N__5523\
        );

    \I__1258\ : Sp12to4
    port map (
            O => \N__5523\,
            I => \N__5520\
        );

    \I__1257\ : Span12Mux_h
    port map (
            O => \N__5520\,
            I => \N__5517\
        );

    \I__1256\ : Span12Mux_v
    port map (
            O => \N__5517\,
            I => \N__5514\
        );

    \I__1255\ : Odrv12
    port map (
            O => \N__5514\,
            I => \TACKn_in\
        );

    \I__1254\ : IoInMux
    port map (
            O => \N__5511\,
            I => \N__5508\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__5508\,
            I => \N__5505\
        );

    \I__1252\ : Span12Mux_s9_v
    port map (
            O => \N__5505\,
            I => \N__5501\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5504\,
            I => \N__5498\
        );

    \I__1250\ : Span12Mux_h
    port map (
            O => \N__5501\,
            I => \N__5495\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5498\,
            I => \N__5492\
        );

    \I__1248\ : Odrv12
    port map (
            O => \N__5495\,
            I => \nBUFEN_c\
        );

    \I__1247\ : Odrv12
    port map (
            O => \N__5492\,
            I => \nBUFEN_c\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5482\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__5486\,
            I => \N__5476\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__5485\,
            I => \N__5463\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__5482\,
            I => \N__5459\
        );

    \I__1242\ : InMux
    port map (
            O => \N__5481\,
            I => \N__5448\
        );

    \I__1241\ : InMux
    port map (
            O => \N__5480\,
            I => \N__5448\
        );

    \I__1240\ : InMux
    port map (
            O => \N__5479\,
            I => \N__5448\
        );

    \I__1239\ : InMux
    port map (
            O => \N__5476\,
            I => \N__5448\
        );

    \I__1238\ : InMux
    port map (
            O => \N__5475\,
            I => \N__5448\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5474\,
            I => \N__5439\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5473\,
            I => \N__5439\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5472\,
            I => \N__5439\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5471\,
            I => \N__5439\
        );

    \I__1233\ : InMux
    port map (
            O => \N__5470\,
            I => \N__5436\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5469\,
            I => \N__5433\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5430\
        );

    \I__1230\ : InMux
    port map (
            O => \N__5467\,
            I => \N__5420\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5466\,
            I => \N__5420\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5463\,
            I => \N__5420\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5462\,
            I => \N__5420\
        );

    \I__1226\ : Span4Mux_v
    port map (
            O => \N__5459\,
            I => \N__5411\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__5448\,
            I => \N__5411\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5439\,
            I => \N__5411\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5436\,
            I => \N__5411\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__5433\,
            I => \N__5407\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5430\,
            I => \N__5404\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5429\,
            I => \N__5400\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5420\,
            I => \N__5395\
        );

    \I__1218\ : Span4Mux_v
    port map (
            O => \N__5411\,
            I => \N__5395\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5410\,
            I => \N__5392\
        );

    \I__1216\ : Span4Mux_v
    port map (
            O => \N__5407\,
            I => \N__5389\
        );

    \I__1215\ : Span4Mux_v
    port map (
            O => \N__5404\,
            I => \N__5386\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5383\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5400\,
            I => \N__5380\
        );

    \I__1212\ : Span4Mux_h
    port map (
            O => \N__5395\,
            I => \N__5377\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5392\,
            I => \N__5374\
        );

    \I__1210\ : Sp12to4
    port map (
            O => \N__5389\,
            I => \N__5371\
        );

    \I__1209\ : Span4Mux_h
    port map (
            O => \N__5386\,
            I => \N__5366\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__5383\,
            I => \N__5366\
        );

    \I__1207\ : Span4Mux_h
    port map (
            O => \N__5380\,
            I => \N__5363\
        );

    \I__1206\ : Span4Mux_h
    port map (
            O => \N__5377\,
            I => \N__5358\
        );

    \I__1205\ : Span4Mux_v
    port map (
            O => \N__5374\,
            I => \N__5358\
        );

    \I__1204\ : Span12Mux_h
    port map (
            O => \N__5371\,
            I => \N__5351\
        );

    \I__1203\ : Sp12to4
    port map (
            O => \N__5366\,
            I => \N__5351\
        );

    \I__1202\ : Sp12to4
    port map (
            O => \N__5363\,
            I => \N__5351\
        );

    \I__1201\ : Sp12to4
    port map (
            O => \N__5358\,
            I => \N__5348\
        );

    \I__1200\ : Span12Mux_v
    port map (
            O => \N__5351\,
            I => \N__5345\
        );

    \I__1199\ : Span12Mux_h
    port map (
            O => \N__5348\,
            I => \N__5342\
        );

    \I__1198\ : Span12Mux_h
    port map (
            O => \N__5345\,
            I => \N__5337\
        );

    \I__1197\ : Span12Mux_v
    port map (
            O => \N__5342\,
            I => \N__5337\
        );

    \I__1196\ : Odrv12
    port map (
            O => \N__5337\,
            I => \RESETn_c\
        );

    \I__1195\ : SRMux
    port map (
            O => \N__5334\,
            I => \N__5331\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5331\,
            I => \N__5328\
        );

    \I__1193\ : Span4Mux_v
    port map (
            O => \N__5328\,
            I => \N__5323\
        );

    \I__1192\ : SRMux
    port map (
            O => \N__5327\,
            I => \N__5320\
        );

    \I__1191\ : SRMux
    port map (
            O => \N__5326\,
            I => \N__5317\
        );

    \I__1190\ : Span4Mux_v
    port map (
            O => \N__5323\,
            I => \N__5310\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5320\,
            I => \N__5310\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__5317\,
            I => \N__5310\
        );

    \I__1187\ : Span4Mux_v
    port map (
            O => \N__5310\,
            I => \N__5307\
        );

    \I__1186\ : Span4Mux_h
    port map (
            O => \N__5307\,
            I => \N__5304\
        );

    \I__1185\ : Odrv4
    port map (
            O => \N__5304\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5301\,
            I => \N__5298\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5298\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5295\,
            I => \N__5292\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5292\,
            I => \N__5289\
        );

    \I__1180\ : Span4Mux_h
    port map (
            O => \N__5289\,
            I => \N__5285\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5288\,
            I => \N__5282\
        );

    \I__1178\ : Odrv4
    port map (
            O => \N__5285\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__5282\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5277\,
            I => \N__5262\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5262\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5262\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5255\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5255\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5255\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5271\,
            I => \N__5248\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5270\,
            I => \N__5248\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5248\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__5262\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5255\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5248\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5238\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__5235\,
            I => \N__5232\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5224\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__5231\,
            I => \N__5220\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__5230\,
            I => \N__5217\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__5229\,
            I => \N__5214\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__5228\,
            I => \N__5211\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__5227\,
            I => \N__5208\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__5224\,
            I => \N__5204\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5223\,
            I => \N__5197\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5197\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5217\,
            I => \N__5197\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5192\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5192\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5187\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5187\
        );

    \I__1147\ : Odrv4
    port map (
            O => \N__5204\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5197\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5192\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__5187\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5178\,
            I => \N__5166\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5177\,
            I => \N__5166\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5159\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5175\,
            I => \N__5159\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5174\,
            I => \N__5159\
        );

    \I__1138\ : InMux
    port map (
            O => \N__5173\,
            I => \N__5152\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5172\,
            I => \N__5152\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5171\,
            I => \N__5152\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5166\,
            I => \N__5149\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__5159\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__5152\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1132\ : Odrv4
    port map (
            O => \N__5149\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5142\,
            I => \N__5138\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5141\,
            I => \N__5135\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__5138\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5135\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__1127\ : ClkMux
    port map (
            O => \N__5130\,
            I => \N__5100\
        );

    \I__1126\ : ClkMux
    port map (
            O => \N__5129\,
            I => \N__5100\
        );

    \I__1125\ : ClkMux
    port map (
            O => \N__5128\,
            I => \N__5100\
        );

    \I__1124\ : ClkMux
    port map (
            O => \N__5127\,
            I => \N__5100\
        );

    \I__1123\ : ClkMux
    port map (
            O => \N__5126\,
            I => \N__5100\
        );

    \I__1122\ : ClkMux
    port map (
            O => \N__5125\,
            I => \N__5100\
        );

    \I__1121\ : ClkMux
    port map (
            O => \N__5124\,
            I => \N__5100\
        );

    \I__1120\ : ClkMux
    port map (
            O => \N__5123\,
            I => \N__5100\
        );

    \I__1119\ : ClkMux
    port map (
            O => \N__5122\,
            I => \N__5100\
        );

    \I__1118\ : ClkMux
    port map (
            O => \N__5121\,
            I => \N__5100\
        );

    \I__1117\ : GlobalMux
    port map (
            O => \N__5100\,
            I => \N__5097\
        );

    \I__1116\ : gio2CtrlBuf
    port map (
            O => \N__5097\,
            I => \CLK6_c_g\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5094\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5091\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5088\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__1112\ : InMux
    port map (
            O => \N__5085\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__5082\,
            I => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5079\,
            I => \bfn_12_7_0_\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5072\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5075\,
            I => \N__5069\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__5072\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__5069\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5064\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__5061\,
            I => \N__5058\
        );

    \I__1103\ : InMux
    port map (
            O => \N__5058\,
            I => \N__5054\
        );

    \I__1102\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5051\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5054\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5051\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__1099\ : InMux
    port map (
            O => \N__5046\,
            I => \N__5043\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5043\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5040\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5033\
        );

    \I__1095\ : InMux
    port map (
            O => \N__5036\,
            I => \N__5030\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__5033\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5030\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__1092\ : InMux
    port map (
            O => \N__5025\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5022\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5019\,
            I => \N__5015\
        );

    \I__1089\ : InMux
    port map (
            O => \N__5018\,
            I => \N__5012\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5015\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__5012\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5007\,
            I => \N__5004\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5004\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5001\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__1083\ : InMux
    port map (
            O => \N__4998\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__1082\ : InMux
    port map (
            O => \N__4995\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__1081\ : CascadeMux
    port map (
            O => \N__4992\,
            I => \N__4988\
        );

    \I__1080\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4985\
        );

    \I__1079\ : InMux
    port map (
            O => \N__4988\,
            I => \N__4982\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__4985\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__4982\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__4977\,
            I => \N__4974\
        );

    \I__1075\ : InMux
    port map (
            O => \N__4974\,
            I => \N__4971\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__4971\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__1073\ : InMux
    port map (
            O => \N__4968\,
            I => \N__4964\
        );

    \I__1072\ : InMux
    port map (
            O => \N__4967\,
            I => \N__4961\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__4964\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__4961\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1069\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4950\
        );

    \I__1068\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4950\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__4950\,
            I => \N__4946\
        );

    \I__1066\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4943\
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__4946\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__4943\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1063\ : CascadeMux
    port map (
            O => \N__4938\,
            I => \N__4932\
        );

    \I__1062\ : InMux
    port map (
            O => \N__4937\,
            I => \N__4927\
        );

    \I__1061\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4927\
        );

    \I__1060\ : InMux
    port map (
            O => \N__4935\,
            I => \N__4924\
        );

    \I__1059\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4921\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__4927\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__4924\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__4921\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1055\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4911\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__4911\,
            I => \N__4907\
        );

    \I__1053\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4904\
        );

    \I__1052\ : Odrv4
    port map (
            O => \N__4907\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__4904\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__1050\ : InMux
    port map (
            O => \N__4899\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__1049\ : InMux
    port map (
            O => \N__4896\,
            I => \N__4892\
        );

    \I__1048\ : InMux
    port map (
            O => \N__4895\,
            I => \N__4889\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__4892\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__4889\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__1045\ : InMux
    port map (
            O => \N__4884\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__1044\ : InMux
    port map (
            O => \N__4881\,
            I => \N__4877\
        );

    \I__1043\ : InMux
    port map (
            O => \N__4880\,
            I => \N__4874\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__4877\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__4874\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4869\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4862\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4859\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__4862\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4859\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__1035\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4851\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__4851\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__1033\ : InMux
    port map (
            O => \N__4848\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__4845\,
            I => \N__4841\
        );

    \I__1031\ : InMux
    port map (
            O => \N__4844\,
            I => \N__4838\
        );

    \I__1030\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4835\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__4838\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__4835\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__1027\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4827\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__4827\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4824\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__4821\,
            I => \N__4818\
        );

    \I__1023\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4814\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4817\,
            I => \N__4811\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__4814\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__4811\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4806\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__1018\ : InMux
    port map (
            O => \N__4803\,
            I => \N__4799\
        );

    \I__1017\ : InMux
    port map (
            O => \N__4802\,
            I => \N__4796\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__4799\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__4796\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4791\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__4788\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4785\,
            I => \N__4781\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4778\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4781\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__4778\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4773\,
            I => \N__4764\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4772\,
            I => \N__4764\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4771\,
            I => \N__4761\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4770\,
            I => \N__4758\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4769\,
            I => \N__4755\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__4764\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__4761\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__4758\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4755\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__999\ : InMux
    port map (
            O => \N__4746\,
            I => \N__4740\
        );

    \I__998\ : InMux
    port map (
            O => \N__4745\,
            I => \N__4737\
        );

    \I__997\ : InMux
    port map (
            O => \N__4744\,
            I => \N__4732\
        );

    \I__996\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4732\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__4740\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4737\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4732\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__992\ : InMux
    port map (
            O => \N__4725\,
            I => \N__4721\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__4724\,
            I => \N__4716\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__4721\,
            I => \N__4713\
        );

    \I__989\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4710\
        );

    \I__988\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4705\
        );

    \I__987\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4705\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__4713\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__4710\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__4705\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__983\ : InMux
    port map (
            O => \N__4698\,
            I => \N__4693\
        );

    \I__982\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4688\
        );

    \I__981\ : InMux
    port map (
            O => \N__4696\,
            I => \N__4688\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4693\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4688\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__978\ : InMux
    port map (
            O => \N__4683\,
            I => \N__4677\
        );

    \I__977\ : InMux
    port map (
            O => \N__4682\,
            I => \N__4674\
        );

    \I__976\ : InMux
    port map (
            O => \N__4681\,
            I => \N__4671\
        );

    \I__975\ : InMux
    port map (
            O => \N__4680\,
            I => \N__4668\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__4677\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4674\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4671\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4668\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__4659\,
            I => \N__4650\
        );

    \I__969\ : InMux
    port map (
            O => \N__4658\,
            I => \N__4645\
        );

    \I__968\ : InMux
    port map (
            O => \N__4657\,
            I => \N__4645\
        );

    \I__967\ : InMux
    port map (
            O => \N__4656\,
            I => \N__4642\
        );

    \I__966\ : InMux
    port map (
            O => \N__4655\,
            I => \N__4633\
        );

    \I__965\ : InMux
    port map (
            O => \N__4654\,
            I => \N__4633\
        );

    \I__964\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4633\
        );

    \I__963\ : InMux
    port map (
            O => \N__4650\,
            I => \N__4633\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__4645\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4642\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4633\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__4626\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\
        );

    \I__958\ : InMux
    port map (
            O => \N__4623\,
            I => \N__4616\
        );

    \I__957\ : InMux
    port map (
            O => \N__4622\,
            I => \N__4616\
        );

    \I__956\ : InMux
    port map (
            O => \N__4621\,
            I => \N__4613\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4616\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4613\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__953\ : InMux
    port map (
            O => \N__4608\,
            I => \N__4601\
        );

    \I__952\ : InMux
    port map (
            O => \N__4607\,
            I => \N__4598\
        );

    \I__951\ : InMux
    port map (
            O => \N__4606\,
            I => \N__4591\
        );

    \I__950\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4591\
        );

    \I__949\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4591\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4601\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4598\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4591\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__945\ : CascadeMux
    port map (
            O => \N__4584\,
            I => \N__4579\
        );

    \I__944\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4575\
        );

    \I__943\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4572\
        );

    \I__942\ : InMux
    port map (
            O => \N__4579\,
            I => \N__4567\
        );

    \I__941\ : InMux
    port map (
            O => \N__4578\,
            I => \N__4567\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4575\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4572\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4567\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__937\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4554\
        );

    \I__936\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4554\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4554\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__934\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4547\
        );

    \I__933\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4544\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4547\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4544\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\
        );

    \I__930\ : CEMux
    port map (
            O => \N__4539\,
            I => \N__4536\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4536\,
            I => \N__4533\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__4533\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__4530\,
            I => \N__4527\
        );

    \I__926\ : InMux
    port map (
            O => \N__4527\,
            I => \N__4520\
        );

    \I__925\ : InMux
    port map (
            O => \N__4526\,
            I => \N__4517\
        );

    \I__924\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4513\
        );

    \I__923\ : InMux
    port map (
            O => \N__4524\,
            I => \N__4510\
        );

    \I__922\ : InMux
    port map (
            O => \N__4523\,
            I => \N__4507\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4520\,
            I => \N__4502\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4517\,
            I => \N__4502\
        );

    \I__919\ : InMux
    port map (
            O => \N__4516\,
            I => \N__4499\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4513\,
            I => \N__4496\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4510\,
            I => \N__4493\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4507\,
            I => \N__4490\
        );

    \I__915\ : Span4Mux_v
    port map (
            O => \N__4502\,
            I => \N__4485\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4499\,
            I => \N__4485\
        );

    \I__913\ : Span4Mux_v
    port map (
            O => \N__4496\,
            I => \N__4482\
        );

    \I__912\ : Span4Mux_v
    port map (
            O => \N__4493\,
            I => \N__4479\
        );

    \I__911\ : Span4Mux_v
    port map (
            O => \N__4490\,
            I => \N__4476\
        );

    \I__910\ : Span4Mux_h
    port map (
            O => \N__4485\,
            I => \N__4472\
        );

    \I__909\ : Sp12to4
    port map (
            O => \N__4482\,
            I => \N__4465\
        );

    \I__908\ : Sp12to4
    port map (
            O => \N__4479\,
            I => \N__4465\
        );

    \I__907\ : Sp12to4
    port map (
            O => \N__4476\,
            I => \N__4465\
        );

    \I__906\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4462\
        );

    \I__905\ : Span4Mux_v
    port map (
            O => \N__4472\,
            I => \N__4459\
        );

    \I__904\ : Span12Mux_h
    port map (
            O => \N__4465\,
            I => \N__4454\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4462\,
            I => \N__4454\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__4459\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__901\ : Odrv12
    port map (
            O => \N__4454\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__900\ : InMux
    port map (
            O => \N__4449\,
            I => \N__4444\
        );

    \I__899\ : InMux
    port map (
            O => \N__4448\,
            I => \N__4441\
        );

    \I__898\ : InMux
    port map (
            O => \N__4447\,
            I => \N__4438\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4444\,
            I => \N__4435\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4441\,
            I => \N__4430\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4438\,
            I => \N__4430\
        );

    \I__894\ : Span4Mux_v
    port map (
            O => \N__4435\,
            I => \N__4427\
        );

    \I__893\ : Span4Mux_v
    port map (
            O => \N__4430\,
            I => \N__4424\
        );

    \I__892\ : Sp12to4
    port map (
            O => \N__4427\,
            I => \N__4419\
        );

    \I__891\ : Sp12to4
    port map (
            O => \N__4424\,
            I => \N__4419\
        );

    \I__890\ : Span12Mux_h
    port map (
            O => \N__4419\,
            I => \N__4416\
        );

    \I__889\ : Span12Mux_v
    port map (
            O => \N__4416\,
            I => \N__4413\
        );

    \I__888\ : Odrv12
    port map (
            O => \N__4413\,
            I => \OVL_c\
        );

    \I__887\ : InMux
    port map (
            O => \N__4410\,
            I => \N__4406\
        );

    \I__886\ : InMux
    port map (
            O => \N__4409\,
            I => \N__4403\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4406\,
            I => \N__4399\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4403\,
            I => \N__4396\
        );

    \I__883\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4393\
        );

    \I__882\ : Span12Mux_h
    port map (
            O => \N__4399\,
            I => \N__4386\
        );

    \I__881\ : Sp12to4
    port map (
            O => \N__4396\,
            I => \N__4386\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4393\,
            I => \N__4386\
        );

    \I__879\ : Odrv12
    port map (
            O => \N__4386\,
            I => \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0\
        );

    \I__878\ : IoInMux
    port map (
            O => \N__4383\,
            I => \N__4380\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__4380\,
            I => \N__4377\
        );

    \I__876\ : Span4Mux_s3_v
    port map (
            O => \N__4377\,
            I => \N__4374\
        );

    \I__875\ : Span4Mux_v
    port map (
            O => \N__4374\,
            I => \N__4371\
        );

    \I__874\ : Span4Mux_v
    port map (
            O => \N__4371\,
            I => \N__4368\
        );

    \I__873\ : Span4Mux_v
    port map (
            O => \N__4368\,
            I => \N__4365\
        );

    \I__872\ : Odrv4
    port map (
            O => \N__4365\,
            I => \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\
        );

    \I__871\ : IoInMux
    port map (
            O => \N__4362\,
            I => \N__4359\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4359\,
            I => \N__4356\
        );

    \I__869\ : Span4Mux_s3_v
    port map (
            O => \N__4356\,
            I => \N__4353\
        );

    \I__868\ : Span4Mux_h
    port map (
            O => \N__4353\,
            I => \N__4350\
        );

    \I__867\ : Odrv4
    port map (
            O => \N__4350\,
            I => \CONSTANT_ONE_NET\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__4347\,
            I => \U409_CIA.N_20_cascade_\
        );

    \I__865\ : InMux
    port map (
            O => \N__4344\,
            I => \N__4340\
        );

    \I__864\ : InMux
    port map (
            O => \N__4343\,
            I => \N__4337\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__4340\,
            I => \U409_CIA.CLKCIA8_0_a2_0\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4337\,
            I => \U409_CIA.CLKCIA8_0_a2_0\
        );

    \I__861\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4329\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4329\,
            I => \U409_CIA.CLKCIA6_0_a2_1\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__4326\,
            I => \U409_CIA.CLKCIAZ0_cascade_\
        );

    \I__858\ : IoInMux
    port map (
            O => \N__4323\,
            I => \N__4320\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4320\,
            I => \N__4317\
        );

    \I__856\ : Span4Mux_s1_v
    port map (
            O => \N__4317\,
            I => \N__4314\
        );

    \I__855\ : Span4Mux_v
    port map (
            O => \N__4314\,
            I => \N__4311\
        );

    \I__854\ : Sp12to4
    port map (
            O => \N__4311\,
            I => \N__4308\
        );

    \I__853\ : Span12Mux_h
    port map (
            O => \N__4308\,
            I => \N__4304\
        );

    \I__852\ : InMux
    port map (
            O => \N__4307\,
            I => \N__4301\
        );

    \I__851\ : Span12Mux_v
    port map (
            O => \N__4304\,
            I => \N__4295\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4301\,
            I => \N__4295\
        );

    \I__849\ : InMux
    port map (
            O => \N__4300\,
            I => \N__4292\
        );

    \I__848\ : Odrv12
    port map (
            O => \N__4295\,
            I => \CLKCIA_c\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4292\,
            I => \CLKCIA_c\
        );

    \I__846\ : InMux
    port map (
            O => \N__4287\,
            I => \N__4284\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4284\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__4281\,
            I => \N__4278\
        );

    \I__843\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4271\
        );

    \I__842\ : InMux
    port map (
            O => \N__4277\,
            I => \N__4271\
        );

    \I__841\ : InMux
    port map (
            O => \N__4276\,
            I => \N__4268\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4271\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4268\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__4263\,
            I => \N__4259\
        );

    \I__837\ : InMux
    port map (
            O => \N__4262\,
            I => \N__4253\
        );

    \I__836\ : InMux
    port map (
            O => \N__4259\,
            I => \N__4246\
        );

    \I__835\ : InMux
    port map (
            O => \N__4258\,
            I => \N__4246\
        );

    \I__834\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4246\
        );

    \I__833\ : InMux
    port map (
            O => \N__4256\,
            I => \N__4243\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4253\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4246\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__4243\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__4236\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__828\ : IoInMux
    port map (
            O => \N__4233\,
            I => \N__4230\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4230\,
            I => \N__4227\
        );

    \I__826\ : Span4Mux_s3_v
    port map (
            O => \N__4227\,
            I => \N__4224\
        );

    \I__825\ : Span4Mux_h
    port map (
            O => \N__4224\,
            I => \N__4221\
        );

    \I__824\ : Sp12to4
    port map (
            O => \N__4221\,
            I => \N__4218\
        );

    \I__823\ : Span12Mux_v
    port map (
            O => \N__4218\,
            I => \N__4214\
        );

    \I__822\ : InMux
    port map (
            O => \N__4217\,
            I => \N__4211\
        );

    \I__821\ : Odrv12
    port map (
            O => \N__4214\,
            I => \TICK50_c\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4211\,
            I => \TICK50_c\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__4206\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__4203\,
            I => \U409_CIA.N_9_cascade_\
        );

    \I__817\ : InMux
    port map (
            O => \N__4200\,
            I => \N__4195\
        );

    \I__816\ : InMux
    port map (
            O => \N__4199\,
            I => \N__4190\
        );

    \I__815\ : InMux
    port map (
            O => \N__4198\,
            I => \N__4190\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4195\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__4190\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__812\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4178\
        );

    \I__811\ : InMux
    port map (
            O => \N__4184\,
            I => \N__4178\
        );

    \I__810\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4175\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4178\,
            I => \N__4170\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4175\,
            I => \N__4170\
        );

    \I__807\ : Odrv12
    port map (
            O => \N__4170\,
            I => \U409_CIA.g0Z0Z_14\
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__4167\,
            I => \N__4163\
        );

    \I__805\ : InMux
    port map (
            O => \N__4166\,
            I => \N__4158\
        );

    \I__804\ : InMux
    port map (
            O => \N__4163\,
            I => \N__4151\
        );

    \I__803\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4151\
        );

    \I__802\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4151\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4158\,
            I => \U409_CIA.VMAZ0\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4151\,
            I => \U409_CIA.VMAZ0\
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__4146\,
            I => \N__4142\
        );

    \I__798\ : InMux
    port map (
            O => \N__4145\,
            I => \N__4136\
        );

    \I__797\ : InMux
    port map (
            O => \N__4142\,
            I => \N__4136\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__4141\,
            I => \N__4133\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__4136\,
            I => \N__4130\
        );

    \I__794\ : InMux
    port map (
            O => \N__4133\,
            I => \N__4127\
        );

    \I__793\ : Span4Mux_v
    port map (
            O => \N__4130\,
            I => \N__4124\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4127\,
            I => \N__4121\
        );

    \I__791\ : Span4Mux_h
    port map (
            O => \N__4124\,
            I => \N__4118\
        );

    \I__790\ : Span4Mux_v
    port map (
            O => \N__4121\,
            I => \N__4115\
        );

    \I__789\ : Sp12to4
    port map (
            O => \N__4118\,
            I => \N__4110\
        );

    \I__788\ : Sp12to4
    port map (
            O => \N__4115\,
            I => \N__4110\
        );

    \I__787\ : Span12Mux_h
    port map (
            O => \N__4110\,
            I => \N__4107\
        );

    \I__786\ : Odrv12
    port map (
            O => \N__4107\,
            I => \U409_CIA.g0Z0Z_13\
        );

    \I__785\ : InMux
    port map (
            O => \N__4104\,
            I => \N__4098\
        );

    \I__784\ : InMux
    port map (
            O => \N__4103\,
            I => \N__4098\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4098\,
            I => \N__4095\
        );

    \I__782\ : Odrv12
    port map (
            O => \N__4095\,
            I => \CIA_ENABLEm\
        );

    \I__781\ : CascadeMux
    port map (
            O => \N__4092\,
            I => \N__4088\
        );

    \I__780\ : InMux
    port map (
            O => \N__4091\,
            I => \N__4083\
        );

    \I__779\ : InMux
    port map (
            O => \N__4088\,
            I => \N__4080\
        );

    \I__778\ : InMux
    port map (
            O => \N__4087\,
            I => \N__4077\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__4086\,
            I => \N__4074\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4083\,
            I => \N__4071\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4080\,
            I => \N__4066\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4077\,
            I => \N__4066\
        );

    \I__773\ : InMux
    port map (
            O => \N__4074\,
            I => \N__4063\
        );

    \I__772\ : Odrv4
    port map (
            O => \N__4071\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__4066\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4063\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__4056\,
            I => \N__4052\
        );

    \I__768\ : InMux
    port map (
            O => \N__4055\,
            I => \N__4048\
        );

    \I__767\ : InMux
    port map (
            O => \N__4052\,
            I => \N__4045\
        );

    \I__766\ : InMux
    port map (
            O => \N__4051\,
            I => \N__4042\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4048\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4045\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__4042\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__762\ : InMux
    port map (
            O => \N__4035\,
            I => \N__4031\
        );

    \I__761\ : InMux
    port map (
            O => \N__4034\,
            I => \N__4028\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4031\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4028\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__4023\,
            I => \N__4020\
        );

    \I__757\ : InMux
    port map (
            O => \N__4020\,
            I => \N__4016\
        );

    \I__756\ : InMux
    port map (
            O => \N__4019\,
            I => \N__4013\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4016\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__4013\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__753\ : InMux
    port map (
            O => \N__4008\,
            I => \N__4004\
        );

    \I__752\ : InMux
    port map (
            O => \N__4007\,
            I => \N__4001\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4004\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__4001\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__3996\,
            I => \N__3991\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__3995\,
            I => \N__3988\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__3994\,
            I => \N__3982\
        );

    \I__746\ : InMux
    port map (
            O => \N__3991\,
            I => \N__3976\
        );

    \I__745\ : InMux
    port map (
            O => \N__3988\,
            I => \N__3976\
        );

    \I__744\ : InMux
    port map (
            O => \N__3987\,
            I => \N__3973\
        );

    \I__743\ : InMux
    port map (
            O => \N__3986\,
            I => \N__3964\
        );

    \I__742\ : InMux
    port map (
            O => \N__3985\,
            I => \N__3964\
        );

    \I__741\ : InMux
    port map (
            O => \N__3982\,
            I => \N__3964\
        );

    \I__740\ : InMux
    port map (
            O => \N__3981\,
            I => \N__3964\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3976\,
            I => \N__3961\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3973\,
            I => \U409_TICK.TICK603_10\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__3964\,
            I => \U409_TICK.TICK603_10\
        );

    \I__736\ : Odrv4
    port map (
            O => \N__3961\,
            I => \U409_TICK.TICK603_10\
        );

    \I__735\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3945\
        );

    \I__734\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3940\
        );

    \I__733\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3940\
        );

    \I__732\ : InMux
    port map (
            O => \N__3951\,
            I => \N__3937\
        );

    \I__731\ : InMux
    port map (
            O => \N__3950\,
            I => \N__3930\
        );

    \I__730\ : InMux
    port map (
            O => \N__3949\,
            I => \N__3930\
        );

    \I__729\ : InMux
    port map (
            O => \N__3948\,
            I => \N__3930\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3945\,
            I => \U409_TICK.TICK603_9\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__3940\,
            I => \U409_TICK.TICK603_9\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__3937\,
            I => \U409_TICK.TICK603_9\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__3930\,
            I => \U409_TICK.TICK603_9\
        );

    \I__724\ : InMux
    port map (
            O => \N__3921\,
            I => \N__3914\
        );

    \I__723\ : InMux
    port map (
            O => \N__3920\,
            I => \N__3911\
        );

    \I__722\ : InMux
    port map (
            O => \N__3919\,
            I => \N__3906\
        );

    \I__721\ : InMux
    port map (
            O => \N__3918\,
            I => \N__3901\
        );

    \I__720\ : InMux
    port map (
            O => \N__3917\,
            I => \N__3901\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3914\,
            I => \N__3896\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__3911\,
            I => \N__3896\
        );

    \I__717\ : InMux
    port map (
            O => \N__3910\,
            I => \N__3891\
        );

    \I__716\ : InMux
    port map (
            O => \N__3909\,
            I => \N__3891\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3906\,
            I => \U409_TICK.TICK603_14\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__3901\,
            I => \U409_TICK.TICK603_14\
        );

    \I__713\ : Odrv4
    port map (
            O => \N__3896\,
            I => \U409_TICK.TICK603_14\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__3891\,
            I => \U409_TICK.TICK603_14\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__3882\,
            I => \U409_TICK.TICK603_10_cascade_\
        );

    \I__710\ : InMux
    port map (
            O => \N__3879\,
            I => \N__3876\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3876\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__708\ : InMux
    port map (
            O => \N__3873\,
            I => \N__3869\
        );

    \I__707\ : InMux
    port map (
            O => \N__3872\,
            I => \N__3866\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3869\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3866\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__704\ : InMux
    port map (
            O => \N__3861\,
            I => \N__3858\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3858\,
            I => \N__3855\
        );

    \I__702\ : Odrv4
    port map (
            O => \N__3855\,
            I => \U409_TICK.TICK503_11\
        );

    \I__701\ : CascadeMux
    port map (
            O => \N__3852\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__3849\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\
        );

    \I__699\ : IoInMux
    port map (
            O => \N__3846\,
            I => \N__3843\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3843\,
            I => \N__3840\
        );

    \I__697\ : IoSpan4Mux
    port map (
            O => \N__3840\,
            I => \N__3837\
        );

    \I__696\ : Span4Mux_s3_v
    port map (
            O => \N__3837\,
            I => \N__3834\
        );

    \I__695\ : Span4Mux_v
    port map (
            O => \N__3834\,
            I => \N__3831\
        );

    \I__694\ : Sp12to4
    port map (
            O => \N__3831\,
            I => \N__3828\
        );

    \I__693\ : Span12Mux_v
    port map (
            O => \N__3828\,
            I => \N__3824\
        );

    \I__692\ : InMux
    port map (
            O => \N__3827\,
            I => \N__3821\
        );

    \I__691\ : Odrv12
    port map (
            O => \N__3824\,
            I => \TACK_OUTn\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3821\,
            I => \TACK_OUTn\
        );

    \I__689\ : InMux
    port map (
            O => \N__3816\,
            I => \N__3807\
        );

    \I__688\ : InMux
    port map (
            O => \N__3815\,
            I => \N__3807\
        );

    \I__687\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3807\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__3807\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__685\ : InMux
    port map (
            O => \N__3804\,
            I => \N__3795\
        );

    \I__684\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3795\
        );

    \I__683\ : InMux
    port map (
            O => \N__3802\,
            I => \N__3795\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__3795\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__681\ : CascadeMux
    port map (
            O => \N__3792\,
            I => \N__3789\
        );

    \I__680\ : InMux
    port map (
            O => \N__3789\,
            I => \N__3786\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3786\,
            I => \N__3783\
        );

    \I__678\ : Odrv4
    port map (
            O => \N__3783\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\
        );

    \I__677\ : InMux
    port map (
            O => \N__3780\,
            I => \N__3777\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3777\,
            I => \N__3774\
        );

    \I__675\ : Span4Mux_v
    port map (
            O => \N__3774\,
            I => \N__3771\
        );

    \I__674\ : Sp12to4
    port map (
            O => \N__3771\,
            I => \N__3768\
        );

    \I__673\ : Span12Mux_h
    port map (
            O => \N__3768\,
            I => \N__3765\
        );

    \I__672\ : Odrv12
    port map (
            O => \N__3765\,
            I => \A_c_13\
        );

    \I__671\ : IoInMux
    port map (
            O => \N__3762\,
            I => \N__3759\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3759\,
            I => \N__3756\
        );

    \I__669\ : Span4Mux_s2_h
    port map (
            O => \N__3756\,
            I => \N__3753\
        );

    \I__668\ : Span4Mux_v
    port map (
            O => \N__3753\,
            I => \N__3750\
        );

    \I__667\ : Span4Mux_h
    port map (
            O => \N__3750\,
            I => \N__3747\
        );

    \I__666\ : Sp12to4
    port map (
            O => \N__3747\,
            I => \N__3744\
        );

    \I__665\ : Span12Mux_h
    port map (
            O => \N__3744\,
            I => \N__3741\
        );

    \I__664\ : Odrv12
    port map (
            O => \N__3741\,
            I => \U409_ADDRESS_DECODE_un1_nCIACS1_i\
        );

    \I__663\ : InMux
    port map (
            O => \N__3738\,
            I => \N__3735\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3735\,
            I => \N__3732\
        );

    \I__661\ : Span4Mux_v
    port map (
            O => \N__3732\,
            I => \N__3729\
        );

    \I__660\ : Sp12to4
    port map (
            O => \N__3729\,
            I => \N__3726\
        );

    \I__659\ : Span12Mux_h
    port map (
            O => \N__3726\,
            I => \N__3723\
        );

    \I__658\ : Odrv12
    port map (
            O => \N__3723\,
            I => \A_c_12\
        );

    \I__657\ : IoInMux
    port map (
            O => \N__3720\,
            I => \N__3717\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3717\,
            I => \N__3714\
        );

    \I__655\ : Span4Mux_s0_h
    port map (
            O => \N__3714\,
            I => \N__3711\
        );

    \I__654\ : Sp12to4
    port map (
            O => \N__3711\,
            I => \N__3708\
        );

    \I__653\ : Span12Mux_s9_v
    port map (
            O => \N__3708\,
            I => \N__3705\
        );

    \I__652\ : Span12Mux_h
    port map (
            O => \N__3705\,
            I => \N__3702\
        );

    \I__651\ : Odrv12
    port map (
            O => \N__3702\,
            I => \U409_ADDRESS_DECODE_un1_nCIACS0_i\
        );

    \I__650\ : CascadeMux
    port map (
            O => \N__3699\,
            I => \N__3696\
        );

    \I__649\ : InMux
    port map (
            O => \N__3696\,
            I => \N__3692\
        );

    \I__648\ : InMux
    port map (
            O => \N__3695\,
            I => \N__3688\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3692\,
            I => \N__3685\
        );

    \I__646\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3682\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3688\,
            I => \N__3679\
        );

    \I__644\ : Span4Mux_h
    port map (
            O => \N__3685\,
            I => \N__3674\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__3682\,
            I => \N__3674\
        );

    \I__642\ : Span4Mux_v
    port map (
            O => \N__3679\,
            I => \N__3671\
        );

    \I__641\ : Span4Mux_v
    port map (
            O => \N__3674\,
            I => \N__3668\
        );

    \I__640\ : Sp12to4
    port map (
            O => \N__3671\,
            I => \N__3663\
        );

    \I__639\ : Sp12to4
    port map (
            O => \N__3668\,
            I => \N__3663\
        );

    \I__638\ : Span12Mux_h
    port map (
            O => \N__3663\,
            I => \N__3660\
        );

    \I__637\ : Span12Mux_v
    port map (
            O => \N__3660\,
            I => \N__3657\
        );

    \I__636\ : Odrv12
    port map (
            O => \N__3657\,
            I => \TSn_c\
        );

    \I__635\ : IoInMux
    port map (
            O => \N__3654\,
            I => \N__3648\
        );

    \I__634\ : InMux
    port map (
            O => \N__3653\,
            I => \N__3645\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__3652\,
            I => \N__3642\
        );

    \I__632\ : CascadeMux
    port map (
            O => \N__3651\,
            I => \N__3637\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3648\,
            I => \N__3634\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3645\,
            I => \N__3631\
        );

    \I__629\ : InMux
    port map (
            O => \N__3642\,
            I => \N__3628\
        );

    \I__628\ : InMux
    port map (
            O => \N__3641\,
            I => \N__3623\
        );

    \I__627\ : InMux
    port map (
            O => \N__3640\,
            I => \N__3623\
        );

    \I__626\ : InMux
    port map (
            O => \N__3637\,
            I => \N__3620\
        );

    \I__625\ : IoSpan4Mux
    port map (
            O => \N__3634\,
            I => \N__3617\
        );

    \I__624\ : Span4Mux_h
    port map (
            O => \N__3631\,
            I => \N__3612\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3628\,
            I => \N__3612\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3623\,
            I => \N__3607\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3620\,
            I => \N__3607\
        );

    \I__620\ : Span4Mux_s0_v
    port map (
            O => \N__3617\,
            I => \N__3604\
        );

    \I__619\ : Span4Mux_v
    port map (
            O => \N__3612\,
            I => \N__3601\
        );

    \I__618\ : Span4Mux_v
    port map (
            O => \N__3607\,
            I => \N__3598\
        );

    \I__617\ : Sp12to4
    port map (
            O => \N__3604\,
            I => \N__3595\
        );

    \I__616\ : Span4Mux_v
    port map (
            O => \N__3601\,
            I => \N__3592\
        );

    \I__615\ : Sp12to4
    port map (
            O => \N__3598\,
            I => \N__3589\
        );

    \I__614\ : Span12Mux_v
    port map (
            O => \N__3595\,
            I => \N__3586\
        );

    \I__613\ : Sp12to4
    port map (
            O => \N__3592\,
            I => \N__3583\
        );

    \I__612\ : Span12Mux_h
    port map (
            O => \N__3589\,
            I => \N__3580\
        );

    \I__611\ : Span12Mux_v
    port map (
            O => \N__3586\,
            I => \N__3577\
        );

    \I__610\ : Span12Mux_h
    port map (
            O => \N__3583\,
            I => \N__3574\
        );

    \I__609\ : Span12Mux_v
    port map (
            O => \N__3580\,
            I => \N__3571\
        );

    \I__608\ : Odrv12
    port map (
            O => \N__3577\,
            I => \CLK40_IN_c\
        );

    \I__607\ : Odrv12
    port map (
            O => \N__3574\,
            I => \CLK40_IN_c\
        );

    \I__606\ : Odrv12
    port map (
            O => \N__3571\,
            I => \CLK40_IN_c\
        );

    \I__605\ : InMux
    port map (
            O => \N__3564\,
            I => \N__3561\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3561\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__603\ : InMux
    port map (
            O => \N__3558\,
            I => \N__3554\
        );

    \I__602\ : InMux
    port map (
            O => \N__3557\,
            I => \N__3551\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3554\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3551\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__599\ : InMux
    port map (
            O => \N__3546\,
            I => \N__3542\
        );

    \I__598\ : InMux
    port map (
            O => \N__3545\,
            I => \N__3539\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3542\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3539\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__595\ : CascadeMux
    port map (
            O => \N__3534\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_\
        );

    \I__594\ : InMux
    port map (
            O => \N__3531\,
            I => \N__3527\
        );

    \I__593\ : InMux
    port map (
            O => \N__3530\,
            I => \N__3524\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3527\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3524\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__590\ : InMux
    port map (
            O => \N__3519\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__589\ : InMux
    port map (
            O => \N__3516\,
            I => \N__3512\
        );

    \I__588\ : InMux
    port map (
            O => \N__3515\,
            I => \N__3509\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3512\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__3509\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__585\ : InMux
    port map (
            O => \N__3504\,
            I => \N__3501\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3501\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__583\ : InMux
    port map (
            O => \N__3498\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__582\ : InMux
    port map (
            O => \N__3495\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__581\ : InMux
    port map (
            O => \N__3492\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__580\ : InMux
    port map (
            O => \N__3489\,
            I => \N__3485\
        );

    \I__579\ : InMux
    port map (
            O => \N__3488\,
            I => \N__3482\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3485\,
            I => \N__3479\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3482\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__576\ : Odrv4
    port map (
            O => \N__3479\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__575\ : InMux
    port map (
            O => \N__3474\,
            I => \N__3468\
        );

    \I__574\ : InMux
    port map (
            O => \N__3473\,
            I => \N__3461\
        );

    \I__573\ : InMux
    port map (
            O => \N__3472\,
            I => \N__3461\
        );

    \I__572\ : InMux
    port map (
            O => \N__3471\,
            I => \N__3461\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3468\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3461\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__569\ : SRMux
    port map (
            O => \N__3456\,
            I => \N__3453\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3453\,
            I => \N__3450\
        );

    \I__567\ : Span4Mux_h
    port map (
            O => \N__3450\,
            I => \N__3447\
        );

    \I__566\ : Odrv4
    port map (
            O => \N__3447\,
            I => \U409_TRANSFER_ACK.RESETn_c_i\
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__3444\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__3441\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__563\ : InMux
    port map (
            O => \N__3438\,
            I => \N__3434\
        );

    \I__562\ : InMux
    port map (
            O => \N__3437\,
            I => \N__3431\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3434\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3431\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__559\ : InMux
    port map (
            O => \N__3426\,
            I => \N__3423\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__3423\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__557\ : InMux
    port map (
            O => \N__3420\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__556\ : InMux
    port map (
            O => \N__3417\,
            I => \N__3413\
        );

    \I__555\ : InMux
    port map (
            O => \N__3416\,
            I => \N__3410\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3413\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3410\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__552\ : InMux
    port map (
            O => \N__3405\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__3402\,
            I => \N__3398\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__3401\,
            I => \N__3395\
        );

    \I__549\ : InMux
    port map (
            O => \N__3398\,
            I => \N__3392\
        );

    \I__548\ : InMux
    port map (
            O => \N__3395\,
            I => \N__3389\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3392\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3389\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__545\ : InMux
    port map (
            O => \N__3384\,
            I => \N__3381\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3381\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__543\ : InMux
    port map (
            O => \N__3378\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__542\ : InMux
    port map (
            O => \N__3375\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__541\ : InMux
    port map (
            O => \N__3372\,
            I => \N__3368\
        );

    \I__540\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3365\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3368\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3365\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__537\ : CascadeMux
    port map (
            O => \N__3360\,
            I => \N__3357\
        );

    \I__536\ : InMux
    port map (
            O => \N__3357\,
            I => \N__3354\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3354\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__534\ : InMux
    port map (
            O => \N__3351\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__533\ : InMux
    port map (
            O => \N__3348\,
            I => \N__3344\
        );

    \I__532\ : InMux
    port map (
            O => \N__3347\,
            I => \N__3341\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3344\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3341\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__529\ : InMux
    port map (
            O => \N__3336\,
            I => \N__3333\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3333\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__527\ : InMux
    port map (
            O => \N__3330\,
            I => \bfn_10_7_0_\
        );

    \I__526\ : InMux
    port map (
            O => \N__3327\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__525\ : InMux
    port map (
            O => \N__3324\,
            I => \N__3321\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3321\,
            I => \N__3317\
        );

    \I__523\ : InMux
    port map (
            O => \N__3320\,
            I => \N__3314\
        );

    \I__522\ : Odrv4
    port map (
            O => \N__3317\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3314\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__520\ : InMux
    port map (
            O => \N__3309\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__519\ : InMux
    port map (
            O => \N__3306\,
            I => \N__3302\
        );

    \I__518\ : InMux
    port map (
            O => \N__3305\,
            I => \N__3299\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3302\,
            I => \N__3296\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3299\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__515\ : Odrv4
    port map (
            O => \N__3296\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__514\ : InMux
    port map (
            O => \N__3291\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__3288\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__3285\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__511\ : IoInMux
    port map (
            O => \N__3282\,
            I => \N__3279\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3279\,
            I => \N__3276\
        );

    \I__509\ : Span4Mux_s2_v
    port map (
            O => \N__3276\,
            I => \N__3273\
        );

    \I__508\ : Span4Mux_v
    port map (
            O => \N__3273\,
            I => \N__3270\
        );

    \I__507\ : Span4Mux_v
    port map (
            O => \N__3270\,
            I => \N__3267\
        );

    \I__506\ : Span4Mux_h
    port map (
            O => \N__3267\,
            I => \N__3263\
        );

    \I__505\ : InMux
    port map (
            O => \N__3266\,
            I => \N__3260\
        );

    \I__504\ : Odrv4
    port map (
            O => \N__3263\,
            I => \TICK60_c\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3260\,
            I => \TICK60_c\
        );

    \I__502\ : InMux
    port map (
            O => \N__3255\,
            I => \N__3252\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3252\,
            I => \U409_TICK.TICK603_8\
        );

    \I__500\ : InMux
    port map (
            O => \N__3249\,
            I => \N__3245\
        );

    \I__499\ : InMux
    port map (
            O => \N__3248\,
            I => \N__3242\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3245\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3242\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__496\ : InMux
    port map (
            O => \N__3237\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__495\ : InMux
    port map (
            O => \N__3234\,
            I => \N__3230\
        );

    \I__494\ : InMux
    port map (
            O => \N__3233\,
            I => \N__3227\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3230\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3227\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__491\ : InMux
    port map (
            O => \N__3222\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__3219\,
            I => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0_cascade_\
        );

    \I__489\ : InMux
    port map (
            O => \N__3216\,
            I => \N__3213\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3213\,
            I => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa\
        );

    \I__487\ : InMux
    port map (
            O => \N__3210\,
            I => \N__3207\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3207\,
            I => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0\
        );

    \I__485\ : CascadeMux
    port map (
            O => \N__3204\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_\
        );

    \I__484\ : InMux
    port map (
            O => \N__3201\,
            I => \N__3189\
        );

    \I__483\ : InMux
    port map (
            O => \N__3200\,
            I => \N__3189\
        );

    \I__482\ : InMux
    port map (
            O => \N__3199\,
            I => \N__3189\
        );

    \I__481\ : InMux
    port map (
            O => \N__3198\,
            I => \N__3189\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3189\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__479\ : CascadeMux
    port map (
            O => \N__3186\,
            I => \N__3180\
        );

    \I__478\ : InMux
    port map (
            O => \N__3185\,
            I => \N__3174\
        );

    \I__477\ : InMux
    port map (
            O => \N__3184\,
            I => \N__3174\
        );

    \I__476\ : InMux
    port map (
            O => \N__3183\,
            I => \N__3167\
        );

    \I__475\ : InMux
    port map (
            O => \N__3180\,
            I => \N__3167\
        );

    \I__474\ : InMux
    port map (
            O => \N__3179\,
            I => \N__3167\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3174\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3167\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__471\ : InMux
    port map (
            O => \N__3162\,
            I => \N__3159\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3159\,
            I => \N__3156\
        );

    \I__469\ : Span12Mux_h
    port map (
            O => \N__3156\,
            I => \N__3153\
        );

    \I__468\ : Odrv12
    port map (
            O => \N__3153\,
            I => \U409_ADDRESS_DECODE.HIROMZ0\
        );

    \I__467\ : InMux
    port map (
            O => \N__3150\,
            I => \N__3147\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3147\,
            I => \U409_ADDRESS_DECODE_un1_ROMEN_0\
        );

    \I__465\ : CascadeMux
    port map (
            O => \N__3144\,
            I => \U409_ADDRESS_DECODE_un1_ROMEN_0_cascade_\
        );

    \I__464\ : IoInMux
    port map (
            O => \N__3141\,
            I => \N__3138\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__3138\,
            I => \N__3135\
        );

    \I__462\ : Span4Mux_s0_v
    port map (
            O => \N__3135\,
            I => \N__3132\
        );

    \I__461\ : Span4Mux_v
    port map (
            O => \N__3132\,
            I => \N__3129\
        );

    \I__460\ : Sp12to4
    port map (
            O => \N__3129\,
            I => \N__3126\
        );

    \I__459\ : Span12Mux_h
    port map (
            O => \N__3126\,
            I => \N__3123\
        );

    \I__458\ : Odrv12
    port map (
            O => \N__3123\,
            I => \ROMENm_i\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__3120\,
            I => \U409_TICK.TICK603_11_cascade_\
        );

    \I__456\ : CascadeMux
    port map (
            O => \N__3117\,
            I => \U409_TRANSFER_ACK.m9_bm_cascade_\
        );

    \I__455\ : InMux
    port map (
            O => \N__3114\,
            I => \N__3111\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__3111\,
            I => \U409_TRANSFER_ACK.N_4\
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__3108\,
            I => \N__3104\
        );

    \I__452\ : CascadeMux
    port map (
            O => \N__3107\,
            I => \N__3101\
        );

    \I__451\ : InMux
    port map (
            O => \N__3104\,
            I => \N__3093\
        );

    \I__450\ : InMux
    port map (
            O => \N__3101\,
            I => \N__3093\
        );

    \I__449\ : InMux
    port map (
            O => \N__3100\,
            I => \N__3093\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3093\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__3090\,
            I => \U409_TRANSFER_ACK.N_4_cascade_\
        );

    \I__446\ : InMux
    port map (
            O => \N__3087\,
            I => \N__3084\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3084\,
            I => \U409_TRANSFER_ACK.m9_am\
        );

    \I__444\ : InMux
    port map (
            O => \N__3081\,
            I => \N__3077\
        );

    \I__443\ : InMux
    port map (
            O => \N__3080\,
            I => \N__3074\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__3077\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3074\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__440\ : InMux
    port map (
            O => \N__3069\,
            I => \N__3064\
        );

    \I__439\ : InMux
    port map (
            O => \N__3068\,
            I => \N__3059\
        );

    \I__438\ : InMux
    port map (
            O => \N__3067\,
            I => \N__3059\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__3064\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3059\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__435\ : InMux
    port map (
            O => \N__3054\,
            I => \N__3048\
        );

    \I__434\ : InMux
    port map (
            O => \N__3053\,
            I => \N__3040\
        );

    \I__433\ : InMux
    port map (
            O => \N__3052\,
            I => \N__3040\
        );

    \I__432\ : InMux
    port map (
            O => \N__3051\,
            I => \N__3040\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3048\,
            I => \N__3037\
        );

    \I__430\ : InMux
    port map (
            O => \N__3047\,
            I => \N__3034\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3040\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__428\ : Odrv4
    port map (
            O => \N__3037\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3034\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__426\ : InMux
    port map (
            O => \N__3027\,
            I => \N__3023\
        );

    \I__425\ : InMux
    port map (
            O => \N__3026\,
            I => \N__3020\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3023\,
            I => \U409_TRANSFER_ACK.N_97\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__3020\,
            I => \U409_TRANSFER_ACK.N_97\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__3015\,
            I => \N__3012\
        );

    \I__421\ : InMux
    port map (
            O => \N__3012\,
            I => \N__3008\
        );

    \I__420\ : InMux
    port map (
            O => \N__3011\,
            I => \N__3003\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3008\,
            I => \N__3000\
        );

    \I__418\ : InMux
    port map (
            O => \N__3007\,
            I => \N__2995\
        );

    \I__417\ : InMux
    port map (
            O => \N__3006\,
            I => \N__2995\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3003\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__415\ : Odrv4
    port map (
            O => \N__3000\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2995\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__2988\,
            I => \U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_\
        );

    \I__412\ : CascadeMux
    port map (
            O => \N__2985\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0_cascade_\
        );

    \I__411\ : InMux
    port map (
            O => \N__2982\,
            I => \N__2979\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__2979\,
            I => \N__2976\
        );

    \I__409\ : Odrv12
    port map (
            O => \N__2976\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\
        );

    \I__408\ : IoInMux
    port map (
            O => \N__2973\,
            I => \N__2970\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2970\,
            I => \N__2967\
        );

    \I__406\ : IoSpan4Mux
    port map (
            O => \N__2967\,
            I => \N__2964\
        );

    \I__405\ : Span4Mux_s0_v
    port map (
            O => \N__2964\,
            I => \N__2961\
        );

    \I__404\ : Span4Mux_v
    port map (
            O => \N__2961\,
            I => \N__2958\
        );

    \I__403\ : Sp12to4
    port map (
            O => \N__2958\,
            I => \N__2955\
        );

    \I__402\ : Odrv12
    port map (
            O => \N__2955\,
            I => \PORTSIZE_0_i\
        );

    \I__401\ : InMux
    port map (
            O => \N__2952\,
            I => \N__2949\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2949\,
            I => \N__2946\
        );

    \I__399\ : Span4Mux_v
    port map (
            O => \N__2946\,
            I => \N__2942\
        );

    \I__398\ : InMux
    port map (
            O => \N__2945\,
            I => \N__2939\
        );

    \I__397\ : Sp12to4
    port map (
            O => \N__2942\,
            I => \N__2934\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2939\,
            I => \N__2934\
        );

    \I__395\ : Odrv12
    port map (
            O => \N__2934\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\
        );

    \I__394\ : CascadeMux
    port map (
            O => \N__2931\,
            I => \N__2925\
        );

    \I__393\ : InMux
    port map (
            O => \N__2930\,
            I => \N__2918\
        );

    \I__392\ : InMux
    port map (
            O => \N__2929\,
            I => \N__2918\
        );

    \I__391\ : InMux
    port map (
            O => \N__2928\,
            I => \N__2915\
        );

    \I__390\ : InMux
    port map (
            O => \N__2925\,
            I => \N__2910\
        );

    \I__389\ : InMux
    port map (
            O => \N__2924\,
            I => \N__2910\
        );

    \I__388\ : InMux
    port map (
            O => \N__2923\,
            I => \N__2907\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2918\,
            I => \N__2902\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2915\,
            I => \N__2902\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2910\,
            I => \N__2899\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__2907\,
            I => \N__2896\
        );

    \I__383\ : Span4Mux_v
    port map (
            O => \N__2902\,
            I => \N__2893\
        );

    \I__382\ : Span4Mux_v
    port map (
            O => \N__2899\,
            I => \N__2890\
        );

    \I__381\ : Span4Mux_v
    port map (
            O => \N__2896\,
            I => \N__2887\
        );

    \I__380\ : Sp12to4
    port map (
            O => \N__2893\,
            I => \N__2884\
        );

    \I__379\ : Span4Mux_h
    port map (
            O => \N__2890\,
            I => \N__2881\
        );

    \I__378\ : Span4Mux_h
    port map (
            O => \N__2887\,
            I => \N__2878\
        );

    \I__377\ : Odrv12
    port map (
            O => \N__2884\,
            I => \A_c_23\
        );

    \I__376\ : Odrv4
    port map (
            O => \N__2881\,
            I => \A_c_23\
        );

    \I__375\ : Odrv4
    port map (
            O => \N__2878\,
            I => \A_c_23\
        );

    \I__374\ : IoInMux
    port map (
            O => \N__2871\,
            I => \N__2868\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2868\,
            I => \N__2865\
        );

    \I__372\ : IoSpan4Mux
    port map (
            O => \N__2865\,
            I => \N__2862\
        );

    \I__371\ : IoSpan4Mux
    port map (
            O => \N__2862\,
            I => \N__2859\
        );

    \I__370\ : Span4Mux_s2_v
    port map (
            O => \N__2859\,
            I => \N__2856\
        );

    \I__369\ : Sp12to4
    port map (
            O => \N__2856\,
            I => \N__2853\
        );

    \I__368\ : Span12Mux_v
    port map (
            O => \N__2853\,
            I => \N__2850\
        );

    \I__367\ : Odrv12
    port map (
            O => \N__2850\,
            I => \U409_ADDRESS_DECODE_un1_nREGSPACE_i\
        );

    \I__366\ : CascadeMux
    port map (
            O => \N__2847\,
            I => \U409_TRANSFER_ACK.i6_mux_0_cascade_\
        );

    \I__365\ : CascadeMux
    port map (
            O => \N__2844\,
            I => \U409_CIA.g0Z0Z_2_cascade_\
        );

    \I__364\ : InMux
    port map (
            O => \N__2841\,
            I => \N__2835\
        );

    \I__363\ : InMux
    port map (
            O => \N__2840\,
            I => \N__2835\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2835\,
            I => \N__2832\
        );

    \I__361\ : Span4Mux_v
    port map (
            O => \N__2832\,
            I => \N__2829\
        );

    \I__360\ : Span4Mux_h
    port map (
            O => \N__2829\,
            I => \N__2826\
        );

    \I__359\ : Odrv4
    port map (
            O => \N__2826\,
            I => \A_c_30\
        );

    \I__358\ : InMux
    port map (
            O => \N__2823\,
            I => \N__2817\
        );

    \I__357\ : InMux
    port map (
            O => \N__2822\,
            I => \N__2817\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2817\,
            I => \N__2814\
        );

    \I__355\ : Span4Mux_v
    port map (
            O => \N__2814\,
            I => \N__2811\
        );

    \I__354\ : Span4Mux_v
    port map (
            O => \N__2811\,
            I => \N__2808\
        );

    \I__353\ : Sp12to4
    port map (
            O => \N__2808\,
            I => \N__2805\
        );

    \I__352\ : Odrv12
    port map (
            O => \N__2805\,
            I => \A_c_28\
        );

    \I__351\ : InMux
    port map (
            O => \N__2802\,
            I => \N__2796\
        );

    \I__350\ : InMux
    port map (
            O => \N__2801\,
            I => \N__2796\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2796\,
            I => \N__2793\
        );

    \I__348\ : Span4Mux_h
    port map (
            O => \N__2793\,
            I => \N__2790\
        );

    \I__347\ : Span4Mux_v
    port map (
            O => \N__2790\,
            I => \N__2787\
        );

    \I__346\ : Odrv4
    port map (
            O => \N__2787\,
            I => \A_c_29\
        );

    \I__345\ : CascadeMux
    port map (
            O => \N__2784\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_\
        );

    \I__344\ : InMux
    port map (
            O => \N__2781\,
            I => \N__2778\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2778\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\
        );

    \I__342\ : InMux
    port map (
            O => \N__2775\,
            I => \N__2769\
        );

    \I__341\ : InMux
    port map (
            O => \N__2774\,
            I => \N__2769\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2769\,
            I => \N__2766\
        );

    \I__339\ : Span4Mux_h
    port map (
            O => \N__2766\,
            I => \N__2763\
        );

    \I__338\ : Span4Mux_v
    port map (
            O => \N__2763\,
            I => \N__2760\
        );

    \I__337\ : Odrv4
    port map (
            O => \N__2760\,
            I => \A_c_24\
        );

    \I__336\ : CascadeMux
    port map (
            O => \N__2757\,
            I => \N__2753\
        );

    \I__335\ : InMux
    port map (
            O => \N__2756\,
            I => \N__2748\
        );

    \I__334\ : InMux
    port map (
            O => \N__2753\,
            I => \N__2748\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2748\,
            I => \N__2745\
        );

    \I__332\ : Span4Mux_v
    port map (
            O => \N__2745\,
            I => \N__2742\
        );

    \I__331\ : Span4Mux_v
    port map (
            O => \N__2742\,
            I => \N__2739\
        );

    \I__330\ : Sp12to4
    port map (
            O => \N__2739\,
            I => \N__2736\
        );

    \I__329\ : Odrv12
    port map (
            O => \N__2736\,
            I => \A_c_26\
        );

    \I__328\ : CascadeMux
    port map (
            O => \N__2733\,
            I => \N__2730\
        );

    \I__327\ : InMux
    port map (
            O => \N__2730\,
            I => \N__2724\
        );

    \I__326\ : InMux
    port map (
            O => \N__2729\,
            I => \N__2724\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2724\,
            I => \N__2721\
        );

    \I__324\ : Span4Mux_v
    port map (
            O => \N__2721\,
            I => \N__2718\
        );

    \I__323\ : Sp12to4
    port map (
            O => \N__2718\,
            I => \N__2715\
        );

    \I__322\ : Odrv12
    port map (
            O => \N__2715\,
            I => \A_c_31\
        );

    \I__321\ : InMux
    port map (
            O => \N__2712\,
            I => \N__2708\
        );

    \I__320\ : InMux
    port map (
            O => \N__2711\,
            I => \N__2705\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2708\,
            I => \N__2700\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2705\,
            I => \N__2700\
        );

    \I__317\ : Span4Mux_v
    port map (
            O => \N__2700\,
            I => \N__2697\
        );

    \I__316\ : Span4Mux_h
    port map (
            O => \N__2697\,
            I => \N__2694\
        );

    \I__315\ : Odrv4
    port map (
            O => \N__2694\,
            I => \A_c_27\
        );

    \I__314\ : InMux
    port map (
            O => \N__2691\,
            I => \N__2688\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2688\,
            I => \U409_CIA.g0Z0Z_10\
        );

    \I__312\ : InMux
    port map (
            O => \N__2685\,
            I => \N__2674\
        );

    \I__311\ : InMux
    port map (
            O => \N__2684\,
            I => \N__2674\
        );

    \I__310\ : InMux
    port map (
            O => \N__2683\,
            I => \N__2674\
        );

    \I__309\ : InMux
    port map (
            O => \N__2682\,
            I => \N__2671\
        );

    \I__308\ : InMux
    port map (
            O => \N__2681\,
            I => \N__2668\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2674\,
            I => \N__2665\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2671\,
            I => \N__2662\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2668\,
            I => \N__2655\
        );

    \I__304\ : Sp12to4
    port map (
            O => \N__2665\,
            I => \N__2655\
        );

    \I__303\ : Sp12to4
    port map (
            O => \N__2662\,
            I => \N__2655\
        );

    \I__302\ : Span12Mux_v
    port map (
            O => \N__2655\,
            I => \N__2652\
        );

    \I__301\ : Odrv12
    port map (
            O => \N__2652\,
            I => \A_c_22\
        );

    \I__300\ : InMux
    port map (
            O => \N__2649\,
            I => \N__2641\
        );

    \I__299\ : InMux
    port map (
            O => \N__2648\,
            I => \N__2641\
        );

    \I__298\ : InMux
    port map (
            O => \N__2647\,
            I => \N__2636\
        );

    \I__297\ : InMux
    port map (
            O => \N__2646\,
            I => \N__2636\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2641\,
            I => \N__2633\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2636\,
            I => \N__2630\
        );

    \I__294\ : Span4Mux_v
    port map (
            O => \N__2633\,
            I => \N__2627\
        );

    \I__293\ : Span12Mux_v
    port map (
            O => \N__2630\,
            I => \N__2624\
        );

    \I__292\ : Span4Mux_h
    port map (
            O => \N__2627\,
            I => \N__2621\
        );

    \I__291\ : Odrv12
    port map (
            O => \N__2624\,
            I => \A_c_21\
        );

    \I__290\ : Odrv4
    port map (
            O => \N__2621\,
            I => \A_c_21\
        );

    \I__289\ : CascadeMux
    port map (
            O => \N__2616\,
            I => \N__2613\
        );

    \I__288\ : InMux
    port map (
            O => \N__2613\,
            I => \N__2610\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__2610\,
            I => \N__2607\
        );

    \I__286\ : Span4Mux_v
    port map (
            O => \N__2607\,
            I => \N__2604\
        );

    \I__285\ : Odrv4
    port map (
            O => \N__2604\,
            I => \U409_CIA.g0Z0Z_8\
        );

    \I__284\ : CascadeMux
    port map (
            O => \N__2601\,
            I => \N__2598\
        );

    \I__283\ : InMux
    port map (
            O => \N__2598\,
            I => \N__2592\
        );

    \I__282\ : InMux
    port map (
            O => \N__2597\,
            I => \N__2592\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2592\,
            I => \N__2589\
        );

    \I__280\ : Span4Mux_v
    port map (
            O => \N__2589\,
            I => \N__2586\
        );

    \I__279\ : Span4Mux_h
    port map (
            O => \N__2586\,
            I => \N__2583\
        );

    \I__278\ : Span4Mux_v
    port map (
            O => \N__2583\,
            I => \N__2580\
        );

    \I__277\ : Odrv4
    port map (
            O => \N__2580\,
            I => \A_c_16\
        );

    \I__276\ : CascadeMux
    port map (
            O => \N__2577\,
            I => \N__2573\
        );

    \I__275\ : InMux
    port map (
            O => \N__2576\,
            I => \N__2570\
        );

    \I__274\ : InMux
    port map (
            O => \N__2573\,
            I => \N__2567\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__2570\,
            I => \N__2564\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2567\,
            I => \N__2561\
        );

    \I__271\ : Span4Mux_v
    port map (
            O => \N__2564\,
            I => \N__2556\
        );

    \I__270\ : Span4Mux_v
    port map (
            O => \N__2561\,
            I => \N__2556\
        );

    \I__269\ : Span4Mux_h
    port map (
            O => \N__2556\,
            I => \N__2553\
        );

    \I__268\ : Span4Mux_v
    port map (
            O => \N__2553\,
            I => \N__2550\
        );

    \I__267\ : Span4Mux_v
    port map (
            O => \N__2550\,
            I => \N__2547\
        );

    \I__266\ : Odrv4
    port map (
            O => \N__2547\,
            I => \A_c_18\
        );

    \I__265\ : InMux
    port map (
            O => \N__2544\,
            I => \N__2541\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2541\,
            I => \U409_CIA.g0Z0Z_11\
        );

    \I__263\ : InMux
    port map (
            O => \N__2538\,
            I => \N__2534\
        );

    \I__262\ : InMux
    port map (
            O => \N__2537\,
            I => \N__2531\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2534\,
            I => \N__2526\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2531\,
            I => \N__2526\
        );

    \I__259\ : Sp12to4
    port map (
            O => \N__2526\,
            I => \N__2523\
        );

    \I__258\ : Span12Mux_v
    port map (
            O => \N__2523\,
            I => \N__2520\
        );

    \I__257\ : Odrv12
    port map (
            O => \N__2520\,
            I => \A_c_17\
        );

    \I__256\ : CascadeMux
    port map (
            O => \N__2517\,
            I => \U409_ADDRESS_DECODE.HIROM_0_cascade_\
        );

    \I__255\ : InMux
    port map (
            O => \N__2514\,
            I => \N__2511\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2511\,
            I => \N__2508\
        );

    \I__253\ : Span4Mux_v
    port map (
            O => \N__2508\,
            I => \N__2505\
        );

    \I__252\ : Span4Mux_v
    port map (
            O => \N__2505\,
            I => \N__2500\
        );

    \I__251\ : InMux
    port map (
            O => \N__2504\,
            I => \N__2495\
        );

    \I__250\ : InMux
    port map (
            O => \N__2503\,
            I => \N__2495\
        );

    \I__249\ : Sp12to4
    port map (
            O => \N__2500\,
            I => \N__2492\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__2495\,
            I => \N__2489\
        );

    \I__247\ : Span12Mux_s3_h
    port map (
            O => \N__2492\,
            I => \N__2484\
        );

    \I__246\ : Span12Mux_h
    port map (
            O => \N__2489\,
            I => \N__2484\
        );

    \I__245\ : Span12Mux_v
    port map (
            O => \N__2484\,
            I => \N__2481\
        );

    \I__244\ : Odrv12
    port map (
            O => \N__2481\,
            I => \A_c_19\
        );

    \I__243\ : CascadeMux
    port map (
            O => \N__2478\,
            I => \N__2475\
        );

    \I__242\ : InMux
    port map (
            O => \N__2475\,
            I => \N__2472\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__2472\,
            I => \U409_ADDRESS_DECODE.HIROM_0\
        );

    \I__240\ : InMux
    port map (
            O => \N__2469\,
            I => \N__2466\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__2466\,
            I => \N__2463\
        );

    \I__238\ : Span4Mux_h
    port map (
            O => \N__2463\,
            I => \N__2460\
        );

    \I__237\ : Span4Mux_v
    port map (
            O => \N__2460\,
            I => \N__2455\
        );

    \I__236\ : InMux
    port map (
            O => \N__2459\,
            I => \N__2450\
        );

    \I__235\ : InMux
    port map (
            O => \N__2458\,
            I => \N__2450\
        );

    \I__234\ : Sp12to4
    port map (
            O => \N__2455\,
            I => \N__2445\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__2450\,
            I => \N__2445\
        );

    \I__232\ : Odrv12
    port map (
            O => \N__2445\,
            I => \A_c_20\
        );

    \I__231\ : CascadeMux
    port map (
            O => \N__2442\,
            I => \N__2439\
        );

    \I__230\ : InMux
    port map (
            O => \N__2439\,
            I => \N__2436\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__2436\,
            I => \N__2432\
        );

    \I__228\ : InMux
    port map (
            O => \N__2435\,
            I => \N__2429\
        );

    \I__227\ : Sp12to4
    port map (
            O => \N__2432\,
            I => \N__2424\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__2429\,
            I => \N__2424\
        );

    \I__225\ : Odrv12
    port map (
            O => \N__2424\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEm_6\
        );

    \I__224\ : InMux
    port map (
            O => \N__2421\,
            I => \N__2418\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__2418\,
            I => \N__2415\
        );

    \I__222\ : Span4Mux_v
    port map (
            O => \N__2415\,
            I => \N__2411\
        );

    \I__221\ : InMux
    port map (
            O => \N__2414\,
            I => \N__2408\
        );

    \I__220\ : Span4Mux_v
    port map (
            O => \N__2411\,
            I => \N__2405\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__2408\,
            I => \N__2402\
        );

    \I__218\ : Span4Mux_v
    port map (
            O => \N__2405\,
            I => \N__2397\
        );

    \I__217\ : Span4Mux_v
    port map (
            O => \N__2402\,
            I => \N__2397\
        );

    \I__216\ : Span4Mux_h
    port map (
            O => \N__2397\,
            I => \N__2394\
        );

    \I__215\ : Odrv4
    port map (
            O => \N__2394\,
            I => \A_c_25\
        );

    \I__214\ : ClkMux
    port map (
            O => \N__2391\,
            I => \N__2364\
        );

    \I__213\ : ClkMux
    port map (
            O => \N__2390\,
            I => \N__2364\
        );

    \I__212\ : ClkMux
    port map (
            O => \N__2389\,
            I => \N__2364\
        );

    \I__211\ : ClkMux
    port map (
            O => \N__2388\,
            I => \N__2364\
        );

    \I__210\ : ClkMux
    port map (
            O => \N__2387\,
            I => \N__2364\
        );

    \I__209\ : ClkMux
    port map (
            O => \N__2386\,
            I => \N__2364\
        );

    \I__208\ : ClkMux
    port map (
            O => \N__2385\,
            I => \N__2364\
        );

    \I__207\ : ClkMux
    port map (
            O => \N__2384\,
            I => \N__2364\
        );

    \I__206\ : ClkMux
    port map (
            O => \N__2383\,
            I => \N__2364\
        );

    \I__205\ : GlobalMux
    port map (
            O => \N__2364\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.TACK_EN_iC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            I => \N__2389\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            I => \N__2386\
        );

    \INVU409_TRANSFER_ACK.TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            I => \N__2390\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            I => \N__2388\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            I => \N__2385\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            I => \N__2383\
        );

    \INVU409_TRANSFER_ACK.CIA_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            I => \N__2391\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            I => \N__2387\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            I => \N__2384\
        );

    \IN_MUX_bfv_10_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_6_0_\
        );

    \IN_MUX_bfv_10_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_10_7_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_12_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_12_7_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_9_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2597\,
            in1 => \N__2503\,
            in2 => \N__2577\,
            in3 => \N__2537\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_11_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2421\,
            in1 => \N__2504\,
            in2 => \N__2601\,
            in3 => \N__2576\,
            lcout => \U409_CIA.g0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_14_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2544\,
            in1 => \N__2469\,
            in2 => \N__2616\,
            in3 => \N__2538\,
            lcout => \U409_CIA.g0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2648\,
            in2 => \_gnd_net_\,
            in3 => \N__2458\,
            lcout => \U409_ADDRESS_DECODE.HIROM_0\,
            ltout => \U409_ADDRESS_DECODE.HIROM_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.HIROM_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2923\,
            in1 => \N__2684\,
            in2 => \N__2517\,
            in3 => \N__2514\,
            lcout => \U409_ADDRESS_DECODE.HIROMZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2683\,
            in1 => \N__4475\,
            in2 => \N__2478\,
            in3 => \N__2435\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__2685\,
            in1 => \N__2459\,
            in2 => \N__2442\,
            in3 => \N__2649\,
            lcout => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2414\,
            in1 => \N__2711\,
            in2 => \N__2757\,
            in3 => \N__2774\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_2_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__2802\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2841\,
            lcout => OPEN,
            ltout => \U409_CIA.g0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_13_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__2823\,
            in1 => \N__2691\,
            in2 => \N__2844\,
            in3 => \N__2682\,
            lcout => \U409_CIA.g0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__2729\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2840\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__2822\,
            in1 => \N__2801\,
            in2 => \N__2784\,
            in3 => \N__2781\,
            lcout => \U409_ADDRESS_DECODE_Z2_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_10_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2775\,
            in1 => \N__2756\,
            in2 => \N__2733\,
            in3 => \N__2712\,
            lcout => \U409_CIA.g0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__2681\,
            in1 => \N__2924\,
            in2 => \_gnd_net_\,
            in3 => \N__2646\,
            lcout => \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_8_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__2647\,
            in1 => \_gnd_net_\,
            in2 => \N__2931\,
            in3 => \N__5469\,
            lcout => \U409_CIA.g0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2930\,
            in1 => \N__2945\,
            in2 => \_gnd_net_\,
            in3 => \N__4523\,
            lcout => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\,
            ltout => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5468\,
            in1 => \N__2929\,
            in2 => \N__2985\,
            in3 => \N__2982\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__2952\,
            in1 => \N__2928\,
            in2 => \_gnd_net_\,
            in3 => \N__4516\,
            lcout => \U409_ADDRESS_DECODE_un1_nREGSPACE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3953\,
            in1 => \N__3918\,
            in2 => \N__3996\,
            in3 => \N__3336\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3952\,
            in1 => \N__3917\,
            in2 => \N__3995\,
            in3 => \N__3504\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5429\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5470\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3474\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100110011"
        )
    port map (
            in0 => \N__3473\,
            in1 => \N__3114\,
            in2 => \N__3108\,
            in3 => \N__3051\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.i6_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010001000"
        )
    port map (
            in0 => \N__3052\,
            in1 => \N__5472\,
            in2 => \N__2847\,
            in3 => \N__3011\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5474\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3068\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4307\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5473\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000110111"
        )
    port map (
            in0 => \N__3472\,
            in1 => \N__3007\,
            in2 => \N__3107\,
            in3 => \N__3027\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.m9_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100001001100"
        )
    port map (
            in0 => \N__3053\,
            in1 => \N__5471\,
            in2 => \N__3117\,
            in3 => \N__3087\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3080\,
            in2 => \_gnd_net_\,
            in3 => \N__3067\,
            lcout => \U409_TRANSFER_ACK.N_4\,
            ltout => \U409_TRANSFER_ACK.N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000111110101"
        )
    port map (
            in0 => \N__3006\,
            in1 => \N__3100\,
            in2 => \N__3090\,
            in3 => \N__3471\,
            lcout => \U409_TRANSFER_ACK.m9_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__3047\,
            in1 => \N__3081\,
            in2 => \N__3651\,
            in3 => \N__3069\,
            lcout => \U409_TRANSFER_ACK.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100001000"
        )
    port map (
            in0 => \N__3054\,
            in1 => \N__3026\,
            in2 => \N__3015\,
            in3 => \N__3546\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5475\,
            in2 => \N__2988\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000000100000"
        )
    port map (
            in0 => \N__3184\,
            in1 => \N__3200\,
            in2 => \N__5486\,
            in3 => \N__3216\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__3150\,
            in1 => \N__5480\,
            in2 => \N__4530\,
            in3 => \N__3691\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0\,
            ltout => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3640\,
            in1 => \N__3179\,
            in2 => \N__3219\,
            in3 => \N__3198\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000110100101"
        )
    port map (
            in0 => \N__3199\,
            in1 => \N__3210\,
            in2 => \N__3186\,
            in3 => \N__3641\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__5481\,
            in1 => \N__3183\,
            in2 => \N__3204\,
            in3 => \N__3531\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__3201\,
            in1 => \N__5479\,
            in2 => \_gnd_net_\,
            in3 => \N__3185\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_ROMEN_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__4449\,
            in1 => \N__4402\,
            in2 => \_gnd_net_\,
            in3 => \N__3162\,
            lcout => \U409_ADDRESS_DECODE_un1_ROMEN_0\,
            ltout => \U409_ADDRESS_DECODE_un1_ROMEN_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMENm_i_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__4526\,
            in1 => \_gnd_net_\,
            in2 => \N__3144\,
            in3 => \N__5487\,
            lcout => \ROMENm_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3306\,
            in1 => \N__3249\,
            in2 => \N__4056\,
            in3 => \N__3489\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3255\,
            in1 => \N__3324\,
            in2 => \N__3120\,
            in3 => \N__3234\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3981\,
            in1 => \N__3948\,
            in2 => \N__3288\,
            in3 => \N__3426\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3348\,
            in1 => \N__3372\,
            in2 => \N__3402\,
            in3 => \N__3516\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__3985\,
            in1 => \N__3920\,
            in2 => \N__3285\,
            in3 => \N__3266\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3950\,
            in1 => \N__3910\,
            in2 => \N__3360\,
            in3 => \N__3986\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3909\,
            in1 => \N__3949\,
            in2 => \N__3994\,
            in3 => \N__3384\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__3417\,
            in1 => \N__3438\,
            in2 => \_gnd_net_\,
            in3 => \N__4087\,
            lcout => \U409_TICK.TICK603_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4051\,
            in2 => \N__4086\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_6_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3248\,
            in2 => \_gnd_net_\,
            in3 => \N__3237\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__5126\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3233\,
            in2 => \_gnd_net_\,
            in3 => \N__3222\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__5126\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3437\,
            in2 => \_gnd_net_\,
            in3 => \N__3420\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3416\,
            in2 => \_gnd_net_\,
            in3 => \N__3405\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__5126\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3401\,
            in3 => \N__3378\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4019\,
            in2 => \_gnd_net_\,
            in3 => \N__3375\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__5126\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3371\,
            in2 => \_gnd_net_\,
            in3 => \N__3351\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3347\,
            in2 => \_gnd_net_\,
            in3 => \N__3330\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_10_7_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4007\,
            in2 => \_gnd_net_\,
            in3 => \N__3327\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__5130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3320\,
            in2 => \_gnd_net_\,
            in3 => \N__3309\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__5130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3305\,
            in2 => \_gnd_net_\,
            in3 => \N__3291\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__5130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4034\,
            in2 => \_gnd_net_\,
            in3 => \N__3519\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__5130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3515\,
            in2 => \_gnd_net_\,
            in3 => \N__3498\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3872\,
            in2 => \_gnd_net_\,
            in3 => \N__3495\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3488\,
            in2 => \_gnd_net_\,
            in3 => \N__3492\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__4200\,
            in1 => \N__4183\,
            in2 => \N__4141\,
            in3 => \N__4166\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__3456\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4276\,
            in1 => \N__4720\,
            in2 => \_gnd_net_\,
            in3 => \N__4771\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4682\,
            in2 => \N__3444\,
            in3 => \N__4256\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__5334\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__3653\,
            in1 => \N__4784\,
            in2 => \N__3699\,
            in3 => \N__4621\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4287\,
            in2 => \N__3441\,
            in3 => \N__4746\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__5334\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001110101"
        )
    port map (
            in0 => \N__4623\,
            in1 => \N__3695\,
            in2 => \N__3652\,
            in3 => \N__4657\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5327\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__3558\,
            in1 => \N__4622\,
            in2 => \_gnd_net_\,
            in3 => \N__4785\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5327\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4277\,
            in1 => \N__4772\,
            in2 => \_gnd_net_\,
            in3 => \N__4257\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5327\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__4658\,
            in1 => \N__4583\,
            in2 => \_gnd_net_\,
            in3 => \N__4608\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5327\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__4725\,
            in1 => \N__4773\,
            in2 => \N__4281\,
            in3 => \N__4258\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5327\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__4698\,
            in1 => \N__3564\,
            in2 => \N__4263\,
            in3 => \N__4683\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5327\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4551\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__3557\,
            in1 => \N__3545\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__3802\,
            in1 => \N__3814\,
            in2 => \N__3534\,
            in3 => \N__3530\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001001100"
        )
    port map (
            in0 => \N__5467\,
            in1 => \N__3827\,
            in2 => \N__3849\,
            in3 => \N__3804\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__3803\,
            in1 => \N__3815\,
            in2 => \_gnd_net_\,
            in3 => \N__5466\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__3816\,
            in1 => \_gnd_net_\,
            in2 => \N__5485\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__4448\,
            in1 => \N__4524\,
            in2 => \N__3792\,
            in3 => \N__4409\,
            lcout => \nBUFEN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4104\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3780\,
            lcout => \U409_ADDRESS_DECODE_un1_nCIACS1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4103\,
            in2 => \_gnd_net_\,
            in3 => \N__3738\,
            lcout => \U409_ADDRESS_DECODE_un1_nCIACS0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__3951\,
            in1 => \N__3921\,
            in2 => \N__4092\,
            in3 => \N__3987\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5171\,
            in1 => \N__5273\,
            in2 => \N__5235\,
            in3 => \N__4854\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__4956\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4937\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4914\,
            in1 => \N__4803\,
            in2 => \N__4992\,
            in3 => \N__4955\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5274\,
            in1 => \N__5173\,
            in2 => \N__5229\,
            in3 => \N__4830\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4091\,
            in2 => \_gnd_net_\,
            in3 => \N__4055\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__5272\,
            in1 => \N__5172\,
            in2 => \N__5228\,
            in3 => \N__4936\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__4035\,
            in1 => \N__3873\,
            in2 => \N__4023\,
            in3 => \N__4008\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => \U409_TICK.TICK603_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3954\,
            in1 => \N__3919\,
            in2 => \N__3882\,
            in3 => \N__3879\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5177\,
            in1 => \N__5269\,
            in2 => \N__5227\,
            in3 => \N__5046\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4866\,
            in1 => \N__4896\,
            in2 => \_gnd_net_\,
            in3 => \N__4935\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3861\,
            in1 => \N__5037\,
            in2 => \N__3852\,
            in3 => \N__5076\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__5271\,
            in1 => \N__5207\,
            in2 => \N__4236\,
            in3 => \N__4217\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5019\,
            in1 => \N__4881\,
            in2 => \N__4821\,
            in3 => \N__4968\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5295\,
            in1 => \N__5142\,
            in2 => \N__5061\,
            in3 => \N__4844\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5270\,
            in1 => \N__5178\,
            in2 => \N__4206\,
            in3 => \N__5007\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__5603\,
            in1 => \N__5648\,
            in2 => \_gnd_net_\,
            in3 => \N__5682\,
            lcout => OPEN,
            ltout => \U409_CIA.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__4161\,
            in1 => \N__5604\,
            in2 => \N__4203\,
            in3 => \N__4344\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_HOLD_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__4184\,
            in1 => \N__4162\,
            in2 => \N__4146\,
            in3 => \N__4198\,
            lcout => \U409_CIA.CIA_HOLDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__4199\,
            in1 => \N__4185\,
            in2 => \N__4167\,
            in3 => \N__4145\,
            lcout => \CIA_ENABLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5645\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5697\,
            in1 => \N__5718\,
            in2 => \_gnd_net_\,
            in3 => \N__5739\,
            lcout => \U409_CIA.CLKCIA8_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5647\,
            in2 => \_gnd_net_\,
            in3 => \N__5680\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_1_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5698\,
            in1 => \N__5602\,
            in2 => \N__5745\,
            in3 => \N__5719\,
            lcout => \U409_CIA.CLKCIA6_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_2_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5601\,
            in1 => \N__5644\,
            in2 => \_gnd_net_\,
            in3 => \N__5679\,
            lcout => OPEN,
            ltout => \U409_CIA.N_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_0_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4300\,
            in2 => \N__4347\,
            in3 => \N__4343\,
            lcout => OPEN,
            ltout => \U409_CIA.CLKCIAZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__4332\,
            in1 => \N__5646\,
            in2 => \N__4326\,
            in3 => \N__5681\,
            lcout => \CLKCIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4656\,
            in1 => \N__4582\,
            in2 => \_gnd_net_\,
            in3 => \N__4607\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4605\,
            in1 => \N__4745\,
            in2 => \N__4584\,
            in3 => \N__4654\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4606\,
            in1 => \N__4655\,
            in2 => \_gnd_net_\,
            in3 => \N__4262\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__5326\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4680\,
            in1 => \N__4744\,
            in2 => \N__4659\,
            in3 => \N__4696\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4770\,
            in1 => \N__4719\,
            in2 => \N__4788\,
            in3 => \N__4559\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4769\,
            in1 => \N__4743\,
            in2 => \N__4724\,
            in3 => \N__4697\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4681\,
            in1 => \N__4653\,
            in2 => \N__4626\,
            in3 => \N__4560\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4604\,
            in2 => \_gnd_net_\,
            in3 => \N__4578\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5403\,
            in2 => \_gnd_net_\,
            in3 => \N__4550\,
            lcout => \TACK_EN_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            ce => \N__4539\,
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__4525\,
            in1 => \N__4447\,
            in2 => \_gnd_net_\,
            in3 => \N__4410\,
            lcout => \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4949\,
            in2 => \N__4938\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4910\,
            in2 => \_gnd_net_\,
            in3 => \N__4899\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4895\,
            in2 => \_gnd_net_\,
            in3 => \N__4884\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4880\,
            in2 => \_gnd_net_\,
            in3 => \N__4869\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4865\,
            in2 => \_gnd_net_\,
            in3 => \N__4848\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4845\,
            in3 => \N__4824\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4817\,
            in2 => \_gnd_net_\,
            in3 => \N__4806\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4802\,
            in2 => \_gnd_net_\,
            in3 => \N__4791\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5141\,
            in2 => \_gnd_net_\,
            in3 => \N__5079\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_7_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5075\,
            in2 => \_gnd_net_\,
            in3 => \N__5064\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__5125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5057\,
            in2 => \_gnd_net_\,
            in3 => \N__5040\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5036\,
            in2 => \_gnd_net_\,
            in3 => \N__5025\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__5125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5288\,
            in2 => \_gnd_net_\,
            in3 => \N__5022\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5018\,
            in2 => \_gnd_net_\,
            in3 => \N__5001\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4967\,
            in2 => \_gnd_net_\,
            in3 => \N__4998\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4991\,
            in2 => \_gnd_net_\,
            in3 => \N__4995\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__5174\,
            in1 => \N__5276\,
            in2 => \N__4977\,
            in3 => \N__5223\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5275\,
            in1 => \N__5175\,
            in2 => \N__5230\,
            in3 => \N__5301\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__5277\,
            in1 => \N__5241\,
            in2 => \N__5231\,
            in3 => \N__5176\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5677\,
            in2 => \N__5649\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5740\,
            in2 => \_gnd_net_\,
            in3 => \N__5094\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__5572\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5598\,
            in2 => \_gnd_net_\,
            in3 => \N__5091\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5699\,
            in2 => \_gnd_net_\,
            in3 => \N__5088\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__5572\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5720\,
            in2 => \_gnd_net_\,
            in3 => \N__5085\,
            lcout => OPEN,
            ltout => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__5600\,
            in1 => \N__5642\,
            in2 => \N__5082\,
            in3 => \N__5655\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5572\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5741\,
            in1 => \N__5721\,
            in2 => \N__5703\,
            in3 => \N__5678\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\,
            ltout => \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010110101010"
        )
    port map (
            in0 => \N__5599\,
            in1 => \N__5643\,
            in2 => \N__5613\,
            in3 => \N__5610\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5572\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_iobuf_RNO_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5559\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_353_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__5532\,
            in1 => \N__5504\,
            in2 => \_gnd_net_\,
            in3 => \N__5410\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 14 2024 11:09:01

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U111_TOP" view "INTERFACE"

module U111_TOP (
    D_LL_AMIGA,
    D_LM_AMIGA,
    D_UU_AMIGA,
    D_UM_AMIGA,
    D_UU_040,
    D_LL_040,
    D_LM_040,
    D_UM_040,
    A_AMIGA,
    A_040,
    SIZ,
    TSn,
    RESETn,
    CLKRAMA,
    PORTSIZE,
    CLK40B,
    TBI_CPUn,
    TAn,
    CPUBGn,
    BUFENn,
    RnW,
    CLK80_CPU,
    BUFDIR,
    TCI_CPUn,
    TS_CPUn,
    CLKRAMB,
    CLK40A,
    DMAn,
    CLK40C,
    CLK40_IN,
    TACKn,
    BGn);

    inout [7:0] D_LL_AMIGA;
    inout [7:0] D_LM_AMIGA;
    inout [7:0] D_UU_AMIGA;
    inout [7:0] D_UM_AMIGA;
    inout [7:0] D_UU_040;
    inout [7:0] D_LL_040;
    inout [7:0] D_LM_040;
    inout [7:0] D_UM_040;
    output [1:0] A_AMIGA;
    input [1:0] A_040;
    input [1:0] SIZ;
    output TSn;
    input RESETn;
    output CLKRAMA;
    input PORTSIZE;
    output CLK40B;
    output TBI_CPUn;
    output TAn;
    output CPUBGn;
    output BUFENn;
    input RnW;
    output CLK80_CPU;
    output BUFDIR;
    output TCI_CPUn;
    input TS_CPUn;
    output CLKRAMB;
    output CLK40A;
    output DMAn;
    output CLK40C;
    input CLK40_IN;
    input TACKn;
    input BGn;

    wire N__7858;
    wire N__7842;
    wire N__7841;
    wire N__7840;
    wire N__7833;
    wire N__7832;
    wire N__7831;
    wire N__7824;
    wire N__7823;
    wire N__7822;
    wire N__7815;
    wire N__7814;
    wire N__7813;
    wire N__7806;
    wire N__7805;
    wire N__7804;
    wire N__7797;
    wire N__7796;
    wire N__7795;
    wire N__7788;
    wire N__7787;
    wire N__7786;
    wire N__7779;
    wire N__7778;
    wire N__7777;
    wire N__7770;
    wire N__7769;
    wire N__7768;
    wire N__7761;
    wire N__7760;
    wire N__7759;
    wire N__7752;
    wire N__7751;
    wire N__7750;
    wire N__7743;
    wire N__7742;
    wire N__7741;
    wire N__7734;
    wire N__7733;
    wire N__7732;
    wire N__7725;
    wire N__7724;
    wire N__7723;
    wire N__7716;
    wire N__7715;
    wire N__7714;
    wire N__7707;
    wire N__7706;
    wire N__7705;
    wire N__7698;
    wire N__7697;
    wire N__7696;
    wire N__7689;
    wire N__7688;
    wire N__7687;
    wire N__7680;
    wire N__7679;
    wire N__7678;
    wire N__7671;
    wire N__7670;
    wire N__7669;
    wire N__7662;
    wire N__7661;
    wire N__7660;
    wire N__7653;
    wire N__7652;
    wire N__7651;
    wire N__7644;
    wire N__7643;
    wire N__7642;
    wire N__7635;
    wire N__7634;
    wire N__7633;
    wire N__7626;
    wire N__7625;
    wire N__7624;
    wire N__7617;
    wire N__7616;
    wire N__7615;
    wire N__7608;
    wire N__7607;
    wire N__7606;
    wire N__7599;
    wire N__7598;
    wire N__7597;
    wire N__7590;
    wire N__7589;
    wire N__7588;
    wire N__7581;
    wire N__7580;
    wire N__7579;
    wire N__7572;
    wire N__7571;
    wire N__7570;
    wire N__7563;
    wire N__7562;
    wire N__7561;
    wire N__7554;
    wire N__7553;
    wire N__7552;
    wire N__7545;
    wire N__7544;
    wire N__7543;
    wire N__7536;
    wire N__7535;
    wire N__7534;
    wire N__7527;
    wire N__7526;
    wire N__7525;
    wire N__7518;
    wire N__7517;
    wire N__7516;
    wire N__7509;
    wire N__7508;
    wire N__7507;
    wire N__7500;
    wire N__7499;
    wire N__7498;
    wire N__7491;
    wire N__7490;
    wire N__7489;
    wire N__7482;
    wire N__7481;
    wire N__7480;
    wire N__7473;
    wire N__7472;
    wire N__7471;
    wire N__7464;
    wire N__7463;
    wire N__7462;
    wire N__7455;
    wire N__7454;
    wire N__7453;
    wire N__7446;
    wire N__7445;
    wire N__7444;
    wire N__7437;
    wire N__7436;
    wire N__7435;
    wire N__7428;
    wire N__7427;
    wire N__7426;
    wire N__7419;
    wire N__7418;
    wire N__7417;
    wire N__7410;
    wire N__7409;
    wire N__7408;
    wire N__7401;
    wire N__7400;
    wire N__7399;
    wire N__7392;
    wire N__7391;
    wire N__7390;
    wire N__7383;
    wire N__7382;
    wire N__7381;
    wire N__7374;
    wire N__7373;
    wire N__7372;
    wire N__7365;
    wire N__7364;
    wire N__7363;
    wire N__7356;
    wire N__7355;
    wire N__7354;
    wire N__7347;
    wire N__7346;
    wire N__7345;
    wire N__7338;
    wire N__7337;
    wire N__7336;
    wire N__7329;
    wire N__7328;
    wire N__7327;
    wire N__7320;
    wire N__7319;
    wire N__7318;
    wire N__7311;
    wire N__7310;
    wire N__7309;
    wire N__7302;
    wire N__7301;
    wire N__7300;
    wire N__7293;
    wire N__7292;
    wire N__7291;
    wire N__7284;
    wire N__7283;
    wire N__7282;
    wire N__7275;
    wire N__7274;
    wire N__7273;
    wire N__7266;
    wire N__7265;
    wire N__7264;
    wire N__7257;
    wire N__7256;
    wire N__7255;
    wire N__7248;
    wire N__7247;
    wire N__7246;
    wire N__7239;
    wire N__7238;
    wire N__7237;
    wire N__7230;
    wire N__7229;
    wire N__7228;
    wire N__7221;
    wire N__7220;
    wire N__7219;
    wire N__7212;
    wire N__7211;
    wire N__7210;
    wire N__7203;
    wire N__7202;
    wire N__7201;
    wire N__7194;
    wire N__7193;
    wire N__7192;
    wire N__7185;
    wire N__7184;
    wire N__7183;
    wire N__7176;
    wire N__7175;
    wire N__7174;
    wire N__7167;
    wire N__7166;
    wire N__7165;
    wire N__7158;
    wire N__7157;
    wire N__7156;
    wire N__7149;
    wire N__7148;
    wire N__7147;
    wire N__7140;
    wire N__7139;
    wire N__7138;
    wire N__7131;
    wire N__7130;
    wire N__7129;
    wire N__7122;
    wire N__7121;
    wire N__7120;
    wire N__7113;
    wire N__7112;
    wire N__7111;
    wire N__7104;
    wire N__7103;
    wire N__7102;
    wire N__7095;
    wire N__7094;
    wire N__7093;
    wire N__7086;
    wire N__7085;
    wire N__7084;
    wire N__7077;
    wire N__7076;
    wire N__7075;
    wire N__7068;
    wire N__7067;
    wire N__7066;
    wire N__7059;
    wire N__7058;
    wire N__7057;
    wire N__7050;
    wire N__7049;
    wire N__7048;
    wire N__7031;
    wire N__7030;
    wire N__7027;
    wire N__7024;
    wire N__7023;
    wire N__7020;
    wire N__7017;
    wire N__7014;
    wire N__7011;
    wire N__7008;
    wire N__7005;
    wire N__7002;
    wire N__6999;
    wire N__6996;
    wire N__6993;
    wire N__6990;
    wire N__6987;
    wire N__6984;
    wire N__6979;
    wire N__6974;
    wire N__6971;
    wire N__6970;
    wire N__6969;
    wire N__6968;
    wire N__6967;
    wire N__6966;
    wire N__6965;
    wire N__6964;
    wire N__6963;
    wire N__6960;
    wire N__6959;
    wire N__6938;
    wire N__6935;
    wire N__6932;
    wire N__6929;
    wire N__6928;
    wire N__6927;
    wire N__6924;
    wire N__6921;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6904;
    wire N__6901;
    wire N__6898;
    wire N__6895;
    wire N__6892;
    wire N__6889;
    wire N__6886;
    wire N__6883;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6871;
    wire N__6868;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6856;
    wire N__6853;
    wire N__6850;
    wire N__6847;
    wire N__6844;
    wire N__6841;
    wire N__6838;
    wire N__6835;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6800;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6787;
    wire N__6784;
    wire N__6781;
    wire N__6778;
    wire N__6775;
    wire N__6772;
    wire N__6769;
    wire N__6766;
    wire N__6763;
    wire N__6760;
    wire N__6757;
    wire N__6752;
    wire N__6749;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6710;
    wire N__6707;
    wire N__6704;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6694;
    wire N__6691;
    wire N__6688;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6676;
    wire N__6673;
    wire N__6670;
    wire N__6667;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6641;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6616;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6599;
    wire N__6596;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6584;
    wire N__6581;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6529;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6500;
    wire N__6497;
    wire N__6494;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6467;
    wire N__6464;
    wire N__6461;
    wire N__6458;
    wire N__6455;
    wire N__6452;
    wire N__6449;
    wire N__6446;
    wire N__6443;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6419;
    wire N__6416;
    wire N__6413;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6380;
    wire N__6377;
    wire N__6374;
    wire N__6371;
    wire N__6368;
    wire N__6367;
    wire N__6366;
    wire N__6365;
    wire N__6364;
    wire N__6363;
    wire N__6362;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6350;
    wire N__6347;
    wire N__6342;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6330;
    wire N__6329;
    wire N__6328;
    wire N__6327;
    wire N__6326;
    wire N__6321;
    wire N__6318;
    wire N__6317;
    wire N__6316;
    wire N__6315;
    wire N__6314;
    wire N__6311;
    wire N__6306;
    wire N__6303;
    wire N__6300;
    wire N__6299;
    wire N__6298;
    wire N__6297;
    wire N__6294;
    wire N__6291;
    wire N__6290;
    wire N__6289;
    wire N__6284;
    wire N__6281;
    wire N__6280;
    wire N__6279;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6269;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6249;
    wire N__6248;
    wire N__6247;
    wire N__6244;
    wire N__6241;
    wire N__6238;
    wire N__6235;
    wire N__6234;
    wire N__6233;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6223;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6179;
    wire N__6174;
    wire N__6171;
    wire N__6170;
    wire N__6165;
    wire N__6160;
    wire N__6157;
    wire N__6152;
    wire N__6149;
    wire N__6144;
    wire N__6139;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6122;
    wire N__6115;
    wire N__6104;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6056;
    wire N__6053;
    wire N__6050;
    wire N__6047;
    wire N__6044;
    wire N__6041;
    wire N__6038;
    wire N__6035;
    wire N__6032;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__5998;
    wire N__5995;
    wire N__5992;
    wire N__5989;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5957;
    wire N__5954;
    wire N__5951;
    wire N__5948;
    wire N__5945;
    wire N__5942;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5927;
    wire N__5926;
    wire N__5925;
    wire N__5922;
    wire N__5919;
    wire N__5916;
    wire N__5913;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5897;
    wire N__5894;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5845;
    wire N__5842;
    wire N__5839;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5756;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5729;
    wire N__5726;
    wire N__5723;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5705;
    wire N__5702;
    wire N__5701;
    wire N__5698;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5665;
    wire N__5662;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5624;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5569;
    wire N__5566;
    wire N__5563;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5549;
    wire N__5546;
    wire N__5545;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5532;
    wire N__5529;
    wire N__5526;
    wire N__5523;
    wire N__5518;
    wire N__5513;
    wire N__5512;
    wire N__5507;
    wire N__5506;
    wire N__5505;
    wire N__5504;
    wire N__5503;
    wire N__5502;
    wire N__5501;
    wire N__5500;
    wire N__5497;
    wire N__5488;
    wire N__5487;
    wire N__5486;
    wire N__5485;
    wire N__5484;
    wire N__5481;
    wire N__5478;
    wire N__5477;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5456;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5444;
    wire N__5441;
    wire N__5440;
    wire N__5437;
    wire N__5430;
    wire N__5421;
    wire N__5418;
    wire N__5417;
    wire N__5416;
    wire N__5413;
    wire N__5410;
    wire N__5409;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5397;
    wire N__5394;
    wire N__5391;
    wire N__5386;
    wire N__5381;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5346;
    wire N__5343;
    wire N__5340;
    wire N__5337;
    wire N__5334;
    wire N__5329;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5281;
    wire N__5280;
    wire N__5279;
    wire N__5278;
    wire N__5277;
    wire N__5276;
    wire N__5275;
    wire N__5274;
    wire N__5273;
    wire N__5270;
    wire N__5265;
    wire N__5254;
    wire N__5249;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5233;
    wire N__5232;
    wire N__5231;
    wire N__5230;
    wire N__5227;
    wire N__5224;
    wire N__5221;
    wire N__5218;
    wire N__5215;
    wire N__5210;
    wire N__5205;
    wire N__5202;
    wire N__5195;
    wire N__5194;
    wire N__5193;
    wire N__5190;
    wire N__5189;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5179;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5162;
    wire N__5159;
    wire N__5154;
    wire N__5149;
    wire N__5144;
    wire N__5141;
    wire N__5140;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5130;
    wire N__5127;
    wire N__5124;
    wire N__5121;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5095;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5048;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5040;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5014;
    wire N__5011;
    wire N__5008;
    wire N__5005;
    wire N__5002;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4864;
    wire N__4861;
    wire N__4858;
    wire N__4855;
    wire N__4852;
    wire N__4849;
    wire N__4846;
    wire N__4843;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4798;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4783;
    wire N__4780;
    wire N__4777;
    wire N__4774;
    wire N__4771;
    wire N__4768;
    wire N__4765;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4753;
    wire N__4752;
    wire N__4749;
    wire N__4748;
    wire N__4747;
    wire N__4746;
    wire N__4743;
    wire N__4742;
    wire N__4739;
    wire N__4738;
    wire N__4735;
    wire N__4730;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4706;
    wire N__4703;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4669;
    wire N__4668;
    wire N__4667;
    wire N__4666;
    wire N__4661;
    wire N__4658;
    wire N__4653;
    wire N__4648;
    wire N__4645;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4615;
    wire N__4614;
    wire N__4613;
    wire N__4612;
    wire N__4609;
    wire N__4606;
    wire N__4605;
    wire N__4602;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4588;
    wire N__4583;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4564;
    wire N__4561;
    wire N__4558;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4539;
    wire N__4536;
    wire N__4531;
    wire N__4528;
    wire N__4525;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4488;
    wire N__4483;
    wire N__4480;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4445;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4423;
    wire N__4420;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4401;
    wire N__4398;
    wire N__4393;
    wire N__4390;
    wire N__4387;
    wire N__4384;
    wire N__4381;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4309;
    wire N__4306;
    wire N__4303;
    wire N__4300;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4183;
    wire N__4180;
    wire N__4177;
    wire N__4172;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4133;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4075;
    wire N__4072;
    wire N__4069;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4051;
    wire N__4048;
    wire N__4045;
    wire N__4040;
    wire N__4039;
    wire N__4036;
    wire N__4031;
    wire N__4028;
    wire N__4027;
    wire N__4024;
    wire N__4021;
    wire N__4020;
    wire N__4019;
    wire N__4014;
    wire N__4011;
    wire N__4008;
    wire N__4007;
    wire N__4006;
    wire N__4005;
    wire N__4004;
    wire N__4003;
    wire N__4002;
    wire N__4001;
    wire N__3994;
    wire N__3991;
    wire N__3988;
    wire N__3985;
    wire N__3982;
    wire N__3979;
    wire N__3978;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3970;
    wire N__3969;
    wire N__3956;
    wire N__3953;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3936;
    wire N__3935;
    wire N__3934;
    wire N__3933;
    wire N__3932;
    wire N__3931;
    wire N__3924;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3914;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3900;
    wire N__3897;
    wire N__3894;
    wire N__3891;
    wire N__3890;
    wire N__3889;
    wire N__3888;
    wire N__3887;
    wire N__3884;
    wire N__3881;
    wire N__3880;
    wire N__3877;
    wire N__3872;
    wire N__3871;
    wire N__3856;
    wire N__3853;
    wire N__3850;
    wire N__3847;
    wire N__3844;
    wire N__3839;
    wire N__3836;
    wire N__3835;
    wire N__3834;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3824;
    wire N__3813;
    wire N__3812;
    wire N__3809;
    wire N__3806;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3796;
    wire N__3793;
    wire N__3792;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3760;
    wire N__3755;
    wire N__3750;
    wire N__3745;
    wire N__3740;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3680;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3668;
    wire N__3665;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3631;
    wire N__3628;
    wire N__3625;
    wire N__3620;
    wire N__3617;
    wire N__3614;
    wire N__3611;
    wire N__3608;
    wire N__3607;
    wire N__3604;
    wire N__3601;
    wire N__3598;
    wire N__3593;
    wire N__3590;
    wire N__3587;
    wire N__3584;
    wire N__3581;
    wire N__3580;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3568;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3550;
    wire N__3547;
    wire N__3544;
    wire N__3541;
    wire N__3538;
    wire N__3535;
    wire N__3530;
    wire N__3527;
    wire N__3524;
    wire N__3521;
    wire N__3518;
    wire N__3515;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire N__3497;
    wire N__3494;
    wire N__3491;
    wire N__3490;
    wire N__3487;
    wire N__3484;
    wire N__3481;
    wire N__3478;
    wire N__3477;
    wire N__3472;
    wire N__3469;
    wire N__3464;
    wire N__3461;
    wire N__3458;
    wire N__3455;
    wire N__3452;
    wire N__3449;
    wire N__3446;
    wire N__3443;
    wire N__3440;
    wire N__3437;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3425;
    wire N__3422;
    wire N__3419;
    wire N__3416;
    wire N__3413;
    wire N__3412;
    wire N__3409;
    wire N__3406;
    wire N__3403;
    wire N__3402;
    wire N__3399;
    wire N__3396;
    wire N__3393;
    wire N__3390;
    wire N__3385;
    wire N__3382;
    wire N__3379;
    wire N__3374;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3362;
    wire N__3359;
    wire N__3356;
    wire N__3353;
    wire N__3350;
    wire N__3347;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3337;
    wire N__3336;
    wire N__3333;
    wire N__3330;
    wire N__3327;
    wire N__3324;
    wire N__3319;
    wire N__3316;
    wire N__3313;
    wire N__3310;
    wire N__3305;
    wire N__3302;
    wire N__3299;
    wire N__3296;
    wire N__3293;
    wire N__3290;
    wire N__3287;
    wire N__3284;
    wire N__3281;
    wire N__3278;
    wire N__3275;
    wire N__3272;
    wire N__3269;
    wire N__3266;
    wire N__3263;
    wire N__3260;
    wire N__3257;
    wire N__3254;
    wire N__3251;
    wire N__3248;
    wire N__3245;
    wire N__3242;
    wire N__3239;
    wire N__3236;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3224;
    wire N__3221;
    wire N__3218;
    wire N__3215;
    wire N__3212;
    wire N__3209;
    wire N__3206;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3188;
    wire N__3185;
    wire N__3182;
    wire N__3179;
    wire N__3176;
    wire N__3173;
    wire N__3170;
    wire N__3167;
    wire N__3166;
    wire N__3163;
    wire N__3160;
    wire N__3157;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3128;
    wire N__3125;
    wire N__3122;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3097;
    wire N__3094;
    wire N__3091;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3077;
    wire N__3074;
    wire N__3071;
    wire N__3068;
    wire N__3065;
    wire N__3062;
    wire N__3059;
    wire N__3056;
    wire N__3053;
    wire N__3050;
    wire N__3047;
    wire N__3044;
    wire N__3041;
    wire N__3038;
    wire N__3035;
    wire N__3032;
    wire N__3029;
    wire N__3026;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3011;
    wire N__3008;
    wire N__3005;
    wire N__3002;
    wire N__2999;
    wire N__2996;
    wire N__2993;
    wire N__2990;
    wire N__2987;
    wire N__2984;
    wire N__2981;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2968;
    wire N__2965;
    wire N__2962;
    wire N__2959;
    wire N__2956;
    wire N__2955;
    wire N__2952;
    wire N__2949;
    wire N__2946;
    wire N__2939;
    wire N__2936;
    wire N__2933;
    wire N__2930;
    wire N__2927;
    wire N__2924;
    wire N__2921;
    wire N__2918;
    wire N__2915;
    wire N__2912;
    wire N__2909;
    wire N__2906;
    wire N__2905;
    wire N__2902;
    wire N__2899;
    wire N__2896;
    wire N__2893;
    wire N__2890;
    wire N__2887;
    wire N__2884;
    wire N__2881;
    wire N__2878;
    wire N__2875;
    wire N__2872;
    wire N__2869;
    wire N__2866;
    wire N__2863;
    wire N__2858;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2839;
    wire N__2838;
    wire N__2837;
    wire N__2836;
    wire N__2835;
    wire N__2834;
    wire N__2833;
    wire N__2832;
    wire N__2829;
    wire N__2826;
    wire N__2823;
    wire N__2822;
    wire N__2821;
    wire N__2820;
    wire N__2819;
    wire N__2818;
    wire N__2815;
    wire N__2812;
    wire N__2809;
    wire N__2806;
    wire N__2803;
    wire N__2800;
    wire N__2797;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2785;
    wire N__2784;
    wire N__2783;
    wire N__2782;
    wire N__2781;
    wire N__2780;
    wire N__2779;
    wire N__2778;
    wire N__2775;
    wire N__2772;
    wire N__2769;
    wire N__2756;
    wire N__2747;
    wire N__2744;
    wire N__2741;
    wire N__2738;
    wire N__2735;
    wire N__2732;
    wire N__2729;
    wire N__2726;
    wire N__2723;
    wire N__2714;
    wire N__2713;
    wire N__2712;
    wire N__2711;
    wire N__2710;
    wire N__2699;
    wire N__2688;
    wire N__2685;
    wire N__2682;
    wire N__2679;
    wire N__2676;
    wire N__2675;
    wire N__2674;
    wire N__2673;
    wire N__2672;
    wire N__2671;
    wire N__2668;
    wire N__2657;
    wire N__2654;
    wire N__2651;
    wire N__2648;
    wire N__2645;
    wire N__2642;
    wire N__2639;
    wire N__2628;
    wire N__2625;
    wire N__2618;
    wire N__2617;
    wire N__2614;
    wire N__2611;
    wire N__2606;
    wire N__2603;
    wire N__2600;
    wire N__2597;
    wire N__2594;
    wire N__2591;
    wire N__2588;
    wire N__2585;
    wire N__2582;
    wire N__2579;
    wire N__2576;
    wire N__2573;
    wire N__2570;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2558;
    wire N__2555;
    wire N__2552;
    wire N__2549;
    wire N__2546;
    wire N__2543;
    wire N__2540;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2516;
    wire N__2513;
    wire N__2510;
    wire N__2507;
    wire N__2504;
    wire N__2501;
    wire N__2498;
    wire N__2495;
    wire N__2492;
    wire N__2489;
    wire N__2486;
    wire N__2483;
    wire N__2480;
    wire N__2477;
    wire N__2474;
    wire N__2471;
    wire N__2468;
    wire N__2465;
    wire N__2462;
    wire N__2461;
    wire N__2458;
    wire N__2455;
    wire N__2452;
    wire N__2449;
    wire N__2446;
    wire N__2443;
    wire N__2440;
    wire N__2437;
    wire N__2434;
    wire N__2431;
    wire N__2426;
    wire N__2423;
    wire N__2420;
    wire N__2417;
    wire N__2414;
    wire N__2411;
    wire N__2408;
    wire N__2405;
    wire N__2402;
    wire N__2399;
    wire N__2396;
    wire N__2393;
    wire N__2390;
    wire N__2387;
    wire N__2384;
    wire N__2381;
    wire N__2378;
    wire N__2375;
    wire N__2372;
    wire N__2369;
    wire N__2366;
    wire N__2363;
    wire N__2360;
    wire N__2357;
    wire N__2354;
    wire N__2351;
    wire N__2348;
    wire N__2345;
    wire N__2342;
    wire N__2339;
    wire N__2336;
    wire N__2333;
    wire N__2330;
    wire N__2327;
    wire N__2324;
    wire N__2321;
    wire N__2318;
    wire N__2315;
    wire N__2312;
    wire N__2309;
    wire N__2306;
    wire N__2303;
    wire N__2300;
    wire N__2297;
    wire N__2294;
    wire N__2291;
    wire N__2288;
    wire N__2285;
    wire N__2282;
    wire N__2279;
    wire N__2276;
    wire N__2273;
    wire N__2270;
    wire N__2267;
    wire N__2264;
    wire N__2261;
    wire N__2258;
    wire N__2255;
    wire N__2252;
    wire N__2249;
    wire N__2246;
    wire N__2243;
    wire N__2240;
    wire N__2237;
    wire N__2234;
    wire N__2231;
    wire N__2228;
    wire N__2225;
    wire N__2222;
    wire N__2219;
    wire N__2216;
    wire N__2213;
    wire N__2210;
    wire N__2207;
    wire N__2204;
    wire N__2201;
    wire N__2198;
    wire VCCG0;
    wire GNDG0;
    wire A_040_c_1;
    wire A_040_c_0;
    wire A_AMIGA_c_0;
    wire D_LL_AMIGA_in_2;
    wire un1_D_LL_AMIGA_2;
    wire D_LM_AMIGA_in_2;
    wire un1_D_LM_AMIGA_2;
    wire D_UM_040_in_1;
    wire D_LL_040_in_1;
    wire un1_D_UM_040_1;
    wire RnW_c_i_0;
    wire D_LM_AMIGA_in_4;
    wire un1_D_LM_AMIGA_4;
    wire D_LM_AMIGA_in_5;
    wire un1_D_LM_AMIGA_5;
    wire D_LM_AMIGA_in_6;
    wire un1_D_LM_AMIGA_6;
    wire D_UU_040_in_3;
    wire D_LM_040_in_3;
    wire un1_D_UU_040_3;
    wire D_LL_AMIGA_in_0;
    wire un1_D_LL_AMIGA_0;
    wire D_LL_AMIGA_in_1;
    wire un1_D_LL_AMIGA_1;
    wire D_LM_AMIGA_in_3;
    wire un1_D_LM_AMIGA_3;
    wire D_LM_AMIGA_in_7;
    wire un1_D_LM_AMIGA_7;
    wire A_AMIGA_c_1;
    wire D_UM_040_in_7;
    wire D_LL_040_in_7;
    wire un1_D_UM_040_7;
    wire D_LM_040_in_6;
    wire D_UU_040_in_6;
    wire un1_D_UU_040_6;
    wire D_LL_AMIGA_in_3;
    wire un1_D_LL_AMIGA_3;
    wire un1_D_UM_AMIGA_0;
    wire D_UM_AMIGA_in_0;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net ;
    wire \INVU111_CYCLE_SM.TA_EN_nessC_net ;
    wire \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net ;
    wire D_LM_040_in_1;
    wire D_UU_040_in_1;
    wire un1_D_UU_040_1;
    wire D_UU_AMIGA_in_6;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ;
    wire un1_D_UU_AMIGA_6;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ;
    wire D_UU_AMIGA_in_4;
    wire un1_D_UU_AMIGA_4;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ;
    wire D_UU_AMIGA_in_7;
    wire un1_D_UU_AMIGA_7;
    wire D_LL_AMIGA_in_4;
    wire un1_D_LL_AMIGA_4;
    wire D_LM_AMIGA_in_0;
    wire un1_D_LM_AMIGA_0;
    wire D_LM_AMIGA_in_1;
    wire un1_D_LM_AMIGA_1;
    wire \INVU111_CYCLE_SM.TSnC_net ;
    wire \U111_CYCLE_SM.A_OUTZ0 ;
    wire \U111_CYCLE_SM.LW_CYCLE_r_1_cascade_ ;
    wire \U111_CYCLE_SM.un1_CYCLE_STATE_1_0 ;
    wire \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_cascade_ ;
    wire RESETn_c_i;
    wire \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_0 ;
    wire \U111_CYCLE_SM.TS_EN10 ;
    wire \U111_CYCLE_SM.TS_ENZ0 ;
    wire TSn_c;
    wire \U111_CYCLE_SM.LW_CYCLE_STARTZ0 ;
    wire \INVU111_CYCLE_SM.A_OUTC_net ;
    wire \INVU111_CYCLE_SM.CYCLE_STATE_0C_net ;
    wire RnW_c;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa ;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net ;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ;
    wire D_UM_AMIGA_in_1;
    wire un1_D_UM_AMIGA_1;
    wire D_UU_AMIGA_in_1;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ;
    wire un1_D_UU_AMIGA_1;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ;
    wire D_UM_AMIGA_in_4;
    wire un1_D_UM_AMIGA_4;
    wire D_UU_040_in_0;
    wire D_LM_040_in_0;
    wire un1_D_UU_040_0;
    wire D_UU_040_in_2;
    wire D_LM_040_in_2;
    wire un1_D_UU_040_2;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ;
    wire D_UU_AMIGA_in_0;
    wire un1_D_UU_AMIGA_0;
    wire D_LL_AMIGA_in_6;
    wire un1_D_LL_AMIGA_6;
    wire D_LL_AMIGA_in_5;
    wire un1_D_LL_AMIGA_5;
    wire D_LL_AMIGA_in_7;
    wire un1_D_LL_AMIGA_7;
    wire D_UM_040_in_2;
    wire D_LL_040_in_2;
    wire un1_D_UM_040_2;
    wire un1_D_UM_AMIGA_2;
    wire D_UM_AMIGA_in_2;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net ;
    wire RESETn_c;
    wire \INVU111_CYCLE_SM.CYCLE_STATE_1C_net ;
    wire \U111_CYCLE_SM.TA_ENZ0 ;
    wire TACKn_c;
    wire TAn_0_i;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ;
    wire TS_CPUn_c;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ;
    wire \U111_CYCLE_SM.TS_EN_4 ;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ;
    wire \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0 ;
    wire D_UM_AMIGA_in_3;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ;
    wire un1_D_UM_AMIGA_3;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ;
    wire D_UM_AMIGA_in_7;
    wire un1_D_UM_AMIGA_7;
    wire D_LL_040_in_4;
    wire D_UM_040_in_4;
    wire un1_D_UM_040_4;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ;
    wire D_UU_AMIGA_in_3;
    wire un1_D_UU_AMIGA_3;
    wire D_UM_040_in_5;
    wire D_LL_040_in_5;
    wire un1_D_UM_040_5;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ;
    wire D_UU_AMIGA_in_5;
    wire un1_D_UU_AMIGA_5;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ;
    wire D_UU_AMIGA_in_2;
    wire un1_D_UU_AMIGA_2;
    wire D_UM_AMIGA_in_5;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ;
    wire un1_D_UM_AMIGA_5;
    wire CLK40;
    wire GB_BUFFER_CLK40_THRU_CO;
    wire \U111_CYCLE_SM.LW_CYCLEZ0 ;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ;
    wire D_UM_AMIGA_in_6;
    wire un1_D_UM_AMIGA_6;
    wire CLK80;
    wire GB_BUFFER_CLK80_THRU_CO;
    wire D_LM_040_in_5;
    wire D_UU_040_in_5;
    wire un1_D_UU_040_5;
    wire D_LM_040_in_7;
    wire D_UU_040_in_7;
    wire un1_D_UU_040_7;
    wire D_UM_040_in_0;
    wire D_LL_040_in_0;
    wire un1_D_UM_040_0;
    wire D_LL_040_in_6;
    wire D_UM_040_in_6;
    wire un1_D_UM_040_6;
    wire D_LL_040_in_3;
    wire D_UM_040_in_3;
    wire un1_D_UM_040_3;
    wire SIZ_c_0;
    wire SIZ_c_1;
    wire PORTSIZE_c;
    wire \U111_CYCLE_SM.LW_TRANS_0 ;
    wire D_UU_040_in_4;
    wire \U111_CYCLE_SM.FLIP ;
    wire D_LM_040_in_4;
    wire un1_D_UU_040_4;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    defparam pll_pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll_pll.TEST_MODE=1'b0;
    defparam pll_pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll_pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll_pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll_pll.FILTER_RANGE=3'b011;
    defparam pll_pll.FEEDBACK_PATH="SIMPLE";
    defparam pll_pll.FDA_RELATIVE=4'b0000;
    defparam pll_pll.FDA_FEEDBACK=4'b0000;
    defparam pll_pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll_pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll_pll.DIVR=4'b0000;
    defparam pll_pll.DIVQ=3'b011;
    defparam pll_pll.DIVF=7'b0001111;
    defparam pll_pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40_2F pll_pll (
            .SCLK(),
            .PLLOUTGLOBALA(CLK80),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALB(CLK40),
            .SDI(),
            .PLLOUTCOREA(),
            .BYPASS(),
            .RESETB(N__7030),
            .PLLOUTCOREB(),
            .LOCK(),
            .SDO(),
            .EXTFEEDBACK(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__7858));
    IO_PAD pll_iopad (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__7858),
            .PACKAGEPIN(CLK40_IN));
    defparam D_UM_040_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_3_iopad (
            .OE(N__7842),
            .DIN(N__7841),
            .DOUT(N__7840),
            .PACKAGEPIN(D_UM_040[3]));
    defparam D_UM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_3_preio (
            .PADOEN(N__7842),
            .PADOUT(N__7841),
            .PADIN(N__7840),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3889),
            .DIN0(D_UM_040_in_3),
            .DOUT0(N__5078),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_1_iopad (
            .OE(N__7833),
            .DIN(N__7832),
            .DOUT(N__7831),
            .PACKAGEPIN(D_LL_AMIGA[1]));
    defparam D_LL_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_1_preio (
            .PADOEN(N__7833),
            .PADOUT(N__7832),
            .PADIN(N__7831),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2822),
            .DIN0(D_LL_AMIGA_in_1),
            .DOUT0(N__2905),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_5_iopad (
            .OE(N__7824),
            .DIN(N__7823),
            .DOUT(N__7822),
            .PACKAGEPIN(D_UU_AMIGA[5]));
    defparam D_UU_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_5_preio (
            .PADOEN(N__7824),
            .PADOUT(N__7823),
            .PADIN(N__7822),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2819),
            .DIN0(D_UU_AMIGA_in_5),
            .DOUT0(N__6809),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_ibuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_ibuf_iopad (
            .OE(N__7815),
            .DIN(N__7814),
            .DOUT(N__7813),
            .PACKAGEPIN(TACKn));
    defparam TACKn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TACKn_ibuf_preio (
            .PADOEN(N__7815),
            .PADOUT(N__7814),
            .PADIN(N__7813),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TACKn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_6_iopad (
            .OE(N__7806),
            .DIN(N__7805),
            .DOUT(N__7804),
            .PACKAGEPIN(D_UU_040[6]));
    defparam D_UU_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_6_preio (
            .PADOEN(N__7806),
            .PADOUT(N__7805),
            .PADIN(N__7804),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3936),
            .DIN0(D_UU_040_in_6),
            .DOUT0(N__3449),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam CPUBGn_obuf_iopad.PULLUP=1'b1;
    IO_PAD CPUBGn_obuf_iopad (
            .OE(N__7797),
            .DIN(N__7796),
            .DOUT(N__7795),
            .PACKAGEPIN(CPUBGn));
    defparam CPUBGn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUBGn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CPUBGn_obuf_preio (
            .PADOEN(N__7797),
            .PADOUT(N__7796),
            .PADIN(N__7795),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_7_iopad (
            .OE(N__7788),
            .DIN(N__7787),
            .DOUT(N__7786),
            .PACKAGEPIN(D_LL_040[7]));
    defparam D_LL_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_7_preio (
            .PADOEN(N__7788),
            .PADOUT(N__7787),
            .PADIN(N__7786),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4003),
            .DIN0(D_LL_040_in_7),
            .DOUT0(N__4916),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_4_iopad (
            .OE(N__7779),
            .DIN(N__7778),
            .DOUT(N__7777),
            .PACKAGEPIN(D_LL_AMIGA[4]));
    defparam D_LL_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_4_preio (
            .PADOEN(N__7779),
            .PADOUT(N__7778),
            .PADIN(N__7777),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2821),
            .DIN0(D_LL_AMIGA_in_4),
            .DOUT0(N__6031),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_3_iopad (
            .OE(N__7770),
            .DIN(N__7769),
            .DOUT(N__7768),
            .PACKAGEPIN(D_UM_AMIGA[3]));
    defparam D_UM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_3_preio (
            .PADOEN(N__7770),
            .PADOUT(N__7769),
            .PADIN(N__7768),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2779),
            .DIN0(D_UM_AMIGA_in_3),
            .DOUT0(N__6503),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_3_iopad (
            .OE(N__7761),
            .DIN(N__7760),
            .DOUT(N__7759),
            .PACKAGEPIN(D_UU_040[3]));
    defparam D_UU_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_3_preio (
            .PADOEN(N__7761),
            .PADOUT(N__7760),
            .PADIN(N__7759),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3931),
            .DIN0(D_UU_040_in_3),
            .DOUT0(N__5894),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_1_iopad (
            .OE(N__7752),
            .DIN(N__7751),
            .DOUT(N__7750),
            .PACKAGEPIN(A_040[1]));
    defparam A_040_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_1_preio (
            .PADOEN(N__7752),
            .PADOUT(N__7751),
            .PADIN(N__7750),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_3_iopad (
            .OE(N__7743),
            .DIN(N__7742),
            .DOUT(N__7741),
            .PACKAGEPIN(D_LM_AMIGA[3]));
    defparam D_LM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_3_preio (
            .PADOEN(N__7743),
            .PADOUT(N__7742),
            .PADIN(N__7741),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2617),
            .DIN0(D_LM_AMIGA_in_3),
            .DOUT0(N__2471),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_0_iopad (
            .OE(N__7734),
            .DIN(N__7733),
            .DOUT(N__7732),
            .PACKAGEPIN(D_LM_040[0]));
    defparam D_LM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_0_preio (
            .PADOEN(N__7734),
            .PADOUT(N__7733),
            .PADIN(N__7732),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4004),
            .DIN0(D_LM_040_in_0),
            .DOUT0(N__3704),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_6_iopad (
            .OE(N__7725),
            .DIN(N__7724),
            .DOUT(N__7723),
            .PACKAGEPIN(D_UM_AMIGA[6]));
    defparam D_UM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_6_preio (
            .PADOEN(N__7725),
            .PADOUT(N__7724),
            .PADIN(N__7723),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2818),
            .DIN0(D_UM_AMIGA_in_6),
            .DOUT0(N__6581),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_4_iopad (
            .OE(N__7716),
            .DIN(N__7715),
            .DOUT(N__7714),
            .PACKAGEPIN(D_LM_AMIGA[4]));
    defparam D_LM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_4_preio (
            .PADOEN(N__7716),
            .PADOUT(N__7715),
            .PADIN(N__7714),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2674),
            .DIN0(D_LM_AMIGA_in_4),
            .DOUT0(N__6095),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_1_iopad (
            .OE(N__7707),
            .DIN(N__7706),
            .DOUT(N__7705),
            .PACKAGEPIN(A_AMIGA[1]));
    defparam A_AMIGA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_1_preio (
            .PADOEN(N__7707),
            .PADOUT(N__7706),
            .PADIN(N__7705),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3205),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_7_iopad (
            .OE(N__7698),
            .DIN(N__7697),
            .DOUT(N__7696),
            .PACKAGEPIN(D_LM_040[7]));
    defparam D_LM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_7_preio (
            .PADOEN(N__7698),
            .PADOUT(N__7697),
            .PADIN(N__7696),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3812),
            .DIN0(D_LM_040_in_7),
            .DOUT0(N__3230),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_4_iopad (
            .OE(N__7689),
            .DIN(N__7688),
            .DOUT(N__7687),
            .PACKAGEPIN(D_UM_040[4]));
    defparam D_UM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_4_preio (
            .PADOEN(N__7689),
            .PADOUT(N__7688),
            .PADIN(N__7687),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3932),
            .DIN0(D_UM_040_in_4),
            .DOUT0(N__4376),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_obuf_iopad (
            .OE(N__7680),
            .DIN(N__7679),
            .DOUT(N__7678),
            .PACKAGEPIN(CLK40B));
    defparam CLK40B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_obuf_preio (
            .PADOEN(N__7680),
            .PADOUT(N__7679),
            .PADIN(N__7678),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5546),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_0_iopad (
            .OE(N__7671),
            .DIN(N__7670),
            .DOUT(N__7669),
            .PACKAGEPIN(D_UU_AMIGA[0]));
    defparam D_UU_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_0_preio (
            .PADOEN(N__7671),
            .PADOUT(N__7670),
            .PADIN(N__7669),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2834),
            .DIN0(D_UU_AMIGA_in_0),
            .DOUT0(N__4292),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_0_iopad (
            .OE(N__7662),
            .DIN(N__7661),
            .DOUT(N__7660),
            .PACKAGEPIN(A_040[0]));
    defparam A_040_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_0_preio (
            .PADOEN(N__7662),
            .PADOUT(N__7661),
            .PADIN(N__7660),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_0_iopad (
            .OE(N__7653),
            .DIN(N__7652),
            .DOUT(N__7651),
            .PACKAGEPIN(D_LM_AMIGA[0]));
    defparam D_LM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_0_preio (
            .PADOEN(N__7653),
            .PADOUT(N__7652),
            .PADIN(N__7651),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2783),
            .DIN0(D_LM_AMIGA_in_0),
            .DOUT0(N__4334),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_1_iopad (
            .OE(N__7644),
            .DIN(N__7643),
            .DOUT(N__7642),
            .PACKAGEPIN(D_UM_040[1]));
    defparam D_UM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_1_preio (
            .PADOEN(N__7644),
            .PADOUT(N__7643),
            .PADIN(N__7642),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3887),
            .DIN0(D_UM_040_in_1),
            .DOUT0(N__4520),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBI_CPUn_obuf_iopad (
            .OE(N__7635),
            .DIN(N__7634),
            .DOUT(N__7633),
            .PACKAGEPIN(TBI_CPUn));
    defparam TBI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TBI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TBI_CPUn_obuf_preio (
            .PADOEN(N__7635),
            .PADOUT(N__7634),
            .PADIN(N__7633),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40A_obuf_iopad (
            .OE(N__7626),
            .DIN(N__7625),
            .DOUT(N__7624),
            .PACKAGEPIN(CLK40A));
    defparam CLK40A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40A_obuf_preio (
            .PADOEN(N__7626),
            .PADOUT(N__7625),
            .PADIN(N__7624),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5545),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_3_iopad (
            .OE(N__7617),
            .DIN(N__7616),
            .DOUT(N__7615),
            .PACKAGEPIN(D_LM_040[3]));
    defparam D_LM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_3_preio (
            .PADOEN(N__7617),
            .PADOUT(N__7616),
            .PADIN(N__7615),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3923),
            .DIN0(D_LM_040_in_3),
            .DOUT0(N__2324),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_4_iopad (
            .OE(N__7608),
            .DIN(N__7607),
            .DOUT(N__7606),
            .PACKAGEPIN(D_LL_040[4]));
    defparam D_LL_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_4_preio (
            .PADOEN(N__7608),
            .PADOUT(N__7607),
            .PADIN(N__7606),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4020),
            .DIN0(D_LL_040_in_4),
            .DOUT0(N__3266),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_7_iopad (
            .OE(N__7599),
            .DIN(N__7598),
            .DOUT(N__7597),
            .PACKAGEPIN(D_LL_AMIGA[7]));
    defparam D_LL_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_7_preio (
            .PADOEN(N__7599),
            .PADOUT(N__7598),
            .PADIN(N__7597),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2782),
            .DIN0(D_LL_AMIGA_in_7),
            .DOUT0(N__3173),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_7_iopad (
            .OE(N__7590),
            .DIN(N__7589),
            .DOUT(N__7588),
            .PACKAGEPIN(D_UU_AMIGA[7]));
    defparam D_UU_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_7_preio (
            .PADOEN(N__7590),
            .PADOUT(N__7589),
            .PADIN(N__7588),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2836),
            .DIN0(D_UU_AMIGA_in_7),
            .DOUT0(N__6734),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFDIR_obuf_iopad (
            .OE(N__7581),
            .DIN(N__7580),
            .DOUT(N__7579),
            .PACKAGEPIN(BUFDIR));
    defparam BUFDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFDIR_obuf_preio (
            .PADOEN(N__7581),
            .PADOUT(N__7580),
            .PADIN(N__7579),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4002),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_5_iopad (
            .OE(N__7572),
            .DIN(N__7571),
            .DOUT(N__7570),
            .PACKAGEPIN(D_LM_AMIGA[5]));
    defparam D_LM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_5_preio (
            .PADOEN(N__7572),
            .PADOUT(N__7571),
            .PADIN(N__7570),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2710),
            .DIN0(D_LM_AMIGA_in_5),
            .DOUT0(N__6878),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_4_iopad (
            .OE(N__7563),
            .DIN(N__7562),
            .DOUT(N__7561),
            .PACKAGEPIN(D_UU_040[4]));
    defparam D_UU_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_4_preio (
            .PADOEN(N__7563),
            .PADOUT(N__7562),
            .PADIN(N__7561),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3970),
            .DIN0(D_UU_040_in_4),
            .DOUT0(N__3374),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SIZ_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__7554),
            .DIN(N__7553),
            .DOUT(N__7552),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__7554),
            .PADOUT(N__7553),
            .PADIN(N__7552),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_6_iopad (
            .OE(N__7545),
            .DIN(N__7544),
            .DOUT(N__7543),
            .PACKAGEPIN(D_LM_040[6]));
    defparam D_LM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_6_preio (
            .PADOEN(N__7545),
            .PADOUT(N__7544),
            .PADIN(N__7543),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3792),
            .DIN0(D_LM_040_in_6),
            .DOUT0(N__2516),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_5_iopad (
            .OE(N__7536),
            .DIN(N__7535),
            .DOUT(N__7534),
            .PACKAGEPIN(D_UM_040[5]));
    defparam D_UM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_5_preio (
            .PADOEN(N__7536),
            .PADOUT(N__7535),
            .PADIN(N__7534),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3933),
            .DIN0(D_UM_040_in_5),
            .DOUT0(N__5591),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TS_CPUn_ibuf_iopad (
            .OE(N__7527),
            .DIN(N__7526),
            .DOUT(N__7525),
            .PACKAGEPIN(TS_CPUn));
    defparam TS_CPUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TS_CPUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TS_CPUn_ibuf_preio (
            .PADOEN(N__7527),
            .PADOUT(N__7526),
            .PADIN(N__7525),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TS_CPUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_1_iopad (
            .OE(N__7518),
            .DIN(N__7517),
            .DOUT(N__7516),
            .PACKAGEPIN(D_LL_040[1]));
    defparam D_LL_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_1_preio (
            .PADOEN(N__7518),
            .PADOUT(N__7517),
            .PADIN(N__7516),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4019),
            .DIN0(D_LL_040_in_1),
            .DOUT0(N__2363),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_3_iopad (
            .OE(N__7509),
            .DIN(N__7508),
            .DOUT(N__7507),
            .PACKAGEPIN(D_LL_AMIGA[3]));
    defparam D_LL_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_3_preio (
            .PADOEN(N__7509),
            .PADOUT(N__7508),
            .PADIN(N__7507),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2838),
            .DIN0(D_LL_AMIGA_in_3),
            .DOUT0(N__6565),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_5_iopad (
            .OE(N__7500),
            .DIN(N__7499),
            .DOUT(N__7498),
            .PACKAGEPIN(D_UM_AMIGA[5]));
    defparam D_UM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_5_preio (
            .PADOEN(N__7500),
            .PADOUT(N__7499),
            .PADIN(N__7498),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2835),
            .DIN0(D_UM_AMIGA_in_5),
            .DOUT0(N__5807),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_1_iopad (
            .OE(N__7491),
            .DIN(N__7490),
            .DOUT(N__7489),
            .PACKAGEPIN(D_UU_040[1]));
    defparam D_UU_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_1_preio (
            .PADOEN(N__7491),
            .PADOUT(N__7490),
            .PADIN(N__7489),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3890),
            .DIN0(D_UU_040_in_1),
            .DOUT0(N__4454),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_3_iopad (
            .OE(N__7482),
            .DIN(N__7481),
            .DOUT(N__7480),
            .PACKAGEPIN(D_UU_AMIGA[3]));
    defparam D_UU_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_3_preio (
            .PADOEN(N__7482),
            .PADOUT(N__7481),
            .PADIN(N__7480),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2820),
            .DIN0(D_UU_AMIGA_in_3),
            .DOUT0(N__2426),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_1_iopad (
            .OE(N__7473),
            .DIN(N__7472),
            .DOUT(N__7471),
            .PACKAGEPIN(D_LM_AMIGA[1]));
    defparam D_LM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_1_preio (
            .PADOEN(N__7473),
            .PADOUT(N__7472),
            .PADIN(N__7471),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2671),
            .DIN0(D_LM_AMIGA_in_1),
            .DOUT0(N__3580),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_2_iopad (
            .OE(N__7464),
            .DIN(N__7463),
            .DOUT(N__7462),
            .PACKAGEPIN(D_LM_040[2]));
    defparam D_LM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_2_preio (
            .PADOEN(N__7464),
            .PADOUT(N__7463),
            .PADIN(N__7462),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3978),
            .DIN0(D_LM_040_in_2),
            .DOUT0(N__2213),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_5_iopad (
            .OE(N__7455),
            .DIN(N__7454),
            .DOUT(N__7453),
            .PACKAGEPIN(D_LL_040[5]));
    defparam D_LL_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_5_preio (
            .PADOEN(N__7455),
            .PADOUT(N__7454),
            .PADIN(N__7453),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4005),
            .DIN0(D_LL_040_in_5),
            .DOUT0(N__4955),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_6_iopad (
            .OE(N__7446),
            .DIN(N__7445),
            .DOUT(N__7444),
            .PACKAGEPIN(D_LL_AMIGA[6]));
    defparam D_LL_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_6_preio (
            .PADOEN(N__7446),
            .PADOUT(N__7445),
            .PADIN(N__7444),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2784),
            .DIN0(D_LL_AMIGA_in_6),
            .DOUT0(N__6647),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_6_iopad (
            .OE(N__7437),
            .DIN(N__7436),
            .DOUT(N__7435),
            .PACKAGEPIN(D_UU_AMIGA[6]));
    defparam D_UU_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_6_preio (
            .PADOEN(N__7437),
            .PADOUT(N__7436),
            .PADIN(N__7435),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2837),
            .DIN0(D_UU_AMIGA_in_6),
            .DOUT0(N__3050),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_1_iopad (
            .OE(N__7428),
            .DIN(N__7427),
            .DOUT(N__7426),
            .PACKAGEPIN(D_UM_AMIGA[1]));
    defparam D_UM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_1_preio (
            .PADOEN(N__7428),
            .PADOUT(N__7427),
            .PADIN(N__7426),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2711),
            .DIN0(D_UM_AMIGA_in_1),
            .DOUT0(N__2858),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_5_iopad (
            .OE(N__7419),
            .DIN(N__7418),
            .DOUT(N__7417),
            .PACKAGEPIN(D_UU_040[5]));
    defparam D_UU_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_5_preio (
            .PADOEN(N__7419),
            .PADOUT(N__7418),
            .PADIN(N__7417),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3934),
            .DIN0(D_UU_040_in_5),
            .DOUT0(N__5729),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMA_obuf_iopad (
            .OE(N__7410),
            .DIN(N__7409),
            .DOUT(N__7408),
            .PACKAGEPIN(CLKRAMA));
    defparam CLKRAMA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMA_obuf_preio (
            .PADOEN(N__7410),
            .PADOUT(N__7409),
            .PADIN(N__7408),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6935),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_2_iopad (
            .OE(N__7401),
            .DIN(N__7400),
            .DOUT(N__7399),
            .PACKAGEPIN(D_UM_040[2]));
    defparam D_UM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_2_preio (
            .PADOEN(N__7401),
            .PADOUT(N__7400),
            .PADIN(N__7399),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3833),
            .DIN0(D_UM_040_in_2),
            .DOUT0(N__4814),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_2_iopad (
            .OE(N__7392),
            .DIN(N__7391),
            .DOUT(N__7390),
            .PACKAGEPIN(D_LL_040[2]));
    defparam D_LL_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_2_preio (
            .PADOEN(N__7392),
            .PADOUT(N__7391),
            .PADIN(N__7390),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4007),
            .DIN0(D_LL_040_in_2),
            .DOUT0(N__2243),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TCI_CPUn_obuf_iopad.PULLUP=1'b1;
    IO_PAD TCI_CPUn_obuf_iopad (
            .OE(N__7383),
            .DIN(N__7382),
            .DOUT(N__7381),
            .PACKAGEPIN(TCI_CPUn));
    defparam TCI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TCI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TCI_CPUn_obuf_preio (
            .PADOEN(N__7383),
            .PADOUT(N__7382),
            .PADIN(N__7381),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7023),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMB_obuf_iopad (
            .OE(N__7374),
            .DIN(N__7373),
            .DOUT(N__7372),
            .PACKAGEPIN(CLKRAMB));
    defparam CLKRAMB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMB_obuf_preio (
            .PADOEN(N__7374),
            .PADOUT(N__7373),
            .PADIN(N__7372),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6928),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_2_iopad (
            .OE(N__7365),
            .DIN(N__7364),
            .DOUT(N__7363),
            .PACKAGEPIN(D_LL_AMIGA[2]));
    defparam D_LL_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_2_preio (
            .PADOEN(N__7365),
            .PADOUT(N__7364),
            .PADIN(N__7363),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2839),
            .DIN0(D_LL_AMIGA_in_2),
            .DOUT0(N__4877),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_4_iopad (
            .OE(N__7356),
            .DIN(N__7355),
            .DOUT(N__7354),
            .PACKAGEPIN(D_UM_AMIGA[4]));
    defparam D_UM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_4_preio (
            .PADOEN(N__7356),
            .PADOUT(N__7355),
            .PADIN(N__7354),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2781),
            .DIN0(D_UM_AMIGA_in_4),
            .DOUT0(N__5963),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_2_iopad (
            .OE(N__7347),
            .DIN(N__7346),
            .DOUT(N__7345),
            .PACKAGEPIN(D_UU_AMIGA[2]));
    defparam D_UU_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_2_preio (
            .PADOEN(N__7347),
            .PADOUT(N__7346),
            .PADIN(N__7345),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2833),
            .DIN0(D_UU_AMIGA_in_2),
            .DOUT0(N__4220),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__7338),
            .DIN(N__7337),
            .DOUT(N__7336),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__7338),
            .PADOUT(N__7337),
            .PADIN(N__7336),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_6_iopad (
            .OE(N__7329),
            .DIN(N__7328),
            .DOUT(N__7327),
            .PACKAGEPIN(D_LM_AMIGA[6]));
    defparam D_LM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_6_preio (
            .PADOEN(N__7329),
            .PADOUT(N__7328),
            .PADIN(N__7327),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2713),
            .DIN0(D_LM_AMIGA_in_6),
            .DOUT0(N__3110),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam RnW_ibuf_iopad.PULLUP=1'b1;
    IO_PAD RnW_ibuf_iopad (
            .OE(N__7320),
            .DIN(N__7319),
            .DOUT(N__7318),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__7320),
            .PADOUT(N__7319),
            .PADIN(N__7318),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_5_iopad (
            .OE(N__7311),
            .DIN(N__7310),
            .DOUT(N__7309),
            .PACKAGEPIN(D_LM_040[5]));
    defparam D_LM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_5_preio (
            .PADOEN(N__7311),
            .PADOUT(N__7310),
            .PADIN(N__7309),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3835),
            .DIN0(D_LM_040_in_5),
            .DOUT0(N__2549),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_6_iopad (
            .OE(N__7302),
            .DIN(N__7301),
            .DOUT(N__7300),
            .PACKAGEPIN(D_UM_040[6]));
    defparam D_UM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_6_preio (
            .PADOEN(N__7302),
            .PADOUT(N__7301),
            .PADIN(N__7300),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3796),
            .DIN0(D_UM_040_in_6),
            .DOUT0(N__5318),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TAn_obuf_iopad.PULLUP=1'b1;
    IO_PAD TAn_obuf_iopad (
            .OE(N__7293),
            .DIN(N__7292),
            .DOUT(N__7291),
            .PACKAGEPIN(TAn));
    defparam TAn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TAn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TAn_obuf_preio (
            .PADOEN(N__7293),
            .PADOUT(N__7292),
            .PADIN(N__7291),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4634),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMAn_obuf_iopad (
            .OE(N__7284),
            .DIN(N__7283),
            .DOUT(N__7282),
            .PACKAGEPIN(DMAn));
    defparam DMAn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMAn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMAn_obuf_preio (
            .PADOEN(N__7284),
            .PADOUT(N__7283),
            .PADIN(N__7282),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7031),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_6_iopad (
            .OE(N__7275),
            .DIN(N__7274),
            .DOUT(N__7273),
            .PACKAGEPIN(D_LL_040[6]));
    defparam D_LL_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_6_preio (
            .PADOEN(N__7275),
            .PADOUT(N__7274),
            .PADIN(N__7273),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4006),
            .DIN0(D_LL_040_in_6),
            .DOUT0(N__4109),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_5_iopad (
            .OE(N__7266),
            .DIN(N__7265),
            .DOUT(N__7264),
            .PACKAGEPIN(D_LL_AMIGA[5]));
    defparam D_LL_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_5_preio (
            .PADOEN(N__7266),
            .PADOUT(N__7265),
            .PADIN(N__7264),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2785),
            .DIN0(D_LL_AMIGA_in_5),
            .DOUT0(N__5849),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_0_iopad (
            .OE(N__7257),
            .DIN(N__7256),
            .DOUT(N__7255),
            .PACKAGEPIN(D_UM_AMIGA[0]));
    defparam D_UM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_0_preio (
            .PADOEN(N__7257),
            .PADOUT(N__7256),
            .PADIN(N__7255),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2673),
            .DIN0(D_UM_AMIGA_in_0),
            .DOUT0(N__6662),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_2_iopad (
            .OE(N__7248),
            .DIN(N__7247),
            .DOUT(N__7246),
            .PACKAGEPIN(D_UU_040[2]));
    defparam D_UU_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_2_preio (
            .PADOEN(N__7248),
            .PADOUT(N__7247),
            .PADIN(N__7246),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3969),
            .DIN0(D_UU_040_in_2),
            .DOUT0(N__5657),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_2_iopad (
            .OE(N__7239),
            .DIN(N__7238),
            .DOUT(N__7237),
            .PACKAGEPIN(D_LM_AMIGA[2]));
    defparam D_LM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_2_preio (
            .PADOEN(N__7239),
            .PADOUT(N__7238),
            .PADIN(N__7237),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2672),
            .DIN0(D_LM_AMIGA_in_2),
            .DOUT0(N__4256),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK80_CPU_obuf_iopad (
            .OE(N__7230),
            .DIN(N__7229),
            .DOUT(N__7228),
            .PACKAGEPIN(CLK80_CPU));
    defparam CLK80_CPU_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK80_CPU_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK80_CPU_obuf_preio (
            .PADOEN(N__7230),
            .PADOUT(N__7229),
            .PADIN(N__7228),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6927),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_3_iopad (
            .OE(N__7221),
            .DIN(N__7220),
            .DOUT(N__7219),
            .PACKAGEPIN(D_LL_040[3]));
    defparam D_LL_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_3_preio (
            .PADOEN(N__7221),
            .PADOUT(N__7220),
            .PADIN(N__7219),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4027),
            .DIN0(D_LL_040_in_3),
            .DOUT0(N__3017),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_1_iopad (
            .OE(N__7212),
            .DIN(N__7211),
            .DOUT(N__7210),
            .PACKAGEPIN(D_LM_040[1]));
    defparam D_LM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_1_preio (
            .PADOEN(N__7212),
            .PADOUT(N__7211),
            .PADIN(N__7210),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3977),
            .DIN0(D_LM_040_in_1),
            .DOUT0(N__3668),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TSn_obuf_iopad.PULLUP=1'b1;
    IO_PAD TSn_obuf_iopad (
            .OE(N__7203),
            .DIN(N__7202),
            .DOUT(N__7201),
            .PACKAGEPIN(TSn));
    defparam TSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TSn_obuf_preio (
            .PADOEN(N__7203),
            .PADOUT(N__7202),
            .PADIN(N__7201),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4064),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_7_iopad (
            .OE(N__7194),
            .DIN(N__7193),
            .DOUT(N__7192),
            .PACKAGEPIN(D_UM_AMIGA[7]));
    defparam D_UM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_7_preio (
            .PADOEN(N__7194),
            .PADOUT(N__7193),
            .PADIN(N__7192),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2780),
            .DIN0(D_UM_AMIGA_in_7),
            .DOUT0(N__3128),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_7_iopad (
            .OE(N__7185),
            .DIN(N__7184),
            .DOUT(N__7183),
            .PACKAGEPIN(D_LM_AMIGA[7]));
    defparam D_LM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_7_preio (
            .PADOEN(N__7185),
            .PADOUT(N__7184),
            .PADIN(N__7183),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2712),
            .DIN0(D_LM_AMIGA_in_7),
            .DOUT0(N__6794),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PORTSIZE_ibuf_iopad.PULLUP=1'b1;
    IO_PAD PORTSIZE_ibuf_iopad (
            .OE(N__7176),
            .DIN(N__7175),
            .DOUT(N__7174),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PORTSIZE_ibuf_preio (
            .PADOEN(N__7176),
            .PADOUT(N__7175),
            .PADIN(N__7174),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PORTSIZE_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_0_iopad (
            .OE(N__7167),
            .DIN(N__7166),
            .DOUT(N__7165),
            .PACKAGEPIN(A_AMIGA[0]));
    defparam A_AMIGA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_0_preio (
            .PADOEN(N__7167),
            .PADOUT(N__7166),
            .PADIN(N__7165),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2273),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_4_iopad (
            .OE(N__7158),
            .DIN(N__7157),
            .DOUT(N__7156),
            .PACKAGEPIN(D_LM_040[4]));
    defparam D_LM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_4_preio (
            .PADOEN(N__7158),
            .PADOUT(N__7157),
            .PADIN(N__7156),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3880),
            .DIN0(D_LM_040_in_4),
            .DOUT0(N__2588),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_7_iopad (
            .OE(N__7149),
            .DIN(N__7148),
            .DOUT(N__7147),
            .PACKAGEPIN(D_UM_040[7]));
    defparam D_UM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_7_preio (
            .PADOEN(N__7149),
            .PADOUT(N__7148),
            .PADIN(N__7147),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3888),
            .DIN0(D_UM_040_in_7),
            .DOUT0(N__4997),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__7140),
            .DIN(N__7139),
            .DOUT(N__7138),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__7140),
            .PADOUT(N__7139),
            .PADIN(N__7138),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_1_iopad (
            .OE(N__7131),
            .DIN(N__7130),
            .DOUT(N__7129),
            .PACKAGEPIN(D_UU_AMIGA[1]));
    defparam D_UU_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_1_preio (
            .PADOEN(N__7131),
            .PADOUT(N__7130),
            .PADIN(N__7129),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2778),
            .DIN0(D_UU_AMIGA_in_1),
            .DOUT0(N__3509),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__7122),
            .DIN(N__7121),
            .DOUT(N__7120),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__7122),
            .PADOUT(N__7121),
            .PADIN(N__7120),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5544),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_0_iopad (
            .OE(N__7113),
            .DIN(N__7112),
            .DOUT(N__7111),
            .PACKAGEPIN(D_UM_040[0]));
    defparam D_UM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_0_preio (
            .PADOEN(N__7113),
            .PADOUT(N__7112),
            .PADIN(N__7111),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3834),
            .DIN0(D_UM_040_in_0),
            .DOUT0(N__2996),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_0_iopad (
            .OE(N__7104),
            .DIN(N__7103),
            .DOUT(N__7102),
            .PACKAGEPIN(D_LL_AMIGA[0]));
    defparam D_LL_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_0_preio (
            .PADOEN(N__7104),
            .PADOUT(N__7103),
            .PADIN(N__7102),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2840),
            .DIN0(D_LL_AMIGA_in_0),
            .DOUT0(N__6707),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_4_iopad (
            .OE(N__7095),
            .DIN(N__7094),
            .DOUT(N__7093),
            .PACKAGEPIN(D_UU_AMIGA[4]));
    defparam D_UU_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_4_preio (
            .PADOEN(N__7095),
            .PADOUT(N__7094),
            .PADIN(N__7093),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2832),
            .DIN0(D_UU_AMIGA_in_4),
            .DOUT0(N__6056),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_7_iopad (
            .OE(N__7086),
            .DIN(N__7085),
            .DOUT(N__7084),
            .PACKAGEPIN(D_UU_040[7]));
    defparam D_UU_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_7_preio (
            .PADOEN(N__7086),
            .PADOUT(N__7085),
            .PADIN(N__7084),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3935),
            .DIN0(D_UU_040_in_7),
            .DOUT0(N__3305),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SIZ_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__7077),
            .DIN(N__7076),
            .DOUT(N__7075),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__7077),
            .PADOUT(N__7076),
            .PADIN(N__7075),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_0_iopad (
            .OE(N__7068),
            .DIN(N__7067),
            .DOUT(N__7066),
            .PACKAGEPIN(D_LL_040[0]));
    defparam D_LL_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_0_preio (
            .PADOEN(N__7068),
            .PADOUT(N__7067),
            .PADIN(N__7066),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4028),
            .DIN0(D_LL_040_in_0),
            .DOUT0(N__2393),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_2_iopad (
            .OE(N__7059),
            .DIN(N__7058),
            .DOUT(N__7057),
            .PACKAGEPIN(D_UM_AMIGA[2]));
    defparam D_UM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_2_preio (
            .PADOEN(N__7059),
            .PADOUT(N__7058),
            .PADIN(N__7057),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2675),
            .DIN0(D_UM_AMIGA_in_2),
            .DOUT0(N__4835),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_0_iopad (
            .OE(N__7050),
            .DIN(N__7049),
            .DOUT(N__7048),
            .PACKAGEPIN(D_UU_040[0]));
    defparam D_UU_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_0_preio (
            .PADOEN(N__7050),
            .PADOUT(N__7049),
            .PADIN(N__7048),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3871),
            .DIN0(D_UU_040_in_0),
            .DOUT0(N__4148),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__1804 (
            .O(N__7031),
            .I(N__7027));
    IoInMux I__1803 (
            .O(N__7030),
            .I(N__7024));
    LocalMux I__1802 (
            .O(N__7027),
            .I(N__7020));
    LocalMux I__1801 (
            .O(N__7024),
            .I(N__7017));
    IoInMux I__1800 (
            .O(N__7023),
            .I(N__7014));
    Span4Mux_s3_v I__1799 (
            .O(N__7020),
            .I(N__7011));
    IoSpan4Mux I__1798 (
            .O(N__7017),
            .I(N__7008));
    LocalMux I__1797 (
            .O(N__7014),
            .I(N__7005));
    Span4Mux_h I__1796 (
            .O(N__7011),
            .I(N__7002));
    Span4Mux_s1_v I__1795 (
            .O(N__7008),
            .I(N__6999));
    Span4Mux_s2_h I__1794 (
            .O(N__7005),
            .I(N__6996));
    Sp12to4 I__1793 (
            .O(N__7002),
            .I(N__6993));
    Span4Mux_v I__1792 (
            .O(N__6999),
            .I(N__6990));
    Span4Mux_h I__1791 (
            .O(N__6996),
            .I(N__6987));
    Span12Mux_h I__1790 (
            .O(N__6993),
            .I(N__6984));
    Span4Mux_v I__1789 (
            .O(N__6990),
            .I(N__6979));
    Span4Mux_v I__1788 (
            .O(N__6987),
            .I(N__6979));
    Odrv12 I__1787 (
            .O(N__6984),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1786 (
            .O(N__6979),
            .I(CONSTANT_ONE_NET));
    InMux I__1785 (
            .O(N__6974),
            .I(N__6971));
    LocalMux I__1784 (
            .O(N__6971),
            .I(N__6960));
    ClkMux I__1783 (
            .O(N__6970),
            .I(N__6938));
    ClkMux I__1782 (
            .O(N__6969),
            .I(N__6938));
    ClkMux I__1781 (
            .O(N__6968),
            .I(N__6938));
    ClkMux I__1780 (
            .O(N__6967),
            .I(N__6938));
    ClkMux I__1779 (
            .O(N__6966),
            .I(N__6938));
    ClkMux I__1778 (
            .O(N__6965),
            .I(N__6938));
    ClkMux I__1777 (
            .O(N__6964),
            .I(N__6938));
    ClkMux I__1776 (
            .O(N__6963),
            .I(N__6938));
    Glb2LocalMux I__1775 (
            .O(N__6960),
            .I(N__6938));
    ClkMux I__1774 (
            .O(N__6959),
            .I(N__6938));
    GlobalMux I__1773 (
            .O(N__6938),
            .I(CLK80));
    IoInMux I__1772 (
            .O(N__6935),
            .I(N__6932));
    LocalMux I__1771 (
            .O(N__6932),
            .I(N__6929));
    IoSpan4Mux I__1770 (
            .O(N__6929),
            .I(N__6924));
    IoInMux I__1769 (
            .O(N__6928),
            .I(N__6921));
    IoInMux I__1768 (
            .O(N__6927),
            .I(N__6918));
    IoSpan4Mux I__1767 (
            .O(N__6924),
            .I(N__6915));
    LocalMux I__1766 (
            .O(N__6921),
            .I(N__6912));
    LocalMux I__1765 (
            .O(N__6918),
            .I(N__6909));
    Span4Mux_s3_v I__1764 (
            .O(N__6915),
            .I(N__6904));
    Span4Mux_s3_v I__1763 (
            .O(N__6912),
            .I(N__6904));
    IoSpan4Mux I__1762 (
            .O(N__6909),
            .I(N__6901));
    Span4Mux_v I__1761 (
            .O(N__6904),
            .I(N__6898));
    Span4Mux_s3_h I__1760 (
            .O(N__6901),
            .I(N__6895));
    Span4Mux_v I__1759 (
            .O(N__6898),
            .I(N__6892));
    Span4Mux_h I__1758 (
            .O(N__6895),
            .I(N__6889));
    Span4Mux_v I__1757 (
            .O(N__6892),
            .I(N__6886));
    Sp12to4 I__1756 (
            .O(N__6889),
            .I(N__6883));
    Odrv4 I__1755 (
            .O(N__6886),
            .I(GB_BUFFER_CLK80_THRU_CO));
    Odrv12 I__1754 (
            .O(N__6883),
            .I(GB_BUFFER_CLK80_THRU_CO));
    IoInMux I__1753 (
            .O(N__6878),
            .I(N__6875));
    LocalMux I__1752 (
            .O(N__6875),
            .I(N__6872));
    IoSpan4Mux I__1751 (
            .O(N__6872),
            .I(N__6868));
    InMux I__1750 (
            .O(N__6871),
            .I(N__6865));
    Span4Mux_s2_h I__1749 (
            .O(N__6868),
            .I(N__6862));
    LocalMux I__1748 (
            .O(N__6865),
            .I(N__6859));
    Span4Mux_v I__1747 (
            .O(N__6862),
            .I(N__6856));
    Span4Mux_v I__1746 (
            .O(N__6859),
            .I(N__6853));
    Sp12to4 I__1745 (
            .O(N__6856),
            .I(N__6850));
    Sp12to4 I__1744 (
            .O(N__6853),
            .I(N__6847));
    Span12Mux_s9_h I__1743 (
            .O(N__6850),
            .I(N__6844));
    Span12Mux_h I__1742 (
            .O(N__6847),
            .I(N__6841));
    Span12Mux_h I__1741 (
            .O(N__6844),
            .I(N__6838));
    Span12Mux_v I__1740 (
            .O(N__6841),
            .I(N__6835));
    Odrv12 I__1739 (
            .O(N__6838),
            .I(D_LM_040_in_5));
    Odrv12 I__1738 (
            .O(N__6835),
            .I(D_LM_040_in_5));
    InMux I__1737 (
            .O(N__6830),
            .I(N__6827));
    LocalMux I__1736 (
            .O(N__6827),
            .I(N__6824));
    Span4Mux_v I__1735 (
            .O(N__6824),
            .I(N__6821));
    Span4Mux_v I__1734 (
            .O(N__6821),
            .I(N__6818));
    Sp12to4 I__1733 (
            .O(N__6818),
            .I(N__6815));
    Span12Mux_h I__1732 (
            .O(N__6815),
            .I(N__6812));
    Odrv12 I__1731 (
            .O(N__6812),
            .I(D_UU_040_in_5));
    IoInMux I__1730 (
            .O(N__6809),
            .I(N__6806));
    LocalMux I__1729 (
            .O(N__6806),
            .I(N__6803));
    Span12Mux_s3_h I__1728 (
            .O(N__6803),
            .I(N__6800));
    Span12Mux_h I__1727 (
            .O(N__6800),
            .I(N__6797));
    Odrv12 I__1726 (
            .O(N__6797),
            .I(un1_D_UU_040_5));
    IoInMux I__1725 (
            .O(N__6794),
            .I(N__6791));
    LocalMux I__1724 (
            .O(N__6791),
            .I(N__6788));
    Span4Mux_s1_h I__1723 (
            .O(N__6788),
            .I(N__6784));
    InMux I__1722 (
            .O(N__6787),
            .I(N__6781));
    Sp12to4 I__1721 (
            .O(N__6784),
            .I(N__6778));
    LocalMux I__1720 (
            .O(N__6781),
            .I(N__6775));
    Span12Mux_s9_v I__1719 (
            .O(N__6778),
            .I(N__6772));
    Span4Mux_v I__1718 (
            .O(N__6775),
            .I(N__6769));
    Span12Mux_h I__1717 (
            .O(N__6772),
            .I(N__6766));
    Span4Mux_h I__1716 (
            .O(N__6769),
            .I(N__6763));
    Span12Mux_h I__1715 (
            .O(N__6766),
            .I(N__6760));
    Sp12to4 I__1714 (
            .O(N__6763),
            .I(N__6757));
    Odrv12 I__1713 (
            .O(N__6760),
            .I(D_LM_040_in_7));
    Odrv12 I__1712 (
            .O(N__6757),
            .I(D_LM_040_in_7));
    InMux I__1711 (
            .O(N__6752),
            .I(N__6749));
    LocalMux I__1710 (
            .O(N__6749),
            .I(N__6746));
    Span4Mux_v I__1709 (
            .O(N__6746),
            .I(N__6743));
    Sp12to4 I__1708 (
            .O(N__6743),
            .I(N__6740));
    Span12Mux_h I__1707 (
            .O(N__6740),
            .I(N__6737));
    Odrv12 I__1706 (
            .O(N__6737),
            .I(D_UU_040_in_7));
    IoInMux I__1705 (
            .O(N__6734),
            .I(N__6731));
    LocalMux I__1704 (
            .O(N__6731),
            .I(N__6728));
    Span12Mux_s11_v I__1703 (
            .O(N__6728),
            .I(N__6725));
    Span12Mux_h I__1702 (
            .O(N__6725),
            .I(N__6722));
    Odrv12 I__1701 (
            .O(N__6722),
            .I(un1_D_UU_040_7));
    InMux I__1700 (
            .O(N__6719),
            .I(N__6716));
    LocalMux I__1699 (
            .O(N__6716),
            .I(N__6713));
    Span12Mux_h I__1698 (
            .O(N__6713),
            .I(N__6710));
    Odrv12 I__1697 (
            .O(N__6710),
            .I(D_UM_040_in_0));
    IoInMux I__1696 (
            .O(N__6707),
            .I(N__6704));
    LocalMux I__1695 (
            .O(N__6704),
            .I(N__6700));
    InMux I__1694 (
            .O(N__6703),
            .I(N__6697));
    IoSpan4Mux I__1693 (
            .O(N__6700),
            .I(N__6694));
    LocalMux I__1692 (
            .O(N__6697),
            .I(N__6691));
    Span4Mux_s2_h I__1691 (
            .O(N__6694),
            .I(N__6688));
    Span4Mux_v I__1690 (
            .O(N__6691),
            .I(N__6685));
    Sp12to4 I__1689 (
            .O(N__6688),
            .I(N__6682));
    Sp12to4 I__1688 (
            .O(N__6685),
            .I(N__6679));
    Span12Mux_h I__1687 (
            .O(N__6682),
            .I(N__6676));
    Span12Mux_v I__1686 (
            .O(N__6679),
            .I(N__6673));
    Span12Mux_h I__1685 (
            .O(N__6676),
            .I(N__6670));
    Span12Mux_h I__1684 (
            .O(N__6673),
            .I(N__6667));
    Odrv12 I__1683 (
            .O(N__6670),
            .I(D_LL_040_in_0));
    Odrv12 I__1682 (
            .O(N__6667),
            .I(D_LL_040_in_0));
    IoInMux I__1681 (
            .O(N__6662),
            .I(N__6659));
    LocalMux I__1680 (
            .O(N__6659),
            .I(N__6656));
    Span12Mux_s4_h I__1679 (
            .O(N__6656),
            .I(N__6653));
    Span12Mux_h I__1678 (
            .O(N__6653),
            .I(N__6650));
    Odrv12 I__1677 (
            .O(N__6650),
            .I(un1_D_UM_040_0));
    IoInMux I__1676 (
            .O(N__6647),
            .I(N__6644));
    LocalMux I__1675 (
            .O(N__6644),
            .I(N__6641));
    IoSpan4Mux I__1674 (
            .O(N__6641),
            .I(N__6637));
    InMux I__1673 (
            .O(N__6640),
            .I(N__6634));
    IoSpan4Mux I__1672 (
            .O(N__6637),
            .I(N__6631));
    LocalMux I__1671 (
            .O(N__6634),
            .I(N__6628));
    Span4Mux_s2_h I__1670 (
            .O(N__6631),
            .I(N__6625));
    Span4Mux_v I__1669 (
            .O(N__6628),
            .I(N__6622));
    Sp12to4 I__1668 (
            .O(N__6625),
            .I(N__6619));
    Sp12to4 I__1667 (
            .O(N__6622),
            .I(N__6616));
    Span12Mux_h I__1666 (
            .O(N__6619),
            .I(N__6613));
    Span12Mux_v I__1665 (
            .O(N__6616),
            .I(N__6610));
    Span12Mux_h I__1664 (
            .O(N__6613),
            .I(N__6607));
    Span12Mux_h I__1663 (
            .O(N__6610),
            .I(N__6604));
    Odrv12 I__1662 (
            .O(N__6607),
            .I(D_LL_040_in_6));
    Odrv12 I__1661 (
            .O(N__6604),
            .I(D_LL_040_in_6));
    InMux I__1660 (
            .O(N__6599),
            .I(N__6596));
    LocalMux I__1659 (
            .O(N__6596),
            .I(N__6593));
    Span4Mux_v I__1658 (
            .O(N__6593),
            .I(N__6590));
    Sp12to4 I__1657 (
            .O(N__6590),
            .I(N__6587));
    Span12Mux_h I__1656 (
            .O(N__6587),
            .I(N__6584));
    Odrv12 I__1655 (
            .O(N__6584),
            .I(D_UM_040_in_6));
    IoInMux I__1654 (
            .O(N__6581),
            .I(N__6578));
    LocalMux I__1653 (
            .O(N__6578),
            .I(N__6575));
    Span12Mux_s6_h I__1652 (
            .O(N__6575),
            .I(N__6572));
    Span12Mux_v I__1651 (
            .O(N__6572),
            .I(N__6569));
    Odrv12 I__1650 (
            .O(N__6569),
            .I(un1_D_UM_040_6));
    InMux I__1649 (
            .O(N__6566),
            .I(N__6562));
    IoInMux I__1648 (
            .O(N__6565),
            .I(N__6559));
    LocalMux I__1647 (
            .O(N__6562),
            .I(N__6556));
    LocalMux I__1646 (
            .O(N__6559),
            .I(N__6553));
    Span4Mux_v I__1645 (
            .O(N__6556),
            .I(N__6550));
    Span4Mux_s3_h I__1644 (
            .O(N__6553),
            .I(N__6547));
    Sp12to4 I__1643 (
            .O(N__6550),
            .I(N__6544));
    Sp12to4 I__1642 (
            .O(N__6547),
            .I(N__6541));
    Span12Mux_h I__1641 (
            .O(N__6544),
            .I(N__6538));
    Span12Mux_v I__1640 (
            .O(N__6541),
            .I(N__6535));
    Span12Mux_v I__1639 (
            .O(N__6538),
            .I(N__6532));
    Span12Mux_h I__1638 (
            .O(N__6535),
            .I(N__6529));
    Span12Mux_v I__1637 (
            .O(N__6532),
            .I(N__6524));
    Span12Mux_h I__1636 (
            .O(N__6529),
            .I(N__6524));
    Odrv12 I__1635 (
            .O(N__6524),
            .I(D_LL_040_in_3));
    InMux I__1634 (
            .O(N__6521),
            .I(N__6518));
    LocalMux I__1633 (
            .O(N__6518),
            .I(N__6515));
    Sp12to4 I__1632 (
            .O(N__6515),
            .I(N__6512));
    Span12Mux_v I__1631 (
            .O(N__6512),
            .I(N__6509));
    Span12Mux_h I__1630 (
            .O(N__6509),
            .I(N__6506));
    Odrv12 I__1629 (
            .O(N__6506),
            .I(D_UM_040_in_3));
    IoInMux I__1628 (
            .O(N__6503),
            .I(N__6500));
    LocalMux I__1627 (
            .O(N__6500),
            .I(N__6497));
    IoSpan4Mux I__1626 (
            .O(N__6497),
            .I(N__6494));
    Span4Mux_s3_h I__1625 (
            .O(N__6494),
            .I(N__6491));
    Sp12to4 I__1624 (
            .O(N__6491),
            .I(N__6488));
    Span12Mux_h I__1623 (
            .O(N__6488),
            .I(N__6485));
    Odrv12 I__1622 (
            .O(N__6485),
            .I(un1_D_UM_040_3));
    InMux I__1621 (
            .O(N__6482),
            .I(N__6479));
    LocalMux I__1620 (
            .O(N__6479),
            .I(N__6476));
    Span4Mux_v I__1619 (
            .O(N__6476),
            .I(N__6473));
    Sp12to4 I__1618 (
            .O(N__6473),
            .I(N__6470));
    Span12Mux_h I__1617 (
            .O(N__6470),
            .I(N__6467));
    Odrv12 I__1616 (
            .O(N__6467),
            .I(SIZ_c_0));
    InMux I__1615 (
            .O(N__6464),
            .I(N__6461));
    LocalMux I__1614 (
            .O(N__6461),
            .I(N__6458));
    Span4Mux_v I__1613 (
            .O(N__6458),
            .I(N__6455));
    Sp12to4 I__1612 (
            .O(N__6455),
            .I(N__6452));
    Span12Mux_h I__1611 (
            .O(N__6452),
            .I(N__6449));
    Odrv12 I__1610 (
            .O(N__6449),
            .I(SIZ_c_1));
    InMux I__1609 (
            .O(N__6446),
            .I(N__6443));
    LocalMux I__1608 (
            .O(N__6443),
            .I(N__6439));
    InMux I__1607 (
            .O(N__6442),
            .I(N__6436));
    Span4Mux_v I__1606 (
            .O(N__6439),
            .I(N__6433));
    LocalMux I__1605 (
            .O(N__6436),
            .I(N__6430));
    Span4Mux_v I__1604 (
            .O(N__6433),
            .I(N__6427));
    Span4Mux_v I__1603 (
            .O(N__6430),
            .I(N__6424));
    Sp12to4 I__1602 (
            .O(N__6427),
            .I(N__6419));
    Sp12to4 I__1601 (
            .O(N__6424),
            .I(N__6419));
    Span12Mux_h I__1600 (
            .O(N__6419),
            .I(N__6416));
    Span12Mux_v I__1599 (
            .O(N__6416),
            .I(N__6413));
    Odrv12 I__1598 (
            .O(N__6413),
            .I(PORTSIZE_c));
    InMux I__1597 (
            .O(N__6410),
            .I(N__6407));
    LocalMux I__1596 (
            .O(N__6407),
            .I(N__6404));
    Span4Mux_h I__1595 (
            .O(N__6404),
            .I(N__6400));
    InMux I__1594 (
            .O(N__6403),
            .I(N__6397));
    Sp12to4 I__1593 (
            .O(N__6400),
            .I(N__6392));
    LocalMux I__1592 (
            .O(N__6397),
            .I(N__6392));
    Span12Mux_v I__1591 (
            .O(N__6392),
            .I(N__6389));
    Odrv12 I__1590 (
            .O(N__6389),
            .I(\U111_CYCLE_SM.LW_TRANS_0 ));
    InMux I__1589 (
            .O(N__6386),
            .I(N__6383));
    LocalMux I__1588 (
            .O(N__6383),
            .I(N__6380));
    Span4Mux_v I__1587 (
            .O(N__6380),
            .I(N__6377));
    Span4Mux_h I__1586 (
            .O(N__6377),
            .I(N__6374));
    Span4Mux_h I__1585 (
            .O(N__6374),
            .I(N__6371));
    Odrv4 I__1584 (
            .O(N__6371),
            .I(D_UU_040_in_4));
    InMux I__1583 (
            .O(N__6368),
            .I(N__6358));
    InMux I__1582 (
            .O(N__6367),
            .I(N__6355));
    InMux I__1581 (
            .O(N__6366),
            .I(N__6350));
    InMux I__1580 (
            .O(N__6365),
            .I(N__6350));
    InMux I__1579 (
            .O(N__6364),
            .I(N__6347));
    InMux I__1578 (
            .O(N__6363),
            .I(N__6342));
    InMux I__1577 (
            .O(N__6362),
            .I(N__6342));
    InMux I__1576 (
            .O(N__6361),
            .I(N__6338));
    LocalMux I__1575 (
            .O(N__6358),
            .I(N__6335));
    LocalMux I__1574 (
            .O(N__6355),
            .I(N__6330));
    LocalMux I__1573 (
            .O(N__6350),
            .I(N__6330));
    LocalMux I__1572 (
            .O(N__6347),
            .I(N__6321));
    LocalMux I__1571 (
            .O(N__6342),
            .I(N__6321));
    InMux I__1570 (
            .O(N__6341),
            .I(N__6318));
    LocalMux I__1569 (
            .O(N__6338),
            .I(N__6311));
    Span4Mux_v I__1568 (
            .O(N__6335),
            .I(N__6306));
    Span4Mux_v I__1567 (
            .O(N__6330),
            .I(N__6306));
    InMux I__1566 (
            .O(N__6329),
            .I(N__6303));
    InMux I__1565 (
            .O(N__6328),
            .I(N__6300));
    InMux I__1564 (
            .O(N__6327),
            .I(N__6294));
    InMux I__1563 (
            .O(N__6326),
            .I(N__6291));
    Span4Mux_v I__1562 (
            .O(N__6321),
            .I(N__6284));
    LocalMux I__1561 (
            .O(N__6318),
            .I(N__6284));
    InMux I__1560 (
            .O(N__6317),
            .I(N__6281));
    InMux I__1559 (
            .O(N__6316),
            .I(N__6276));
    InMux I__1558 (
            .O(N__6315),
            .I(N__6273));
    InMux I__1557 (
            .O(N__6314),
            .I(N__6270));
    Span4Mux_v I__1556 (
            .O(N__6311),
            .I(N__6262));
    Span4Mux_h I__1555 (
            .O(N__6306),
            .I(N__6262));
    LocalMux I__1554 (
            .O(N__6303),
            .I(N__6262));
    LocalMux I__1553 (
            .O(N__6300),
            .I(N__6259));
    InMux I__1552 (
            .O(N__6299),
            .I(N__6256));
    InMux I__1551 (
            .O(N__6298),
            .I(N__6253));
    InMux I__1550 (
            .O(N__6297),
            .I(N__6250));
    LocalMux I__1549 (
            .O(N__6294),
            .I(N__6244));
    LocalMux I__1548 (
            .O(N__6291),
            .I(N__6241));
    InMux I__1547 (
            .O(N__6290),
            .I(N__6238));
    InMux I__1546 (
            .O(N__6289),
            .I(N__6235));
    Span4Mux_v I__1545 (
            .O(N__6284),
            .I(N__6229));
    LocalMux I__1544 (
            .O(N__6281),
            .I(N__6226));
    InMux I__1543 (
            .O(N__6280),
            .I(N__6223));
    InMux I__1542 (
            .O(N__6279),
            .I(N__6220));
    LocalMux I__1541 (
            .O(N__6276),
            .I(N__6217));
    LocalMux I__1540 (
            .O(N__6273),
            .I(N__6214));
    LocalMux I__1539 (
            .O(N__6270),
            .I(N__6211));
    InMux I__1538 (
            .O(N__6269),
            .I(N__6208));
    Span4Mux_v I__1537 (
            .O(N__6262),
            .I(N__6197));
    Span4Mux_h I__1536 (
            .O(N__6259),
            .I(N__6197));
    LocalMux I__1535 (
            .O(N__6256),
            .I(N__6197));
    LocalMux I__1534 (
            .O(N__6253),
            .I(N__6197));
    LocalMux I__1533 (
            .O(N__6250),
            .I(N__6197));
    InMux I__1532 (
            .O(N__6249),
            .I(N__6194));
    InMux I__1531 (
            .O(N__6248),
            .I(N__6191));
    InMux I__1530 (
            .O(N__6247),
            .I(N__6188));
    Span4Mux_h I__1529 (
            .O(N__6244),
            .I(N__6179));
    Span4Mux_v I__1528 (
            .O(N__6241),
            .I(N__6179));
    LocalMux I__1527 (
            .O(N__6238),
            .I(N__6179));
    LocalMux I__1526 (
            .O(N__6235),
            .I(N__6179));
    InMux I__1525 (
            .O(N__6234),
            .I(N__6174));
    InMux I__1524 (
            .O(N__6233),
            .I(N__6174));
    InMux I__1523 (
            .O(N__6232),
            .I(N__6171));
    Span4Mux_h I__1522 (
            .O(N__6229),
            .I(N__6165));
    Span4Mux_v I__1521 (
            .O(N__6226),
            .I(N__6165));
    LocalMux I__1520 (
            .O(N__6223),
            .I(N__6160));
    LocalMux I__1519 (
            .O(N__6220),
            .I(N__6160));
    Span4Mux_v I__1518 (
            .O(N__6217),
            .I(N__6157));
    Span4Mux_v I__1517 (
            .O(N__6214),
            .I(N__6152));
    Span4Mux_v I__1516 (
            .O(N__6211),
            .I(N__6152));
    LocalMux I__1515 (
            .O(N__6208),
            .I(N__6149));
    Span4Mux_v I__1514 (
            .O(N__6197),
            .I(N__6144));
    LocalMux I__1513 (
            .O(N__6194),
            .I(N__6144));
    LocalMux I__1512 (
            .O(N__6191),
            .I(N__6139));
    LocalMux I__1511 (
            .O(N__6188),
            .I(N__6139));
    Span4Mux_h I__1510 (
            .O(N__6179),
            .I(N__6134));
    LocalMux I__1509 (
            .O(N__6174),
            .I(N__6134));
    LocalMux I__1508 (
            .O(N__6171),
            .I(N__6131));
    InMux I__1507 (
            .O(N__6170),
            .I(N__6128));
    Span4Mux_v I__1506 (
            .O(N__6165),
            .I(N__6125));
    Span12Mux_v I__1505 (
            .O(N__6160),
            .I(N__6122));
    Span4Mux_h I__1504 (
            .O(N__6157),
            .I(N__6115));
    Span4Mux_h I__1503 (
            .O(N__6152),
            .I(N__6115));
    Span4Mux_v I__1502 (
            .O(N__6149),
            .I(N__6115));
    Span4Mux_v I__1501 (
            .O(N__6144),
            .I(N__6104));
    Span4Mux_v I__1500 (
            .O(N__6139),
            .I(N__6104));
    Span4Mux_v I__1499 (
            .O(N__6134),
            .I(N__6104));
    Span4Mux_h I__1498 (
            .O(N__6131),
            .I(N__6104));
    LocalMux I__1497 (
            .O(N__6128),
            .I(N__6104));
    Odrv4 I__1496 (
            .O(N__6125),
            .I(\U111_CYCLE_SM.FLIP ));
    Odrv12 I__1495 (
            .O(N__6122),
            .I(\U111_CYCLE_SM.FLIP ));
    Odrv4 I__1494 (
            .O(N__6115),
            .I(\U111_CYCLE_SM.FLIP ));
    Odrv4 I__1493 (
            .O(N__6104),
            .I(\U111_CYCLE_SM.FLIP ));
    IoInMux I__1492 (
            .O(N__6095),
            .I(N__6092));
    LocalMux I__1491 (
            .O(N__6092),
            .I(N__6089));
    Span4Mux_s1_h I__1490 (
            .O(N__6089),
            .I(N__6086));
    Sp12to4 I__1489 (
            .O(N__6086),
            .I(N__6082));
    InMux I__1488 (
            .O(N__6085),
            .I(N__6079));
    Span12Mux_v I__1487 (
            .O(N__6082),
            .I(N__6076));
    LocalMux I__1486 (
            .O(N__6079),
            .I(N__6073));
    Span12Mux_h I__1485 (
            .O(N__6076),
            .I(N__6070));
    Span12Mux_h I__1484 (
            .O(N__6073),
            .I(N__6067));
    Span12Mux_h I__1483 (
            .O(N__6070),
            .I(N__6064));
    Span12Mux_v I__1482 (
            .O(N__6067),
            .I(N__6061));
    Odrv12 I__1481 (
            .O(N__6064),
            .I(D_LM_040_in_4));
    Odrv12 I__1480 (
            .O(N__6061),
            .I(D_LM_040_in_4));
    IoInMux I__1479 (
            .O(N__6056),
            .I(N__6053));
    LocalMux I__1478 (
            .O(N__6053),
            .I(N__6050));
    IoSpan4Mux I__1477 (
            .O(N__6050),
            .I(N__6047));
    IoSpan4Mux I__1476 (
            .O(N__6047),
            .I(N__6044));
    Span4Mux_s2_v I__1475 (
            .O(N__6044),
            .I(N__6041));
    Span4Mux_v I__1474 (
            .O(N__6041),
            .I(N__6038));
    Odrv4 I__1473 (
            .O(N__6038),
            .I(un1_D_UU_040_4));
    InMux I__1472 (
            .O(N__6035),
            .I(N__6032));
    LocalMux I__1471 (
            .O(N__6032),
            .I(N__6028));
    IoInMux I__1470 (
            .O(N__6031),
            .I(N__6025));
    Span4Mux_v I__1469 (
            .O(N__6028),
            .I(N__6022));
    LocalMux I__1468 (
            .O(N__6025),
            .I(N__6019));
    Span4Mux_h I__1467 (
            .O(N__6022),
            .I(N__6016));
    Span4Mux_s2_h I__1466 (
            .O(N__6019),
            .I(N__6013));
    Sp12to4 I__1465 (
            .O(N__6016),
            .I(N__6010));
    Span4Mux_v I__1464 (
            .O(N__6013),
            .I(N__6007));
    Span12Mux_h I__1463 (
            .O(N__6010),
            .I(N__6004));
    Sp12to4 I__1462 (
            .O(N__6007),
            .I(N__6001));
    Span12Mux_v I__1461 (
            .O(N__6004),
            .I(N__5998));
    Span12Mux_h I__1460 (
            .O(N__6001),
            .I(N__5995));
    Span12Mux_v I__1459 (
            .O(N__5998),
            .I(N__5992));
    Span12Mux_h I__1458 (
            .O(N__5995),
            .I(N__5989));
    Odrv12 I__1457 (
            .O(N__5992),
            .I(D_LL_040_in_4));
    Odrv12 I__1456 (
            .O(N__5989),
            .I(D_LL_040_in_4));
    InMux I__1455 (
            .O(N__5984),
            .I(N__5981));
    LocalMux I__1454 (
            .O(N__5981),
            .I(N__5978));
    Span4Mux_v I__1453 (
            .O(N__5978),
            .I(N__5975));
    Span4Mux_h I__1452 (
            .O(N__5975),
            .I(N__5972));
    Sp12to4 I__1451 (
            .O(N__5972),
            .I(N__5969));
    Span12Mux_h I__1450 (
            .O(N__5969),
            .I(N__5966));
    Odrv12 I__1449 (
            .O(N__5966),
            .I(D_UM_040_in_4));
    IoInMux I__1448 (
            .O(N__5963),
            .I(N__5960));
    LocalMux I__1447 (
            .O(N__5960),
            .I(N__5957));
    Span4Mux_s2_h I__1446 (
            .O(N__5957),
            .I(N__5954));
    Span4Mux_h I__1445 (
            .O(N__5954),
            .I(N__5951));
    Span4Mux_h I__1444 (
            .O(N__5951),
            .I(N__5948));
    Span4Mux_h I__1443 (
            .O(N__5948),
            .I(N__5945));
    Odrv4 I__1442 (
            .O(N__5945),
            .I(un1_D_UM_040_4));
    InMux I__1441 (
            .O(N__5942),
            .I(N__5939));
    LocalMux I__1440 (
            .O(N__5939),
            .I(N__5936));
    Odrv12 I__1439 (
            .O(N__5936),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ));
    InMux I__1438 (
            .O(N__5933),
            .I(N__5930));
    LocalMux I__1437 (
            .O(N__5930),
            .I(N__5927));
    Span4Mux_v I__1436 (
            .O(N__5927),
            .I(N__5922));
    InMux I__1435 (
            .O(N__5926),
            .I(N__5919));
    InMux I__1434 (
            .O(N__5925),
            .I(N__5916));
    Sp12to4 I__1433 (
            .O(N__5922),
            .I(N__5913));
    LocalMux I__1432 (
            .O(N__5919),
            .I(N__5908));
    LocalMux I__1431 (
            .O(N__5916),
            .I(N__5908));
    Span12Mux_h I__1430 (
            .O(N__5913),
            .I(N__5905));
    Span12Mux_v I__1429 (
            .O(N__5908),
            .I(N__5902));
    Span12Mux_v I__1428 (
            .O(N__5905),
            .I(N__5897));
    Span12Mux_h I__1427 (
            .O(N__5902),
            .I(N__5897));
    Odrv12 I__1426 (
            .O(N__5897),
            .I(D_UU_AMIGA_in_3));
    IoInMux I__1425 (
            .O(N__5894),
            .I(N__5891));
    LocalMux I__1424 (
            .O(N__5891),
            .I(N__5888));
    Span4Mux_s3_v I__1423 (
            .O(N__5888),
            .I(N__5885));
    Span4Mux_h I__1422 (
            .O(N__5885),
            .I(N__5882));
    Span4Mux_h I__1421 (
            .O(N__5882),
            .I(N__5879));
    Span4Mux_h I__1420 (
            .O(N__5879),
            .I(N__5876));
    Span4Mux_h I__1419 (
            .O(N__5876),
            .I(N__5873));
    Odrv4 I__1418 (
            .O(N__5873),
            .I(un1_D_UU_AMIGA_3));
    InMux I__1417 (
            .O(N__5870),
            .I(N__5867));
    LocalMux I__1416 (
            .O(N__5867),
            .I(N__5864));
    Span4Mux_v I__1415 (
            .O(N__5864),
            .I(N__5861));
    Span4Mux_h I__1414 (
            .O(N__5861),
            .I(N__5858));
    Sp12to4 I__1413 (
            .O(N__5858),
            .I(N__5855));
    Span12Mux_h I__1412 (
            .O(N__5855),
            .I(N__5852));
    Odrv12 I__1411 (
            .O(N__5852),
            .I(D_UM_040_in_5));
    IoInMux I__1410 (
            .O(N__5849),
            .I(N__5846));
    LocalMux I__1409 (
            .O(N__5846),
            .I(N__5842));
    InMux I__1408 (
            .O(N__5845),
            .I(N__5839));
    IoSpan4Mux I__1407 (
            .O(N__5842),
            .I(N__5836));
    LocalMux I__1406 (
            .O(N__5839),
            .I(N__5833));
    Span4Mux_s3_h I__1405 (
            .O(N__5836),
            .I(N__5830));
    Sp12to4 I__1404 (
            .O(N__5833),
            .I(N__5827));
    Sp12to4 I__1403 (
            .O(N__5830),
            .I(N__5824));
    Span12Mux_v I__1402 (
            .O(N__5827),
            .I(N__5821));
    Span12Mux_v I__1401 (
            .O(N__5824),
            .I(N__5818));
    Span12Mux_v I__1400 (
            .O(N__5821),
            .I(N__5813));
    Span12Mux_h I__1399 (
            .O(N__5818),
            .I(N__5813));
    Span12Mux_h I__1398 (
            .O(N__5813),
            .I(N__5810));
    Odrv12 I__1397 (
            .O(N__5810),
            .I(D_LL_040_in_5));
    IoInMux I__1396 (
            .O(N__5807),
            .I(N__5804));
    LocalMux I__1395 (
            .O(N__5804),
            .I(N__5801));
    IoSpan4Mux I__1394 (
            .O(N__5801),
            .I(N__5798));
    IoSpan4Mux I__1393 (
            .O(N__5798),
            .I(N__5795));
    Span4Mux_s2_v I__1392 (
            .O(N__5795),
            .I(N__5792));
    Span4Mux_v I__1391 (
            .O(N__5792),
            .I(N__5789));
    Odrv4 I__1390 (
            .O(N__5789),
            .I(un1_D_UM_040_5));
    InMux I__1389 (
            .O(N__5786),
            .I(N__5783));
    LocalMux I__1388 (
            .O(N__5783),
            .I(N__5780));
    Span4Mux_v I__1387 (
            .O(N__5780),
            .I(N__5777));
    Odrv4 I__1386 (
            .O(N__5777),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ));
    InMux I__1385 (
            .O(N__5774),
            .I(N__5771));
    LocalMux I__1384 (
            .O(N__5771),
            .I(N__5768));
    Span4Mux_v I__1383 (
            .O(N__5768),
            .I(N__5764));
    InMux I__1382 (
            .O(N__5767),
            .I(N__5761));
    Span4Mux_v I__1381 (
            .O(N__5764),
            .I(N__5756));
    LocalMux I__1380 (
            .O(N__5761),
            .I(N__5756));
    Span4Mux_h I__1379 (
            .O(N__5756),
            .I(N__5752));
    InMux I__1378 (
            .O(N__5755),
            .I(N__5749));
    Span4Mux_v I__1377 (
            .O(N__5752),
            .I(N__5746));
    LocalMux I__1376 (
            .O(N__5749),
            .I(N__5743));
    Span4Mux_h I__1375 (
            .O(N__5746),
            .I(N__5740));
    Span12Mux_v I__1374 (
            .O(N__5743),
            .I(N__5737));
    Span4Mux_h I__1373 (
            .O(N__5740),
            .I(N__5734));
    Odrv12 I__1372 (
            .O(N__5737),
            .I(D_UU_AMIGA_in_5));
    Odrv4 I__1371 (
            .O(N__5734),
            .I(D_UU_AMIGA_in_5));
    IoInMux I__1370 (
            .O(N__5729),
            .I(N__5726));
    LocalMux I__1369 (
            .O(N__5726),
            .I(N__5723));
    Span12Mux_s6_v I__1368 (
            .O(N__5723),
            .I(N__5720));
    Span12Mux_h I__1367 (
            .O(N__5720),
            .I(N__5717));
    Odrv12 I__1366 (
            .O(N__5717),
            .I(un1_D_UU_AMIGA_5));
    InMux I__1365 (
            .O(N__5714),
            .I(N__5711));
    LocalMux I__1364 (
            .O(N__5711),
            .I(N__5708));
    Odrv12 I__1363 (
            .O(N__5708),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ));
    InMux I__1362 (
            .O(N__5705),
            .I(N__5702));
    LocalMux I__1361 (
            .O(N__5702),
            .I(N__5698));
    InMux I__1360 (
            .O(N__5701),
            .I(N__5694));
    Span4Mux_v I__1359 (
            .O(N__5698),
            .I(N__5691));
    InMux I__1358 (
            .O(N__5697),
            .I(N__5688));
    LocalMux I__1357 (
            .O(N__5694),
            .I(N__5685));
    Span4Mux_v I__1356 (
            .O(N__5691),
            .I(N__5680));
    LocalMux I__1355 (
            .O(N__5688),
            .I(N__5680));
    Span4Mux_v I__1354 (
            .O(N__5685),
            .I(N__5677));
    Span4Mux_v I__1353 (
            .O(N__5680),
            .I(N__5674));
    Span4Mux_h I__1352 (
            .O(N__5677),
            .I(N__5671));
    Sp12to4 I__1351 (
            .O(N__5674),
            .I(N__5668));
    Sp12to4 I__1350 (
            .O(N__5671),
            .I(N__5665));
    Span12Mux_h I__1349 (
            .O(N__5668),
            .I(N__5662));
    Odrv12 I__1348 (
            .O(N__5665),
            .I(D_UU_AMIGA_in_2));
    Odrv12 I__1347 (
            .O(N__5662),
            .I(D_UU_AMIGA_in_2));
    IoInMux I__1346 (
            .O(N__5657),
            .I(N__5654));
    LocalMux I__1345 (
            .O(N__5654),
            .I(N__5651));
    Span12Mux_s0_v I__1344 (
            .O(N__5651),
            .I(N__5648));
    Span12Mux_h I__1343 (
            .O(N__5648),
            .I(N__5645));
    Odrv12 I__1342 (
            .O(N__5645),
            .I(un1_D_UU_AMIGA_2));
    InMux I__1341 (
            .O(N__5642),
            .I(N__5639));
    LocalMux I__1340 (
            .O(N__5639),
            .I(N__5636));
    Span4Mux_v I__1339 (
            .O(N__5636),
            .I(N__5632));
    InMux I__1338 (
            .O(N__5635),
            .I(N__5629));
    Span4Mux_v I__1337 (
            .O(N__5632),
            .I(N__5624));
    LocalMux I__1336 (
            .O(N__5629),
            .I(N__5624));
    Span4Mux_v I__1335 (
            .O(N__5624),
            .I(N__5620));
    InMux I__1334 (
            .O(N__5623),
            .I(N__5617));
    Span4Mux_v I__1333 (
            .O(N__5620),
            .I(N__5612));
    LocalMux I__1332 (
            .O(N__5617),
            .I(N__5612));
    Span4Mux_v I__1331 (
            .O(N__5612),
            .I(N__5609));
    Sp12to4 I__1330 (
            .O(N__5609),
            .I(N__5606));
    Span12Mux_h I__1329 (
            .O(N__5606),
            .I(N__5603));
    Odrv12 I__1328 (
            .O(N__5603),
            .I(D_UM_AMIGA_in_5));
    InMux I__1327 (
            .O(N__5600),
            .I(N__5597));
    LocalMux I__1326 (
            .O(N__5597),
            .I(N__5594));
    Odrv12 I__1325 (
            .O(N__5594),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ));
    IoInMux I__1324 (
            .O(N__5591),
            .I(N__5588));
    LocalMux I__1323 (
            .O(N__5588),
            .I(N__5585));
    Span4Mux_s2_v I__1322 (
            .O(N__5585),
            .I(N__5582));
    Span4Mux_h I__1321 (
            .O(N__5582),
            .I(N__5579));
    Span4Mux_v I__1320 (
            .O(N__5579),
            .I(N__5576));
    Sp12to4 I__1319 (
            .O(N__5576),
            .I(N__5573));
    Odrv12 I__1318 (
            .O(N__5573),
            .I(un1_D_UM_AMIGA_5));
    InMux I__1317 (
            .O(N__5570),
            .I(N__5566));
    InMux I__1316 (
            .O(N__5569),
            .I(N__5563));
    LocalMux I__1315 (
            .O(N__5566),
            .I(N__5559));
    LocalMux I__1314 (
            .O(N__5563),
            .I(N__5556));
    ClkMux I__1313 (
            .O(N__5562),
            .I(N__5549));
    Glb2LocalMux I__1312 (
            .O(N__5559),
            .I(N__5549));
    Glb2LocalMux I__1311 (
            .O(N__5556),
            .I(N__5549));
    GlobalMux I__1310 (
            .O(N__5549),
            .I(CLK40));
    IoInMux I__1309 (
            .O(N__5546),
            .I(N__5541));
    IoInMux I__1308 (
            .O(N__5545),
            .I(N__5538));
    IoInMux I__1307 (
            .O(N__5544),
            .I(N__5535));
    LocalMux I__1306 (
            .O(N__5541),
            .I(N__5532));
    LocalMux I__1305 (
            .O(N__5538),
            .I(N__5529));
    LocalMux I__1304 (
            .O(N__5535),
            .I(N__5526));
    Span12Mux_s5_v I__1303 (
            .O(N__5532),
            .I(N__5523));
    Span12Mux_s10_h I__1302 (
            .O(N__5529),
            .I(N__5518));
    Span12Mux_s9_h I__1301 (
            .O(N__5526),
            .I(N__5518));
    Odrv12 I__1300 (
            .O(N__5523),
            .I(GB_BUFFER_CLK40_THRU_CO));
    Odrv12 I__1299 (
            .O(N__5518),
            .I(GB_BUFFER_CLK40_THRU_CO));
    InMux I__1298 (
            .O(N__5513),
            .I(N__5507));
    InMux I__1297 (
            .O(N__5512),
            .I(N__5507));
    LocalMux I__1296 (
            .O(N__5507),
            .I(N__5497));
    InMux I__1295 (
            .O(N__5506),
            .I(N__5488));
    InMux I__1294 (
            .O(N__5505),
            .I(N__5488));
    InMux I__1293 (
            .O(N__5504),
            .I(N__5488));
    InMux I__1292 (
            .O(N__5503),
            .I(N__5488));
    InMux I__1291 (
            .O(N__5502),
            .I(N__5481));
    InMux I__1290 (
            .O(N__5501),
            .I(N__5478));
    InMux I__1289 (
            .O(N__5500),
            .I(N__5473));
    Span4Mux_v I__1288 (
            .O(N__5497),
            .I(N__5470));
    LocalMux I__1287 (
            .O(N__5488),
            .I(N__5467));
    InMux I__1286 (
            .O(N__5487),
            .I(N__5464));
    InMux I__1285 (
            .O(N__5486),
            .I(N__5461));
    InMux I__1284 (
            .O(N__5485),
            .I(N__5456));
    InMux I__1283 (
            .O(N__5484),
            .I(N__5456));
    LocalMux I__1282 (
            .O(N__5481),
            .I(N__5451));
    LocalMux I__1281 (
            .O(N__5478),
            .I(N__5451));
    InMux I__1280 (
            .O(N__5477),
            .I(N__5448));
    InMux I__1279 (
            .O(N__5476),
            .I(N__5445));
    LocalMux I__1278 (
            .O(N__5473),
            .I(N__5441));
    Sp12to4 I__1277 (
            .O(N__5470),
            .I(N__5437));
    Span4Mux_v I__1276 (
            .O(N__5467),
            .I(N__5430));
    LocalMux I__1275 (
            .O(N__5464),
            .I(N__5430));
    LocalMux I__1274 (
            .O(N__5461),
            .I(N__5430));
    LocalMux I__1273 (
            .O(N__5456),
            .I(N__5421));
    Span4Mux_v I__1272 (
            .O(N__5451),
            .I(N__5421));
    LocalMux I__1271 (
            .O(N__5448),
            .I(N__5421));
    LocalMux I__1270 (
            .O(N__5445),
            .I(N__5421));
    InMux I__1269 (
            .O(N__5444),
            .I(N__5418));
    Span4Mux_v I__1268 (
            .O(N__5441),
            .I(N__5413));
    InMux I__1267 (
            .O(N__5440),
            .I(N__5410));
    Span12Mux_h I__1266 (
            .O(N__5437),
            .I(N__5405));
    Span4Mux_v I__1265 (
            .O(N__5430),
            .I(N__5402));
    Span4Mux_v I__1264 (
            .O(N__5421),
            .I(N__5397));
    LocalMux I__1263 (
            .O(N__5418),
            .I(N__5397));
    InMux I__1262 (
            .O(N__5417),
            .I(N__5394));
    InMux I__1261 (
            .O(N__5416),
            .I(N__5391));
    Span4Mux_v I__1260 (
            .O(N__5413),
            .I(N__5386));
    LocalMux I__1259 (
            .O(N__5410),
            .I(N__5386));
    InMux I__1258 (
            .O(N__5409),
            .I(N__5381));
    InMux I__1257 (
            .O(N__5408),
            .I(N__5381));
    Odrv12 I__1256 (
            .O(N__5405),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    Odrv4 I__1255 (
            .O(N__5402),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    Odrv4 I__1254 (
            .O(N__5397),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    LocalMux I__1253 (
            .O(N__5394),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    LocalMux I__1252 (
            .O(N__5391),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    Odrv4 I__1251 (
            .O(N__5386),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    LocalMux I__1250 (
            .O(N__5381),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    InMux I__1249 (
            .O(N__5366),
            .I(N__5363));
    LocalMux I__1248 (
            .O(N__5363),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ));
    InMux I__1247 (
            .O(N__5360),
            .I(N__5357));
    LocalMux I__1246 (
            .O(N__5357),
            .I(N__5354));
    Span4Mux_h I__1245 (
            .O(N__5354),
            .I(N__5350));
    InMux I__1244 (
            .O(N__5353),
            .I(N__5347));
    Span4Mux_v I__1243 (
            .O(N__5350),
            .I(N__5343));
    LocalMux I__1242 (
            .O(N__5347),
            .I(N__5340));
    InMux I__1241 (
            .O(N__5346),
            .I(N__5337));
    Span4Mux_h I__1240 (
            .O(N__5343),
            .I(N__5334));
    Sp12to4 I__1239 (
            .O(N__5340),
            .I(N__5329));
    LocalMux I__1238 (
            .O(N__5337),
            .I(N__5329));
    Sp12to4 I__1237 (
            .O(N__5334),
            .I(N__5324));
    Span12Mux_h I__1236 (
            .O(N__5329),
            .I(N__5324));
    Span12Mux_v I__1235 (
            .O(N__5324),
            .I(N__5321));
    Odrv12 I__1234 (
            .O(N__5321),
            .I(D_UM_AMIGA_in_6));
    IoInMux I__1233 (
            .O(N__5318),
            .I(N__5315));
    LocalMux I__1232 (
            .O(N__5315),
            .I(N__5312));
    Span12Mux_s4_h I__1231 (
            .O(N__5312),
            .I(N__5309));
    Span12Mux_h I__1230 (
            .O(N__5309),
            .I(N__5306));
    Odrv12 I__1229 (
            .O(N__5306),
            .I(un1_D_UM_AMIGA_6));
    CascadeMux I__1228 (
            .O(N__5303),
            .I(N__5300));
    InMux I__1227 (
            .O(N__5300),
            .I(N__5297));
    LocalMux I__1226 (
            .O(N__5297),
            .I(N__5294));
    Span12Mux_h I__1225 (
            .O(N__5294),
            .I(N__5291));
    Span12Mux_v I__1224 (
            .O(N__5291),
            .I(N__5288));
    Odrv12 I__1223 (
            .O(N__5288),
            .I(TS_CPUn_c));
    InMux I__1222 (
            .O(N__5285),
            .I(N__5282));
    LocalMux I__1221 (
            .O(N__5282),
            .I(N__5270));
    InMux I__1220 (
            .O(N__5281),
            .I(N__5265));
    InMux I__1219 (
            .O(N__5280),
            .I(N__5265));
    InMux I__1218 (
            .O(N__5279),
            .I(N__5254));
    InMux I__1217 (
            .O(N__5278),
            .I(N__5254));
    InMux I__1216 (
            .O(N__5277),
            .I(N__5254));
    InMux I__1215 (
            .O(N__5276),
            .I(N__5254));
    InMux I__1214 (
            .O(N__5275),
            .I(N__5254));
    InMux I__1213 (
            .O(N__5274),
            .I(N__5249));
    InMux I__1212 (
            .O(N__5273),
            .I(N__5249));
    Odrv4 I__1211 (
            .O(N__5270),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1210 (
            .O(N__5265),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1209 (
            .O(N__5254),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1208 (
            .O(N__5249),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    InMux I__1207 (
            .O(N__5240),
            .I(N__5237));
    LocalMux I__1206 (
            .O(N__5237),
            .I(\U111_CYCLE_SM.TS_EN_4 ));
    CEMux I__1205 (
            .O(N__5234),
            .I(N__5227));
    CEMux I__1204 (
            .O(N__5233),
            .I(N__5224));
    CEMux I__1203 (
            .O(N__5232),
            .I(N__5221));
    CEMux I__1202 (
            .O(N__5231),
            .I(N__5218));
    CEMux I__1201 (
            .O(N__5230),
            .I(N__5215));
    LocalMux I__1200 (
            .O(N__5227),
            .I(N__5210));
    LocalMux I__1199 (
            .O(N__5224),
            .I(N__5210));
    LocalMux I__1198 (
            .O(N__5221),
            .I(N__5205));
    LocalMux I__1197 (
            .O(N__5218),
            .I(N__5205));
    LocalMux I__1196 (
            .O(N__5215),
            .I(N__5202));
    Odrv4 I__1195 (
            .O(N__5210),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    Odrv4 I__1194 (
            .O(N__5205),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    Odrv4 I__1193 (
            .O(N__5202),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    SRMux I__1192 (
            .O(N__5195),
            .I(N__5190));
    SRMux I__1191 (
            .O(N__5194),
            .I(N__5185));
    SRMux I__1190 (
            .O(N__5193),
            .I(N__5182));
    LocalMux I__1189 (
            .O(N__5190),
            .I(N__5179));
    SRMux I__1188 (
            .O(N__5189),
            .I(N__5176));
    SRMux I__1187 (
            .O(N__5188),
            .I(N__5173));
    LocalMux I__1186 (
            .O(N__5185),
            .I(N__5170));
    LocalMux I__1185 (
            .O(N__5182),
            .I(N__5167));
    Span4Mux_h I__1184 (
            .O(N__5179),
            .I(N__5162));
    LocalMux I__1183 (
            .O(N__5176),
            .I(N__5162));
    LocalMux I__1182 (
            .O(N__5173),
            .I(N__5159));
    Span4Mux_h I__1181 (
            .O(N__5170),
            .I(N__5154));
    Span4Mux_h I__1180 (
            .O(N__5167),
            .I(N__5154));
    Span4Mux_h I__1179 (
            .O(N__5162),
            .I(N__5149));
    Span4Mux_h I__1178 (
            .O(N__5159),
            .I(N__5149));
    Odrv4 I__1177 (
            .O(N__5154),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0 ));
    Odrv4 I__1176 (
            .O(N__5149),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0 ));
    InMux I__1175 (
            .O(N__5144),
            .I(N__5141));
    LocalMux I__1174 (
            .O(N__5141),
            .I(N__5136));
    InMux I__1173 (
            .O(N__5140),
            .I(N__5133));
    InMux I__1172 (
            .O(N__5139),
            .I(N__5130));
    Span4Mux_v I__1171 (
            .O(N__5136),
            .I(N__5127));
    LocalMux I__1170 (
            .O(N__5133),
            .I(N__5124));
    LocalMux I__1169 (
            .O(N__5130),
            .I(N__5121));
    Span4Mux_v I__1168 (
            .O(N__5127),
            .I(N__5118));
    Span4Mux_v I__1167 (
            .O(N__5124),
            .I(N__5115));
    Span4Mux_h I__1166 (
            .O(N__5121),
            .I(N__5112));
    Sp12to4 I__1165 (
            .O(N__5118),
            .I(N__5109));
    Span4Mux_v I__1164 (
            .O(N__5115),
            .I(N__5106));
    Span4Mux_v I__1163 (
            .O(N__5112),
            .I(N__5103));
    Span12Mux_h I__1162 (
            .O(N__5109),
            .I(N__5100));
    Sp12to4 I__1161 (
            .O(N__5106),
            .I(N__5095));
    Sp12to4 I__1160 (
            .O(N__5103),
            .I(N__5095));
    Span12Mux_v I__1159 (
            .O(N__5100),
            .I(N__5090));
    Span12Mux_h I__1158 (
            .O(N__5095),
            .I(N__5090));
    Odrv12 I__1157 (
            .O(N__5090),
            .I(D_UM_AMIGA_in_3));
    InMux I__1156 (
            .O(N__5087),
            .I(N__5084));
    LocalMux I__1155 (
            .O(N__5084),
            .I(N__5081));
    Odrv12 I__1154 (
            .O(N__5081),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ));
    IoInMux I__1153 (
            .O(N__5078),
            .I(N__5075));
    LocalMux I__1152 (
            .O(N__5075),
            .I(N__5072));
    Span4Mux_s2_h I__1151 (
            .O(N__5072),
            .I(N__5069));
    Span4Mux_h I__1150 (
            .O(N__5069),
            .I(N__5066));
    Sp12to4 I__1149 (
            .O(N__5066),
            .I(N__5063));
    Span12Mux_s9_v I__1148 (
            .O(N__5063),
            .I(N__5060));
    Odrv12 I__1147 (
            .O(N__5060),
            .I(un1_D_UM_AMIGA_3));
    InMux I__1146 (
            .O(N__5057),
            .I(N__5054));
    LocalMux I__1145 (
            .O(N__5054),
            .I(N__5051));
    Odrv12 I__1144 (
            .O(N__5051),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ));
    InMux I__1143 (
            .O(N__5048),
            .I(N__5044));
    InMux I__1142 (
            .O(N__5047),
            .I(N__5041));
    LocalMux I__1141 (
            .O(N__5044),
            .I(N__5037));
    LocalMux I__1140 (
            .O(N__5041),
            .I(N__5034));
    InMux I__1139 (
            .O(N__5040),
            .I(N__5031));
    Span4Mux_v I__1138 (
            .O(N__5037),
            .I(N__5028));
    Span4Mux_h I__1137 (
            .O(N__5034),
            .I(N__5025));
    LocalMux I__1136 (
            .O(N__5031),
            .I(N__5022));
    Sp12to4 I__1135 (
            .O(N__5028),
            .I(N__5019));
    Span4Mux_v I__1134 (
            .O(N__5025),
            .I(N__5014));
    Span4Mux_h I__1133 (
            .O(N__5022),
            .I(N__5014));
    Span12Mux_h I__1132 (
            .O(N__5019),
            .I(N__5011));
    Span4Mux_v I__1131 (
            .O(N__5014),
            .I(N__5008));
    Span12Mux_v I__1130 (
            .O(N__5011),
            .I(N__5005));
    Sp12to4 I__1129 (
            .O(N__5008),
            .I(N__5002));
    Odrv12 I__1128 (
            .O(N__5005),
            .I(D_UM_AMIGA_in_7));
    Odrv12 I__1127 (
            .O(N__5002),
            .I(D_UM_AMIGA_in_7));
    IoInMux I__1126 (
            .O(N__4997),
            .I(N__4994));
    LocalMux I__1125 (
            .O(N__4994),
            .I(N__4991));
    Span4Mux_s1_h I__1124 (
            .O(N__4991),
            .I(N__4988));
    Span4Mux_h I__1123 (
            .O(N__4988),
            .I(N__4985));
    Sp12to4 I__1122 (
            .O(N__4985),
            .I(N__4982));
    Span12Mux_s10_v I__1121 (
            .O(N__4982),
            .I(N__4979));
    Span12Mux_h I__1120 (
            .O(N__4979),
            .I(N__4976));
    Odrv12 I__1119 (
            .O(N__4976),
            .I(un1_D_UM_AMIGA_7));
    InMux I__1118 (
            .O(N__4973),
            .I(N__4970));
    LocalMux I__1117 (
            .O(N__4970),
            .I(N__4967));
    Span4Mux_v I__1116 (
            .O(N__4967),
            .I(N__4964));
    Sp12to4 I__1115 (
            .O(N__4964),
            .I(N__4961));
    Span12Mux_h I__1114 (
            .O(N__4961),
            .I(N__4958));
    Odrv12 I__1113 (
            .O(N__4958),
            .I(D_LL_AMIGA_in_5));
    IoInMux I__1112 (
            .O(N__4955),
            .I(N__4952));
    LocalMux I__1111 (
            .O(N__4952),
            .I(N__4949));
    IoSpan4Mux I__1110 (
            .O(N__4949),
            .I(N__4946));
    Span4Mux_s3_h I__1109 (
            .O(N__4946),
            .I(N__4943));
    Sp12to4 I__1108 (
            .O(N__4943),
            .I(N__4940));
    Span12Mux_h I__1107 (
            .O(N__4940),
            .I(N__4937));
    Odrv12 I__1106 (
            .O(N__4937),
            .I(un1_D_LL_AMIGA_5));
    InMux I__1105 (
            .O(N__4934),
            .I(N__4931));
    LocalMux I__1104 (
            .O(N__4931),
            .I(N__4928));
    Span4Mux_v I__1103 (
            .O(N__4928),
            .I(N__4925));
    Sp12to4 I__1102 (
            .O(N__4925),
            .I(N__4922));
    Span12Mux_h I__1101 (
            .O(N__4922),
            .I(N__4919));
    Odrv12 I__1100 (
            .O(N__4919),
            .I(D_LL_AMIGA_in_7));
    IoInMux I__1099 (
            .O(N__4916),
            .I(N__4913));
    LocalMux I__1098 (
            .O(N__4913),
            .I(N__4910));
    Span4Mux_s2_h I__1097 (
            .O(N__4910),
            .I(N__4907));
    Span4Mux_v I__1096 (
            .O(N__4907),
            .I(N__4904));
    Span4Mux_v I__1095 (
            .O(N__4904),
            .I(N__4901));
    Sp12to4 I__1094 (
            .O(N__4901),
            .I(N__4898));
    Span12Mux_s9_h I__1093 (
            .O(N__4898),
            .I(N__4895));
    Odrv12 I__1092 (
            .O(N__4895),
            .I(un1_D_LL_AMIGA_7));
    InMux I__1091 (
            .O(N__4892),
            .I(N__4889));
    LocalMux I__1090 (
            .O(N__4889),
            .I(N__4886));
    Sp12to4 I__1089 (
            .O(N__4886),
            .I(N__4883));
    Span12Mux_h I__1088 (
            .O(N__4883),
            .I(N__4880));
    Odrv12 I__1087 (
            .O(N__4880),
            .I(D_UM_040_in_2));
    IoInMux I__1086 (
            .O(N__4877),
            .I(N__4874));
    LocalMux I__1085 (
            .O(N__4874),
            .I(N__4870));
    InMux I__1084 (
            .O(N__4873),
            .I(N__4867));
    IoSpan4Mux I__1083 (
            .O(N__4870),
            .I(N__4864));
    LocalMux I__1082 (
            .O(N__4867),
            .I(N__4861));
    Span4Mux_s2_h I__1081 (
            .O(N__4864),
            .I(N__4858));
    Span4Mux_v I__1080 (
            .O(N__4861),
            .I(N__4855));
    Sp12to4 I__1079 (
            .O(N__4858),
            .I(N__4852));
    Sp12to4 I__1078 (
            .O(N__4855),
            .I(N__4849));
    Span12Mux_h I__1077 (
            .O(N__4852),
            .I(N__4846));
    Span12Mux_h I__1076 (
            .O(N__4849),
            .I(N__4843));
    Span12Mux_h I__1075 (
            .O(N__4846),
            .I(N__4838));
    Span12Mux_v I__1074 (
            .O(N__4843),
            .I(N__4838));
    Odrv12 I__1073 (
            .O(N__4838),
            .I(D_LL_040_in_2));
    IoInMux I__1072 (
            .O(N__4835),
            .I(N__4832));
    LocalMux I__1071 (
            .O(N__4832),
            .I(N__4829));
    Span4Mux_s3_h I__1070 (
            .O(N__4829),
            .I(N__4826));
    Span4Mux_v I__1069 (
            .O(N__4826),
            .I(N__4823));
    Sp12to4 I__1068 (
            .O(N__4823),
            .I(N__4820));
    Span12Mux_s10_h I__1067 (
            .O(N__4820),
            .I(N__4817));
    Odrv12 I__1066 (
            .O(N__4817),
            .I(un1_D_UM_040_2));
    IoInMux I__1065 (
            .O(N__4814),
            .I(N__4811));
    LocalMux I__1064 (
            .O(N__4811),
            .I(N__4808));
    Span12Mux_s5_h I__1063 (
            .O(N__4808),
            .I(N__4805));
    Span12Mux_h I__1062 (
            .O(N__4805),
            .I(N__4802));
    Odrv12 I__1061 (
            .O(N__4802),
            .I(un1_D_UM_AMIGA_2));
    InMux I__1060 (
            .O(N__4799),
            .I(N__4794));
    InMux I__1059 (
            .O(N__4798),
            .I(N__4791));
    InMux I__1058 (
            .O(N__4797),
            .I(N__4788));
    LocalMux I__1057 (
            .O(N__4794),
            .I(N__4783));
    LocalMux I__1056 (
            .O(N__4791),
            .I(N__4783));
    LocalMux I__1055 (
            .O(N__4788),
            .I(N__4780));
    Span4Mux_v I__1054 (
            .O(N__4783),
            .I(N__4777));
    Sp12to4 I__1053 (
            .O(N__4780),
            .I(N__4774));
    Sp12to4 I__1052 (
            .O(N__4777),
            .I(N__4771));
    Span12Mux_v I__1051 (
            .O(N__4774),
            .I(N__4768));
    Span12Mux_h I__1050 (
            .O(N__4771),
            .I(N__4765));
    Odrv12 I__1049 (
            .O(N__4768),
            .I(D_UM_AMIGA_in_2));
    Odrv12 I__1048 (
            .O(N__4765),
            .I(D_UM_AMIGA_in_2));
    InMux I__1047 (
            .O(N__4760),
            .I(N__4757));
    LocalMux I__1046 (
            .O(N__4757),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ));
    CascadeMux I__1045 (
            .O(N__4754),
            .I(N__4749));
    CascadeMux I__1044 (
            .O(N__4753),
            .I(N__4743));
    CascadeMux I__1043 (
            .O(N__4752),
            .I(N__4739));
    InMux I__1042 (
            .O(N__4749),
            .I(N__4735));
    InMux I__1041 (
            .O(N__4748),
            .I(N__4730));
    InMux I__1040 (
            .O(N__4747),
            .I(N__4730));
    InMux I__1039 (
            .O(N__4746),
            .I(N__4723));
    InMux I__1038 (
            .O(N__4743),
            .I(N__4723));
    InMux I__1037 (
            .O(N__4742),
            .I(N__4723));
    InMux I__1036 (
            .O(N__4739),
            .I(N__4720));
    InMux I__1035 (
            .O(N__4738),
            .I(N__4717));
    LocalMux I__1034 (
            .O(N__4735),
            .I(N__4706));
    LocalMux I__1033 (
            .O(N__4730),
            .I(N__4706));
    LocalMux I__1032 (
            .O(N__4723),
            .I(N__4706));
    LocalMux I__1031 (
            .O(N__4720),
            .I(N__4706));
    LocalMux I__1030 (
            .O(N__4717),
            .I(N__4706));
    Span4Mux_v I__1029 (
            .O(N__4706),
            .I(N__4703));
    Span4Mux_h I__1028 (
            .O(N__4703),
            .I(N__4699));
    InMux I__1027 (
            .O(N__4702),
            .I(N__4696));
    Sp12to4 I__1026 (
            .O(N__4699),
            .I(N__4693));
    LocalMux I__1025 (
            .O(N__4696),
            .I(N__4690));
    Span12Mux_s11_h I__1024 (
            .O(N__4693),
            .I(N__4685));
    Span12Mux_v I__1023 (
            .O(N__4690),
            .I(N__4685));
    Span12Mux_v I__1022 (
            .O(N__4685),
            .I(N__4682));
    Odrv12 I__1021 (
            .O(N__4682),
            .I(RESETn_c));
    InMux I__1020 (
            .O(N__4679),
            .I(N__4676));
    LocalMux I__1019 (
            .O(N__4676),
            .I(N__4673));
    Odrv4 I__1018 (
            .O(N__4673),
            .I(\U111_CYCLE_SM.TA_ENZ0 ));
    InMux I__1017 (
            .O(N__4670),
            .I(N__4661));
    InMux I__1016 (
            .O(N__4669),
            .I(N__4661));
    InMux I__1015 (
            .O(N__4668),
            .I(N__4658));
    InMux I__1014 (
            .O(N__4667),
            .I(N__4653));
    InMux I__1013 (
            .O(N__4666),
            .I(N__4653));
    LocalMux I__1012 (
            .O(N__4661),
            .I(N__4648));
    LocalMux I__1011 (
            .O(N__4658),
            .I(N__4648));
    LocalMux I__1010 (
            .O(N__4653),
            .I(N__4645));
    Sp12to4 I__1009 (
            .O(N__4648),
            .I(N__4640));
    Sp12to4 I__1008 (
            .O(N__4645),
            .I(N__4640));
    Span12Mux_v I__1007 (
            .O(N__4640),
            .I(N__4637));
    Odrv12 I__1006 (
            .O(N__4637),
            .I(TACKn_c));
    IoInMux I__1005 (
            .O(N__4634),
            .I(N__4631));
    LocalMux I__1004 (
            .O(N__4631),
            .I(N__4628));
    Span4Mux_s3_v I__1003 (
            .O(N__4628),
            .I(N__4625));
    Sp12to4 I__1002 (
            .O(N__4625),
            .I(N__4622));
    Span12Mux_h I__1001 (
            .O(N__4622),
            .I(N__4619));
    Odrv12 I__1000 (
            .O(N__4619),
            .I(TAn_0_i));
    CascadeMux I__999 (
            .O(N__4616),
            .I(N__4609));
    CascadeMux I__998 (
            .O(N__4615),
            .I(N__4606));
    CascadeMux I__997 (
            .O(N__4614),
            .I(N__4602));
    InMux I__996 (
            .O(N__4613),
            .I(N__4598));
    InMux I__995 (
            .O(N__4612),
            .I(N__4595));
    InMux I__994 (
            .O(N__4609),
            .I(N__4588));
    InMux I__993 (
            .O(N__4606),
            .I(N__4588));
    InMux I__992 (
            .O(N__4605),
            .I(N__4588));
    InMux I__991 (
            .O(N__4602),
            .I(N__4583));
    InMux I__990 (
            .O(N__4601),
            .I(N__4583));
    LocalMux I__989 (
            .O(N__4598),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__988 (
            .O(N__4595),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__987 (
            .O(N__4588),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__986 (
            .O(N__4583),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    InMux I__985 (
            .O(N__4574),
            .I(N__4571));
    LocalMux I__984 (
            .O(N__4571),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ));
    InMux I__983 (
            .O(N__4568),
            .I(N__4565));
    LocalMux I__982 (
            .O(N__4565),
            .I(N__4561));
    InMux I__981 (
            .O(N__4564),
            .I(N__4558));
    Span4Mux_v I__980 (
            .O(N__4561),
            .I(N__4554));
    LocalMux I__979 (
            .O(N__4558),
            .I(N__4551));
    InMux I__978 (
            .O(N__4557),
            .I(N__4548));
    Sp12to4 I__977 (
            .O(N__4554),
            .I(N__4545));
    Span4Mux_v I__976 (
            .O(N__4551),
            .I(N__4542));
    LocalMux I__975 (
            .O(N__4548),
            .I(N__4539));
    Span12Mux_h I__974 (
            .O(N__4545),
            .I(N__4536));
    Sp12to4 I__973 (
            .O(N__4542),
            .I(N__4531));
    Span12Mux_v I__972 (
            .O(N__4539),
            .I(N__4531));
    Span12Mux_v I__971 (
            .O(N__4536),
            .I(N__4528));
    Span12Mux_h I__970 (
            .O(N__4531),
            .I(N__4525));
    Odrv12 I__969 (
            .O(N__4528),
            .I(D_UM_AMIGA_in_1));
    Odrv12 I__968 (
            .O(N__4525),
            .I(D_UM_AMIGA_in_1));
    IoInMux I__967 (
            .O(N__4520),
            .I(N__4517));
    LocalMux I__966 (
            .O(N__4517),
            .I(N__4514));
    Span4Mux_s2_h I__965 (
            .O(N__4514),
            .I(N__4511));
    Sp12to4 I__964 (
            .O(N__4511),
            .I(N__4508));
    Span12Mux_s11_v I__963 (
            .O(N__4508),
            .I(N__4505));
    Span12Mux_h I__962 (
            .O(N__4505),
            .I(N__4502));
    Odrv12 I__961 (
            .O(N__4502),
            .I(un1_D_UM_AMIGA_1));
    InMux I__960 (
            .O(N__4499),
            .I(N__4496));
    LocalMux I__959 (
            .O(N__4496),
            .I(N__4492));
    InMux I__958 (
            .O(N__4495),
            .I(N__4489));
    Span4Mux_v I__957 (
            .O(N__4492),
            .I(N__4483));
    LocalMux I__956 (
            .O(N__4489),
            .I(N__4483));
    InMux I__955 (
            .O(N__4488),
            .I(N__4480));
    Span4Mux_v I__954 (
            .O(N__4483),
            .I(N__4475));
    LocalMux I__953 (
            .O(N__4480),
            .I(N__4475));
    Span4Mux_h I__952 (
            .O(N__4475),
            .I(N__4472));
    Span4Mux_v I__951 (
            .O(N__4472),
            .I(N__4469));
    Sp12to4 I__950 (
            .O(N__4469),
            .I(N__4466));
    Odrv12 I__949 (
            .O(N__4466),
            .I(D_UU_AMIGA_in_1));
    InMux I__948 (
            .O(N__4463),
            .I(N__4460));
    LocalMux I__947 (
            .O(N__4460),
            .I(N__4457));
    Odrv4 I__946 (
            .O(N__4457),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ));
    IoInMux I__945 (
            .O(N__4454),
            .I(N__4451));
    LocalMux I__944 (
            .O(N__4451),
            .I(N__4448));
    IoSpan4Mux I__943 (
            .O(N__4448),
            .I(N__4445));
    IoSpan4Mux I__942 (
            .O(N__4445),
            .I(N__4442));
    Sp12to4 I__941 (
            .O(N__4442),
            .I(N__4439));
    Span12Mux_s9_h I__940 (
            .O(N__4439),
            .I(N__4436));
    Odrv12 I__939 (
            .O(N__4436),
            .I(un1_D_UU_AMIGA_1));
    InMux I__938 (
            .O(N__4433),
            .I(N__4430));
    LocalMux I__937 (
            .O(N__4430),
            .I(N__4427));
    Odrv12 I__936 (
            .O(N__4427),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ));
    InMux I__935 (
            .O(N__4424),
            .I(N__4420));
    InMux I__934 (
            .O(N__4423),
            .I(N__4416));
    LocalMux I__933 (
            .O(N__4420),
            .I(N__4413));
    InMux I__932 (
            .O(N__4419),
            .I(N__4410));
    LocalMux I__931 (
            .O(N__4416),
            .I(N__4407));
    Span4Mux_h I__930 (
            .O(N__4413),
            .I(N__4404));
    LocalMux I__929 (
            .O(N__4410),
            .I(N__4401));
    Span12Mux_v I__928 (
            .O(N__4407),
            .I(N__4398));
    Span4Mux_v I__927 (
            .O(N__4404),
            .I(N__4393));
    Span4Mux_h I__926 (
            .O(N__4401),
            .I(N__4393));
    Span12Mux_h I__925 (
            .O(N__4398),
            .I(N__4390));
    Span4Mux_v I__924 (
            .O(N__4393),
            .I(N__4387));
    Span12Mux_v I__923 (
            .O(N__4390),
            .I(N__4384));
    Sp12to4 I__922 (
            .O(N__4387),
            .I(N__4381));
    Odrv12 I__921 (
            .O(N__4384),
            .I(D_UM_AMIGA_in_4));
    Odrv12 I__920 (
            .O(N__4381),
            .I(D_UM_AMIGA_in_4));
    IoInMux I__919 (
            .O(N__4376),
            .I(N__4373));
    LocalMux I__918 (
            .O(N__4373),
            .I(N__4370));
    Span4Mux_s0_v I__917 (
            .O(N__4370),
            .I(N__4367));
    Span4Mux_v I__916 (
            .O(N__4367),
            .I(N__4364));
    Span4Mux_v I__915 (
            .O(N__4364),
            .I(N__4361));
    Sp12to4 I__914 (
            .O(N__4361),
            .I(N__4358));
    Span12Mux_s11_h I__913 (
            .O(N__4358),
            .I(N__4355));
    Odrv12 I__912 (
            .O(N__4355),
            .I(un1_D_UM_AMIGA_4));
    InMux I__911 (
            .O(N__4352),
            .I(N__4349));
    LocalMux I__910 (
            .O(N__4349),
            .I(N__4346));
    Span4Mux_v I__909 (
            .O(N__4346),
            .I(N__4343));
    Sp12to4 I__908 (
            .O(N__4343),
            .I(N__4340));
    Span12Mux_h I__907 (
            .O(N__4340),
            .I(N__4337));
    Odrv12 I__906 (
            .O(N__4337),
            .I(D_UU_040_in_0));
    IoInMux I__905 (
            .O(N__4334),
            .I(N__4331));
    LocalMux I__904 (
            .O(N__4331),
            .I(N__4328));
    IoSpan4Mux I__903 (
            .O(N__4328),
            .I(N__4324));
    InMux I__902 (
            .O(N__4327),
            .I(N__4321));
    IoSpan4Mux I__901 (
            .O(N__4324),
            .I(N__4318));
    LocalMux I__900 (
            .O(N__4321),
            .I(N__4315));
    Span4Mux_s2_h I__899 (
            .O(N__4318),
            .I(N__4312));
    Span12Mux_v I__898 (
            .O(N__4315),
            .I(N__4309));
    Sp12to4 I__897 (
            .O(N__4312),
            .I(N__4306));
    Span12Mux_h I__896 (
            .O(N__4309),
            .I(N__4303));
    Span12Mux_h I__895 (
            .O(N__4306),
            .I(N__4300));
    Span12Mux_v I__894 (
            .O(N__4303),
            .I(N__4295));
    Span12Mux_h I__893 (
            .O(N__4300),
            .I(N__4295));
    Odrv12 I__892 (
            .O(N__4295),
            .I(D_LM_040_in_0));
    IoInMux I__891 (
            .O(N__4292),
            .I(N__4289));
    LocalMux I__890 (
            .O(N__4289),
            .I(N__4286));
    IoSpan4Mux I__889 (
            .O(N__4286),
            .I(N__4283));
    Sp12to4 I__888 (
            .O(N__4283),
            .I(N__4280));
    Span12Mux_s6_v I__887 (
            .O(N__4280),
            .I(N__4277));
    Odrv12 I__886 (
            .O(N__4277),
            .I(un1_D_UU_040_0));
    InMux I__885 (
            .O(N__4274),
            .I(N__4271));
    LocalMux I__884 (
            .O(N__4271),
            .I(N__4268));
    Sp12to4 I__883 (
            .O(N__4268),
            .I(N__4265));
    Span12Mux_s7_v I__882 (
            .O(N__4265),
            .I(N__4262));
    Span12Mux_h I__881 (
            .O(N__4262),
            .I(N__4259));
    Odrv12 I__880 (
            .O(N__4259),
            .I(D_UU_040_in_2));
    IoInMux I__879 (
            .O(N__4256),
            .I(N__4252));
    InMux I__878 (
            .O(N__4255),
            .I(N__4249));
    LocalMux I__877 (
            .O(N__4252),
            .I(N__4246));
    LocalMux I__876 (
            .O(N__4249),
            .I(N__4243));
    Span12Mux_s9_h I__875 (
            .O(N__4246),
            .I(N__4240));
    Span12Mux_v I__874 (
            .O(N__4243),
            .I(N__4237));
    Span12Mux_v I__873 (
            .O(N__4240),
            .I(N__4234));
    Span12Mux_h I__872 (
            .O(N__4237),
            .I(N__4231));
    Span12Mux_h I__871 (
            .O(N__4234),
            .I(N__4228));
    Span12Mux_v I__870 (
            .O(N__4231),
            .I(N__4225));
    Odrv12 I__869 (
            .O(N__4228),
            .I(D_LM_040_in_2));
    Odrv12 I__868 (
            .O(N__4225),
            .I(D_LM_040_in_2));
    IoInMux I__867 (
            .O(N__4220),
            .I(N__4217));
    LocalMux I__866 (
            .O(N__4217),
            .I(N__4214));
    IoSpan4Mux I__865 (
            .O(N__4214),
            .I(N__4211));
    IoSpan4Mux I__864 (
            .O(N__4211),
            .I(N__4208));
    Span4Mux_s3_v I__863 (
            .O(N__4208),
            .I(N__4205));
    Odrv4 I__862 (
            .O(N__4205),
            .I(un1_D_UU_040_2));
    InMux I__861 (
            .O(N__4202),
            .I(N__4199));
    LocalMux I__860 (
            .O(N__4199),
            .I(N__4196));
    Span4Mux_v I__859 (
            .O(N__4196),
            .I(N__4193));
    Odrv4 I__858 (
            .O(N__4193),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ));
    InMux I__857 (
            .O(N__4190),
            .I(N__4187));
    LocalMux I__856 (
            .O(N__4187),
            .I(N__4184));
    Span4Mux_h I__855 (
            .O(N__4184),
            .I(N__4180));
    InMux I__854 (
            .O(N__4183),
            .I(N__4177));
    Span4Mux_v I__853 (
            .O(N__4180),
            .I(N__4172));
    LocalMux I__852 (
            .O(N__4177),
            .I(N__4172));
    Span4Mux_v I__851 (
            .O(N__4172),
            .I(N__4168));
    InMux I__850 (
            .O(N__4171),
            .I(N__4165));
    Span4Mux_v I__849 (
            .O(N__4168),
            .I(N__4160));
    LocalMux I__848 (
            .O(N__4165),
            .I(N__4160));
    Span4Mux_v I__847 (
            .O(N__4160),
            .I(N__4157));
    Span4Mux_h I__846 (
            .O(N__4157),
            .I(N__4154));
    Span4Mux_h I__845 (
            .O(N__4154),
            .I(N__4151));
    Odrv4 I__844 (
            .O(N__4151),
            .I(D_UU_AMIGA_in_0));
    IoInMux I__843 (
            .O(N__4148),
            .I(N__4145));
    LocalMux I__842 (
            .O(N__4145),
            .I(N__4142));
    IoSpan4Mux I__841 (
            .O(N__4142),
            .I(N__4139));
    Span4Mux_s2_v I__840 (
            .O(N__4139),
            .I(N__4136));
    Span4Mux_v I__839 (
            .O(N__4136),
            .I(N__4133));
    Sp12to4 I__838 (
            .O(N__4133),
            .I(N__4130));
    Odrv12 I__837 (
            .O(N__4130),
            .I(un1_D_UU_AMIGA_0));
    InMux I__836 (
            .O(N__4127),
            .I(N__4124));
    LocalMux I__835 (
            .O(N__4124),
            .I(N__4121));
    Span4Mux_v I__834 (
            .O(N__4121),
            .I(N__4118));
    Sp12to4 I__833 (
            .O(N__4118),
            .I(N__4115));
    Span12Mux_h I__832 (
            .O(N__4115),
            .I(N__4112));
    Odrv12 I__831 (
            .O(N__4112),
            .I(D_LL_AMIGA_in_6));
    IoInMux I__830 (
            .O(N__4109),
            .I(N__4106));
    LocalMux I__829 (
            .O(N__4106),
            .I(N__4103));
    Span4Mux_s2_h I__828 (
            .O(N__4103),
            .I(N__4100));
    Span4Mux_v I__827 (
            .O(N__4100),
            .I(N__4097));
    Span4Mux_v I__826 (
            .O(N__4097),
            .I(N__4094));
    Sp12to4 I__825 (
            .O(N__4094),
            .I(N__4091));
    Span12Mux_s9_h I__824 (
            .O(N__4091),
            .I(N__4088));
    Odrv12 I__823 (
            .O(N__4088),
            .I(un1_D_LL_AMIGA_6));
    InMux I__822 (
            .O(N__4085),
            .I(N__4082));
    LocalMux I__821 (
            .O(N__4082),
            .I(\U111_CYCLE_SM.TS_EN10 ));
    CascadeMux I__820 (
            .O(N__4079),
            .I(N__4076));
    InMux I__819 (
            .O(N__4076),
            .I(N__4072));
    InMux I__818 (
            .O(N__4075),
            .I(N__4069));
    LocalMux I__817 (
            .O(N__4072),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    LocalMux I__816 (
            .O(N__4069),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    IoInMux I__815 (
            .O(N__4064),
            .I(N__4061));
    LocalMux I__814 (
            .O(N__4061),
            .I(N__4058));
    IoSpan4Mux I__813 (
            .O(N__4058),
            .I(N__4055));
    Span4Mux_s2_v I__812 (
            .O(N__4055),
            .I(N__4052));
    Sp12to4 I__811 (
            .O(N__4052),
            .I(N__4048));
    InMux I__810 (
            .O(N__4051),
            .I(N__4045));
    Odrv12 I__809 (
            .O(N__4048),
            .I(TSn_c));
    LocalMux I__808 (
            .O(N__4045),
            .I(TSn_c));
    CascadeMux I__807 (
            .O(N__4040),
            .I(N__4036));
    InMux I__806 (
            .O(N__4039),
            .I(N__4031));
    InMux I__805 (
            .O(N__4036),
            .I(N__4031));
    LocalMux I__804 (
            .O(N__4031),
            .I(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ));
    IoInMux I__803 (
            .O(N__4028),
            .I(N__4024));
    IoInMux I__802 (
            .O(N__4027),
            .I(N__4021));
    LocalMux I__801 (
            .O(N__4024),
            .I(N__4014));
    LocalMux I__800 (
            .O(N__4021),
            .I(N__4014));
    IoInMux I__799 (
            .O(N__4020),
            .I(N__4011));
    IoInMux I__798 (
            .O(N__4019),
            .I(N__4008));
    IoSpan4Mux I__797 (
            .O(N__4014),
            .I(N__3994));
    LocalMux I__796 (
            .O(N__4011),
            .I(N__3994));
    LocalMux I__795 (
            .O(N__4008),
            .I(N__3994));
    IoInMux I__794 (
            .O(N__4007),
            .I(N__3991));
    IoInMux I__793 (
            .O(N__4006),
            .I(N__3988));
    IoInMux I__792 (
            .O(N__4005),
            .I(N__3985));
    IoInMux I__791 (
            .O(N__4004),
            .I(N__3982));
    IoInMux I__790 (
            .O(N__4003),
            .I(N__3979));
    IoInMux I__789 (
            .O(N__4002),
            .I(N__3974));
    InMux I__788 (
            .O(N__4001),
            .I(N__3971));
    IoSpan4Mux I__787 (
            .O(N__3994),
            .I(N__3956));
    LocalMux I__786 (
            .O(N__3991),
            .I(N__3956));
    LocalMux I__785 (
            .O(N__3988),
            .I(N__3956));
    LocalMux I__784 (
            .O(N__3985),
            .I(N__3956));
    LocalMux I__783 (
            .O(N__3982),
            .I(N__3956));
    LocalMux I__782 (
            .O(N__3979),
            .I(N__3956));
    IoInMux I__781 (
            .O(N__3978),
            .I(N__3953));
    IoInMux I__780 (
            .O(N__3977),
            .I(N__3950));
    LocalMux I__779 (
            .O(N__3974),
            .I(N__3947));
    LocalMux I__778 (
            .O(N__3971),
            .I(N__3944));
    IoInMux I__777 (
            .O(N__3970),
            .I(N__3940));
    IoInMux I__776 (
            .O(N__3969),
            .I(N__3937));
    IoSpan4Mux I__775 (
            .O(N__3956),
            .I(N__3924));
    LocalMux I__774 (
            .O(N__3953),
            .I(N__3924));
    LocalMux I__773 (
            .O(N__3950),
            .I(N__3924));
    Span4Mux_s3_v I__772 (
            .O(N__3947),
            .I(N__3920));
    Span4Mux_h I__771 (
            .O(N__3944),
            .I(N__3917));
    InMux I__770 (
            .O(N__3943),
            .I(N__3914));
    LocalMux I__769 (
            .O(N__3940),
            .I(N__3909));
    LocalMux I__768 (
            .O(N__3937),
            .I(N__3909));
    IoInMux I__767 (
            .O(N__3936),
            .I(N__3906));
    IoInMux I__766 (
            .O(N__3935),
            .I(N__3903));
    IoInMux I__765 (
            .O(N__3934),
            .I(N__3900));
    IoInMux I__764 (
            .O(N__3933),
            .I(N__3897));
    IoInMux I__763 (
            .O(N__3932),
            .I(N__3894));
    IoInMux I__762 (
            .O(N__3931),
            .I(N__3891));
    IoSpan4Mux I__761 (
            .O(N__3924),
            .I(N__3884));
    IoInMux I__760 (
            .O(N__3923),
            .I(N__3881));
    Span4Mux_v I__759 (
            .O(N__3920),
            .I(N__3877));
    Span4Mux_h I__758 (
            .O(N__3917),
            .I(N__3872));
    LocalMux I__757 (
            .O(N__3914),
            .I(N__3872));
    IoSpan4Mux I__756 (
            .O(N__3909),
            .I(N__3856));
    LocalMux I__755 (
            .O(N__3906),
            .I(N__3856));
    LocalMux I__754 (
            .O(N__3903),
            .I(N__3856));
    LocalMux I__753 (
            .O(N__3900),
            .I(N__3856));
    LocalMux I__752 (
            .O(N__3897),
            .I(N__3856));
    LocalMux I__751 (
            .O(N__3894),
            .I(N__3856));
    LocalMux I__750 (
            .O(N__3891),
            .I(N__3856));
    IoInMux I__749 (
            .O(N__3890),
            .I(N__3853));
    IoInMux I__748 (
            .O(N__3889),
            .I(N__3850));
    IoInMux I__747 (
            .O(N__3888),
            .I(N__3847));
    IoInMux I__746 (
            .O(N__3887),
            .I(N__3844));
    IoSpan4Mux I__745 (
            .O(N__3884),
            .I(N__3839));
    LocalMux I__744 (
            .O(N__3881),
            .I(N__3839));
    IoInMux I__743 (
            .O(N__3880),
            .I(N__3836));
    Span4Mux_v I__742 (
            .O(N__3877),
            .I(N__3830));
    Span4Mux_v I__741 (
            .O(N__3872),
            .I(N__3827));
    IoInMux I__740 (
            .O(N__3871),
            .I(N__3824));
    IoSpan4Mux I__739 (
            .O(N__3856),
            .I(N__3813));
    LocalMux I__738 (
            .O(N__3853),
            .I(N__3813));
    LocalMux I__737 (
            .O(N__3850),
            .I(N__3813));
    LocalMux I__736 (
            .O(N__3847),
            .I(N__3813));
    LocalMux I__735 (
            .O(N__3844),
            .I(N__3813));
    IoSpan4Mux I__734 (
            .O(N__3839),
            .I(N__3809));
    LocalMux I__733 (
            .O(N__3836),
            .I(N__3806));
    IoInMux I__732 (
            .O(N__3835),
            .I(N__3803));
    IoInMux I__731 (
            .O(N__3834),
            .I(N__3800));
    IoInMux I__730 (
            .O(N__3833),
            .I(N__3797));
    Sp12to4 I__729 (
            .O(N__3830),
            .I(N__3793));
    Sp12to4 I__728 (
            .O(N__3827),
            .I(N__3789));
    LocalMux I__727 (
            .O(N__3824),
            .I(N__3786));
    IoSpan4Mux I__726 (
            .O(N__3813),
            .I(N__3783));
    IoInMux I__725 (
            .O(N__3812),
            .I(N__3780));
    IoSpan4Mux I__724 (
            .O(N__3809),
            .I(N__3769));
    IoSpan4Mux I__723 (
            .O(N__3806),
            .I(N__3769));
    LocalMux I__722 (
            .O(N__3803),
            .I(N__3769));
    LocalMux I__721 (
            .O(N__3800),
            .I(N__3769));
    LocalMux I__720 (
            .O(N__3797),
            .I(N__3769));
    IoInMux I__719 (
            .O(N__3796),
            .I(N__3766));
    Span12Mux_h I__718 (
            .O(N__3793),
            .I(N__3763));
    IoInMux I__717 (
            .O(N__3792),
            .I(N__3760));
    Span12Mux_h I__716 (
            .O(N__3789),
            .I(N__3755));
    Span12Mux_s11_v I__715 (
            .O(N__3786),
            .I(N__3755));
    IoSpan4Mux I__714 (
            .O(N__3783),
            .I(N__3750));
    LocalMux I__713 (
            .O(N__3780),
            .I(N__3750));
    IoSpan4Mux I__712 (
            .O(N__3769),
            .I(N__3745));
    LocalMux I__711 (
            .O(N__3766),
            .I(N__3745));
    Span12Mux_h I__710 (
            .O(N__3763),
            .I(N__3740));
    LocalMux I__709 (
            .O(N__3760),
            .I(N__3740));
    Odrv12 I__708 (
            .O(N__3755),
            .I(RnW_c));
    Odrv4 I__707 (
            .O(N__3750),
            .I(RnW_c));
    Odrv4 I__706 (
            .O(N__3745),
            .I(RnW_c));
    Odrv12 I__705 (
            .O(N__3740),
            .I(RnW_c));
    CascadeMux I__704 (
            .O(N__3731),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_ ));
    CascadeMux I__703 (
            .O(N__3728),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_ ));
    InMux I__702 (
            .O(N__3725),
            .I(N__3722));
    LocalMux I__701 (
            .O(N__3722),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa ));
    InMux I__700 (
            .O(N__3719),
            .I(N__3716));
    LocalMux I__699 (
            .O(N__3716),
            .I(N__3713));
    Span12Mux_v I__698 (
            .O(N__3713),
            .I(N__3710));
    Span12Mux_h I__697 (
            .O(N__3710),
            .I(N__3707));
    Odrv12 I__696 (
            .O(N__3707),
            .I(D_LM_AMIGA_in_0));
    IoInMux I__695 (
            .O(N__3704),
            .I(N__3701));
    LocalMux I__694 (
            .O(N__3701),
            .I(N__3698));
    Span4Mux_s3_h I__693 (
            .O(N__3698),
            .I(N__3695));
    Span4Mux_v I__692 (
            .O(N__3695),
            .I(N__3692));
    Span4Mux_v I__691 (
            .O(N__3692),
            .I(N__3689));
    Span4Mux_h I__690 (
            .O(N__3689),
            .I(N__3686));
    Sp12to4 I__689 (
            .O(N__3686),
            .I(N__3683));
    Odrv12 I__688 (
            .O(N__3683),
            .I(un1_D_LM_AMIGA_0));
    InMux I__687 (
            .O(N__3680),
            .I(N__3677));
    LocalMux I__686 (
            .O(N__3677),
            .I(N__3674));
    Span12Mux_h I__685 (
            .O(N__3674),
            .I(N__3671));
    Odrv12 I__684 (
            .O(N__3671),
            .I(D_LM_AMIGA_in_1));
    IoInMux I__683 (
            .O(N__3668),
            .I(N__3665));
    LocalMux I__682 (
            .O(N__3665),
            .I(N__3662));
    Span4Mux_s0_h I__681 (
            .O(N__3662),
            .I(N__3659));
    Span4Mux_h I__680 (
            .O(N__3659),
            .I(N__3656));
    Span4Mux_h I__679 (
            .O(N__3656),
            .I(N__3653));
    Sp12to4 I__678 (
            .O(N__3653),
            .I(N__3650));
    Span12Mux_v I__677 (
            .O(N__3650),
            .I(N__3647));
    Odrv12 I__676 (
            .O(N__3647),
            .I(un1_D_LM_AMIGA_1));
    InMux I__675 (
            .O(N__3644),
            .I(N__3641));
    LocalMux I__674 (
            .O(N__3641),
            .I(N__3638));
    Span4Mux_v I__673 (
            .O(N__3638),
            .I(N__3635));
    Sp12to4 I__672 (
            .O(N__3635),
            .I(N__3632));
    Span12Mux_h I__671 (
            .O(N__3632),
            .I(N__3628));
    InMux I__670 (
            .O(N__3631),
            .I(N__3625));
    Odrv12 I__669 (
            .O(N__3628),
            .I(\U111_CYCLE_SM.A_OUTZ0 ));
    LocalMux I__668 (
            .O(N__3625),
            .I(\U111_CYCLE_SM.A_OUTZ0 ));
    CascadeMux I__667 (
            .O(N__3620),
            .I(\U111_CYCLE_SM.LW_CYCLE_r_1_cascade_ ));
    InMux I__666 (
            .O(N__3617),
            .I(N__3614));
    LocalMux I__665 (
            .O(N__3614),
            .I(\U111_CYCLE_SM.un1_CYCLE_STATE_1_0 ));
    CascadeMux I__664 (
            .O(N__3611),
            .I(\U111_CYCLE_SM.un1_CYCLE_STATE_1_0_cascade_ ));
    InMux I__663 (
            .O(N__3608),
            .I(N__3604));
    SRMux I__662 (
            .O(N__3607),
            .I(N__3601));
    LocalMux I__661 (
            .O(N__3604),
            .I(N__3598));
    LocalMux I__660 (
            .O(N__3601),
            .I(RESETn_c_i));
    Odrv12 I__659 (
            .O(N__3598),
            .I(RESETn_c_i));
    CEMux I__658 (
            .O(N__3593),
            .I(N__3590));
    LocalMux I__657 (
            .O(N__3590),
            .I(N__3587));
    Span4Mux_v I__656 (
            .O(N__3587),
            .I(N__3584));
    Odrv4 I__655 (
            .O(N__3584),
            .I(\U111_CYCLE_SM.un1_CYCLE_STATE_1_0_0 ));
    InMux I__654 (
            .O(N__3581),
            .I(N__3577));
    IoInMux I__653 (
            .O(N__3580),
            .I(N__3574));
    LocalMux I__652 (
            .O(N__3577),
            .I(N__3571));
    LocalMux I__651 (
            .O(N__3574),
            .I(N__3568));
    Span4Mux_h I__650 (
            .O(N__3571),
            .I(N__3565));
    Span4Mux_s3_h I__649 (
            .O(N__3568),
            .I(N__3562));
    Span4Mux_h I__648 (
            .O(N__3565),
            .I(N__3559));
    Sp12to4 I__647 (
            .O(N__3562),
            .I(N__3556));
    Sp12to4 I__646 (
            .O(N__3559),
            .I(N__3553));
    Span12Mux_v I__645 (
            .O(N__3556),
            .I(N__3550));
    Span12Mux_v I__644 (
            .O(N__3553),
            .I(N__3547));
    Span12Mux_h I__643 (
            .O(N__3550),
            .I(N__3544));
    Span12Mux_v I__642 (
            .O(N__3547),
            .I(N__3541));
    Span12Mux_h I__641 (
            .O(N__3544),
            .I(N__3538));
    Span12Mux_h I__640 (
            .O(N__3541),
            .I(N__3535));
    Odrv12 I__639 (
            .O(N__3538),
            .I(D_LM_040_in_1));
    Odrv12 I__638 (
            .O(N__3535),
            .I(D_LM_040_in_1));
    InMux I__637 (
            .O(N__3530),
            .I(N__3527));
    LocalMux I__636 (
            .O(N__3527),
            .I(N__3524));
    Span4Mux_v I__635 (
            .O(N__3524),
            .I(N__3521));
    Span4Mux_v I__634 (
            .O(N__3521),
            .I(N__3518));
    Sp12to4 I__633 (
            .O(N__3518),
            .I(N__3515));
    Span12Mux_h I__632 (
            .O(N__3515),
            .I(N__3512));
    Odrv12 I__631 (
            .O(N__3512),
            .I(D_UU_040_in_1));
    IoInMux I__630 (
            .O(N__3509),
            .I(N__3506));
    LocalMux I__629 (
            .O(N__3506),
            .I(N__3503));
    Span4Mux_s3_h I__628 (
            .O(N__3503),
            .I(N__3500));
    Sp12to4 I__627 (
            .O(N__3500),
            .I(N__3497));
    Span12Mux_s8_v I__626 (
            .O(N__3497),
            .I(N__3494));
    Odrv12 I__625 (
            .O(N__3494),
            .I(un1_D_UU_040_1));
    InMux I__624 (
            .O(N__3491),
            .I(N__3487));
    InMux I__623 (
            .O(N__3490),
            .I(N__3484));
    LocalMux I__622 (
            .O(N__3487),
            .I(N__3481));
    LocalMux I__621 (
            .O(N__3484),
            .I(N__3478));
    Span4Mux_v I__620 (
            .O(N__3481),
            .I(N__3472));
    Span4Mux_v I__619 (
            .O(N__3478),
            .I(N__3472));
    InMux I__618 (
            .O(N__3477),
            .I(N__3469));
    Sp12to4 I__617 (
            .O(N__3472),
            .I(N__3464));
    LocalMux I__616 (
            .O(N__3469),
            .I(N__3464));
    Span12Mux_h I__615 (
            .O(N__3464),
            .I(N__3461));
    Odrv12 I__614 (
            .O(N__3461),
            .I(D_UU_AMIGA_in_6));
    InMux I__613 (
            .O(N__3458),
            .I(N__3455));
    LocalMux I__612 (
            .O(N__3455),
            .I(N__3452));
    Odrv12 I__611 (
            .O(N__3452),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ));
    IoInMux I__610 (
            .O(N__3449),
            .I(N__3446));
    LocalMux I__609 (
            .O(N__3446),
            .I(N__3443));
    Span4Mux_s3_v I__608 (
            .O(N__3443),
            .I(N__3440));
    Span4Mux_h I__607 (
            .O(N__3440),
            .I(N__3437));
    Span4Mux_h I__606 (
            .O(N__3437),
            .I(N__3434));
    Span4Mux_h I__605 (
            .O(N__3434),
            .I(N__3431));
    Span4Mux_v I__604 (
            .O(N__3431),
            .I(N__3428));
    Odrv4 I__603 (
            .O(N__3428),
            .I(un1_D_UU_AMIGA_6));
    InMux I__602 (
            .O(N__3425),
            .I(N__3422));
    LocalMux I__601 (
            .O(N__3422),
            .I(N__3419));
    Odrv12 I__600 (
            .O(N__3419),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ));
    InMux I__599 (
            .O(N__3416),
            .I(N__3413));
    LocalMux I__598 (
            .O(N__3413),
            .I(N__3409));
    InMux I__597 (
            .O(N__3412),
            .I(N__3406));
    Span4Mux_v I__596 (
            .O(N__3409),
            .I(N__3403));
    LocalMux I__595 (
            .O(N__3406),
            .I(N__3399));
    Span4Mux_v I__594 (
            .O(N__3403),
            .I(N__3396));
    InMux I__593 (
            .O(N__3402),
            .I(N__3393));
    Span4Mux_h I__592 (
            .O(N__3399),
            .I(N__3390));
    Sp12to4 I__591 (
            .O(N__3396),
            .I(N__3385));
    LocalMux I__590 (
            .O(N__3393),
            .I(N__3385));
    Sp12to4 I__589 (
            .O(N__3390),
            .I(N__3382));
    Span12Mux_h I__588 (
            .O(N__3385),
            .I(N__3379));
    Odrv12 I__587 (
            .O(N__3382),
            .I(D_UU_AMIGA_in_4));
    Odrv12 I__586 (
            .O(N__3379),
            .I(D_UU_AMIGA_in_4));
    IoInMux I__585 (
            .O(N__3374),
            .I(N__3371));
    LocalMux I__584 (
            .O(N__3371),
            .I(N__3368));
    Span4Mux_s3_v I__583 (
            .O(N__3368),
            .I(N__3365));
    Span4Mux_v I__582 (
            .O(N__3365),
            .I(N__3362));
    Sp12to4 I__581 (
            .O(N__3362),
            .I(N__3359));
    Odrv12 I__580 (
            .O(N__3359),
            .I(un1_D_UU_AMIGA_4));
    InMux I__579 (
            .O(N__3356),
            .I(N__3353));
    LocalMux I__578 (
            .O(N__3353),
            .I(N__3350));
    Odrv12 I__577 (
            .O(N__3350),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ));
    InMux I__576 (
            .O(N__3347),
            .I(N__3343));
    InMux I__575 (
            .O(N__3346),
            .I(N__3340));
    LocalMux I__574 (
            .O(N__3343),
            .I(N__3337));
    LocalMux I__573 (
            .O(N__3340),
            .I(N__3333));
    Span4Mux_v I__572 (
            .O(N__3337),
            .I(N__3330));
    InMux I__571 (
            .O(N__3336),
            .I(N__3327));
    Span4Mux_v I__570 (
            .O(N__3333),
            .I(N__3324));
    Sp12to4 I__569 (
            .O(N__3330),
            .I(N__3319));
    LocalMux I__568 (
            .O(N__3327),
            .I(N__3319));
    Sp12to4 I__567 (
            .O(N__3324),
            .I(N__3316));
    Span12Mux_h I__566 (
            .O(N__3319),
            .I(N__3313));
    Span12Mux_h I__565 (
            .O(N__3316),
            .I(N__3310));
    Odrv12 I__564 (
            .O(N__3313),
            .I(D_UU_AMIGA_in_7));
    Odrv12 I__563 (
            .O(N__3310),
            .I(D_UU_AMIGA_in_7));
    IoInMux I__562 (
            .O(N__3305),
            .I(N__3302));
    LocalMux I__561 (
            .O(N__3302),
            .I(N__3299));
    IoSpan4Mux I__560 (
            .O(N__3299),
            .I(N__3296));
    Sp12to4 I__559 (
            .O(N__3296),
            .I(N__3293));
    Span12Mux_s6_v I__558 (
            .O(N__3293),
            .I(N__3290));
    Span12Mux_h I__557 (
            .O(N__3290),
            .I(N__3287));
    Odrv12 I__556 (
            .O(N__3287),
            .I(un1_D_UU_AMIGA_7));
    InMux I__555 (
            .O(N__3284),
            .I(N__3281));
    LocalMux I__554 (
            .O(N__3281),
            .I(N__3278));
    Span4Mux_v I__553 (
            .O(N__3278),
            .I(N__3275));
    Sp12to4 I__552 (
            .O(N__3275),
            .I(N__3272));
    Span12Mux_h I__551 (
            .O(N__3272),
            .I(N__3269));
    Odrv12 I__550 (
            .O(N__3269),
            .I(D_LL_AMIGA_in_4));
    IoInMux I__549 (
            .O(N__3266),
            .I(N__3263));
    LocalMux I__548 (
            .O(N__3263),
            .I(N__3260));
    IoSpan4Mux I__547 (
            .O(N__3260),
            .I(N__3257));
    IoSpan4Mux I__546 (
            .O(N__3257),
            .I(N__3254));
    Sp12to4 I__545 (
            .O(N__3254),
            .I(N__3251));
    Span12Mux_s9_h I__544 (
            .O(N__3251),
            .I(N__3248));
    Odrv12 I__543 (
            .O(N__3248),
            .I(un1_D_LL_AMIGA_4));
    InMux I__542 (
            .O(N__3245),
            .I(N__3242));
    LocalMux I__541 (
            .O(N__3242),
            .I(N__3239));
    Sp12to4 I__540 (
            .O(N__3239),
            .I(N__3236));
    Span12Mux_v I__539 (
            .O(N__3236),
            .I(N__3233));
    Odrv12 I__538 (
            .O(N__3233),
            .I(D_LM_AMIGA_in_7));
    IoInMux I__537 (
            .O(N__3230),
            .I(N__3227));
    LocalMux I__536 (
            .O(N__3227),
            .I(N__3224));
    IoSpan4Mux I__535 (
            .O(N__3224),
            .I(N__3221));
    Span4Mux_s0_h I__534 (
            .O(N__3221),
            .I(N__3218));
    Sp12to4 I__533 (
            .O(N__3218),
            .I(N__3215));
    Span12Mux_h I__532 (
            .O(N__3215),
            .I(N__3212));
    Odrv12 I__531 (
            .O(N__3212),
            .I(un1_D_LM_AMIGA_7));
    InMux I__530 (
            .O(N__3209),
            .I(N__3206));
    LocalMux I__529 (
            .O(N__3206),
            .I(N__3202));
    IoInMux I__528 (
            .O(N__3205),
            .I(N__3199));
    Span12Mux_v I__527 (
            .O(N__3202),
            .I(N__3196));
    LocalMux I__526 (
            .O(N__3199),
            .I(N__3193));
    Odrv12 I__525 (
            .O(N__3196),
            .I(A_AMIGA_c_1));
    Odrv12 I__524 (
            .O(N__3193),
            .I(A_AMIGA_c_1));
    InMux I__523 (
            .O(N__3188),
            .I(N__3185));
    LocalMux I__522 (
            .O(N__3185),
            .I(N__3182));
    Span12Mux_v I__521 (
            .O(N__3182),
            .I(N__3179));
    Span12Mux_h I__520 (
            .O(N__3179),
            .I(N__3176));
    Odrv12 I__519 (
            .O(N__3176),
            .I(D_UM_040_in_7));
    IoInMux I__518 (
            .O(N__3173),
            .I(N__3170));
    LocalMux I__517 (
            .O(N__3170),
            .I(N__3167));
    IoSpan4Mux I__516 (
            .O(N__3167),
            .I(N__3163));
    InMux I__515 (
            .O(N__3166),
            .I(N__3160));
    Span4Mux_s3_h I__514 (
            .O(N__3163),
            .I(N__3157));
    LocalMux I__513 (
            .O(N__3160),
            .I(N__3154));
    Sp12to4 I__512 (
            .O(N__3157),
            .I(N__3151));
    Span12Mux_v I__511 (
            .O(N__3154),
            .I(N__3148));
    Span12Mux_v I__510 (
            .O(N__3151),
            .I(N__3145));
    Span12Mux_v I__509 (
            .O(N__3148),
            .I(N__3142));
    Span12Mux_h I__508 (
            .O(N__3145),
            .I(N__3139));
    Span12Mux_h I__507 (
            .O(N__3142),
            .I(N__3136));
    Span12Mux_h I__506 (
            .O(N__3139),
            .I(N__3133));
    Odrv12 I__505 (
            .O(N__3136),
            .I(D_LL_040_in_7));
    Odrv12 I__504 (
            .O(N__3133),
            .I(D_LL_040_in_7));
    IoInMux I__503 (
            .O(N__3128),
            .I(N__3125));
    LocalMux I__502 (
            .O(N__3125),
            .I(N__3122));
    Span4Mux_s3_h I__501 (
            .O(N__3122),
            .I(N__3119));
    Span4Mux_h I__500 (
            .O(N__3119),
            .I(N__3116));
    Span4Mux_h I__499 (
            .O(N__3116),
            .I(N__3113));
    Odrv4 I__498 (
            .O(N__3113),
            .I(un1_D_UM_040_7));
    IoInMux I__497 (
            .O(N__3110),
            .I(N__3107));
    LocalMux I__496 (
            .O(N__3107),
            .I(N__3103));
    InMux I__495 (
            .O(N__3106),
            .I(N__3100));
    Span4Mux_s2_h I__494 (
            .O(N__3103),
            .I(N__3097));
    LocalMux I__493 (
            .O(N__3100),
            .I(N__3094));
    Span4Mux_v I__492 (
            .O(N__3097),
            .I(N__3091));
    Span4Mux_v I__491 (
            .O(N__3094),
            .I(N__3088));
    Sp12to4 I__490 (
            .O(N__3091),
            .I(N__3085));
    Span4Mux_v I__489 (
            .O(N__3088),
            .I(N__3082));
    Span12Mux_h I__488 (
            .O(N__3085),
            .I(N__3077));
    Sp12to4 I__487 (
            .O(N__3082),
            .I(N__3077));
    Span12Mux_h I__486 (
            .O(N__3077),
            .I(N__3074));
    Odrv12 I__485 (
            .O(N__3074),
            .I(D_LM_040_in_6));
    InMux I__484 (
            .O(N__3071),
            .I(N__3068));
    LocalMux I__483 (
            .O(N__3068),
            .I(N__3065));
    Span4Mux_v I__482 (
            .O(N__3065),
            .I(N__3062));
    Span4Mux_h I__481 (
            .O(N__3062),
            .I(N__3059));
    Sp12to4 I__480 (
            .O(N__3059),
            .I(N__3056));
    Span12Mux_h I__479 (
            .O(N__3056),
            .I(N__3053));
    Odrv12 I__478 (
            .O(N__3053),
            .I(D_UU_040_in_6));
    IoInMux I__477 (
            .O(N__3050),
            .I(N__3047));
    LocalMux I__476 (
            .O(N__3047),
            .I(N__3044));
    IoSpan4Mux I__475 (
            .O(N__3044),
            .I(N__3041));
    IoSpan4Mux I__474 (
            .O(N__3041),
            .I(N__3038));
    Span4Mux_s3_v I__473 (
            .O(N__3038),
            .I(N__3035));
    Odrv4 I__472 (
            .O(N__3035),
            .I(un1_D_UU_040_6));
    InMux I__471 (
            .O(N__3032),
            .I(N__3029));
    LocalMux I__470 (
            .O(N__3029),
            .I(N__3026));
    Span4Mux_v I__469 (
            .O(N__3026),
            .I(N__3023));
    Sp12to4 I__468 (
            .O(N__3023),
            .I(N__3020));
    Odrv12 I__467 (
            .O(N__3020),
            .I(D_LL_AMIGA_in_3));
    IoInMux I__466 (
            .O(N__3017),
            .I(N__3014));
    LocalMux I__465 (
            .O(N__3014),
            .I(N__3011));
    IoSpan4Mux I__464 (
            .O(N__3011),
            .I(N__3008));
    Sp12to4 I__463 (
            .O(N__3008),
            .I(N__3005));
    Span12Mux_s7_v I__462 (
            .O(N__3005),
            .I(N__3002));
    Span12Mux_h I__461 (
            .O(N__3002),
            .I(N__2999));
    Odrv12 I__460 (
            .O(N__2999),
            .I(un1_D_LL_AMIGA_3));
    IoInMux I__459 (
            .O(N__2996),
            .I(N__2993));
    LocalMux I__458 (
            .O(N__2993),
            .I(N__2990));
    IoSpan4Mux I__457 (
            .O(N__2990),
            .I(N__2987));
    Sp12to4 I__456 (
            .O(N__2987),
            .I(N__2984));
    Span12Mux_s7_h I__455 (
            .O(N__2984),
            .I(N__2981));
    Span12Mux_h I__454 (
            .O(N__2981),
            .I(N__2978));
    Odrv12 I__453 (
            .O(N__2978),
            .I(un1_D_UM_AMIGA_0));
    InMux I__452 (
            .O(N__2975),
            .I(N__2972));
    LocalMux I__451 (
            .O(N__2972),
            .I(N__2969));
    Span4Mux_v I__450 (
            .O(N__2969),
            .I(N__2965));
    InMux I__449 (
            .O(N__2968),
            .I(N__2962));
    Span4Mux_v I__448 (
            .O(N__2965),
            .I(N__2959));
    LocalMux I__447 (
            .O(N__2962),
            .I(N__2956));
    Span4Mux_v I__446 (
            .O(N__2959),
            .I(N__2952));
    Span4Mux_v I__445 (
            .O(N__2956),
            .I(N__2949));
    InMux I__444 (
            .O(N__2955),
            .I(N__2946));
    Sp12to4 I__443 (
            .O(N__2952),
            .I(N__2939));
    Sp12to4 I__442 (
            .O(N__2949),
            .I(N__2939));
    LocalMux I__441 (
            .O(N__2946),
            .I(N__2939));
    Span12Mux_h I__440 (
            .O(N__2939),
            .I(N__2936));
    Odrv12 I__439 (
            .O(N__2936),
            .I(D_UM_AMIGA_in_0));
    InMux I__438 (
            .O(N__2933),
            .I(N__2930));
    LocalMux I__437 (
            .O(N__2930),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ));
    InMux I__436 (
            .O(N__2927),
            .I(N__2924));
    LocalMux I__435 (
            .O(N__2924),
            .I(N__2921));
    Sp12to4 I__434 (
            .O(N__2921),
            .I(N__2918));
    Span12Mux_v I__433 (
            .O(N__2918),
            .I(N__2915));
    Span12Mux_h I__432 (
            .O(N__2915),
            .I(N__2912));
    Odrv12 I__431 (
            .O(N__2912),
            .I(D_UM_040_in_1));
    InMux I__430 (
            .O(N__2909),
            .I(N__2906));
    LocalMux I__429 (
            .O(N__2906),
            .I(N__2902));
    IoInMux I__428 (
            .O(N__2905),
            .I(N__2899));
    Span4Mux_v I__427 (
            .O(N__2902),
            .I(N__2896));
    LocalMux I__426 (
            .O(N__2899),
            .I(N__2893));
    Span4Mux_v I__425 (
            .O(N__2896),
            .I(N__2890));
    Span4Mux_s3_h I__424 (
            .O(N__2893),
            .I(N__2887));
    Sp12to4 I__423 (
            .O(N__2890),
            .I(N__2884));
    Sp12to4 I__422 (
            .O(N__2887),
            .I(N__2881));
    Span12Mux_h I__421 (
            .O(N__2884),
            .I(N__2878));
    Span12Mux_v I__420 (
            .O(N__2881),
            .I(N__2875));
    Span12Mux_v I__419 (
            .O(N__2878),
            .I(N__2872));
    Span12Mux_h I__418 (
            .O(N__2875),
            .I(N__2869));
    Span12Mux_h I__417 (
            .O(N__2872),
            .I(N__2866));
    Span12Mux_h I__416 (
            .O(N__2869),
            .I(N__2863));
    Odrv12 I__415 (
            .O(N__2866),
            .I(D_LL_040_in_1));
    Odrv12 I__414 (
            .O(N__2863),
            .I(D_LL_040_in_1));
    IoInMux I__413 (
            .O(N__2858),
            .I(N__2855));
    LocalMux I__412 (
            .O(N__2855),
            .I(N__2852));
    IoSpan4Mux I__411 (
            .O(N__2852),
            .I(N__2849));
    Span4Mux_s1_h I__410 (
            .O(N__2849),
            .I(N__2846));
    Span4Mux_h I__409 (
            .O(N__2846),
            .I(N__2843));
    Odrv4 I__408 (
            .O(N__2843),
            .I(un1_D_UM_040_1));
    IoInMux I__407 (
            .O(N__2840),
            .I(N__2829));
    IoInMux I__406 (
            .O(N__2839),
            .I(N__2826));
    IoInMux I__405 (
            .O(N__2838),
            .I(N__2823));
    IoInMux I__404 (
            .O(N__2837),
            .I(N__2815));
    IoInMux I__403 (
            .O(N__2836),
            .I(N__2812));
    IoInMux I__402 (
            .O(N__2835),
            .I(N__2809));
    IoInMux I__401 (
            .O(N__2834),
            .I(N__2806));
    IoInMux I__400 (
            .O(N__2833),
            .I(N__2803));
    IoInMux I__399 (
            .O(N__2832),
            .I(N__2800));
    LocalMux I__398 (
            .O(N__2829),
            .I(N__2797));
    LocalMux I__397 (
            .O(N__2826),
            .I(N__2792));
    LocalMux I__396 (
            .O(N__2823),
            .I(N__2792));
    IoInMux I__395 (
            .O(N__2822),
            .I(N__2789));
    IoInMux I__394 (
            .O(N__2821),
            .I(N__2786));
    IoInMux I__393 (
            .O(N__2820),
            .I(N__2775));
    IoInMux I__392 (
            .O(N__2819),
            .I(N__2772));
    IoInMux I__391 (
            .O(N__2818),
            .I(N__2769));
    LocalMux I__390 (
            .O(N__2815),
            .I(N__2756));
    LocalMux I__389 (
            .O(N__2812),
            .I(N__2756));
    LocalMux I__388 (
            .O(N__2809),
            .I(N__2756));
    LocalMux I__387 (
            .O(N__2806),
            .I(N__2756));
    LocalMux I__386 (
            .O(N__2803),
            .I(N__2756));
    LocalMux I__385 (
            .O(N__2800),
            .I(N__2756));
    IoSpan4Mux I__384 (
            .O(N__2797),
            .I(N__2747));
    IoSpan4Mux I__383 (
            .O(N__2792),
            .I(N__2747));
    LocalMux I__382 (
            .O(N__2789),
            .I(N__2747));
    LocalMux I__381 (
            .O(N__2786),
            .I(N__2747));
    IoInMux I__380 (
            .O(N__2785),
            .I(N__2744));
    IoInMux I__379 (
            .O(N__2784),
            .I(N__2741));
    IoInMux I__378 (
            .O(N__2783),
            .I(N__2738));
    IoInMux I__377 (
            .O(N__2782),
            .I(N__2735));
    IoInMux I__376 (
            .O(N__2781),
            .I(N__2732));
    IoInMux I__375 (
            .O(N__2780),
            .I(N__2729));
    IoInMux I__374 (
            .O(N__2779),
            .I(N__2726));
    IoInMux I__373 (
            .O(N__2778),
            .I(N__2723));
    LocalMux I__372 (
            .O(N__2775),
            .I(N__2714));
    LocalMux I__371 (
            .O(N__2772),
            .I(N__2714));
    LocalMux I__370 (
            .O(N__2769),
            .I(N__2714));
    IoSpan4Mux I__369 (
            .O(N__2756),
            .I(N__2714));
    IoSpan4Mux I__368 (
            .O(N__2747),
            .I(N__2699));
    LocalMux I__367 (
            .O(N__2744),
            .I(N__2699));
    LocalMux I__366 (
            .O(N__2741),
            .I(N__2699));
    LocalMux I__365 (
            .O(N__2738),
            .I(N__2699));
    LocalMux I__364 (
            .O(N__2735),
            .I(N__2699));
    LocalMux I__363 (
            .O(N__2732),
            .I(N__2688));
    LocalMux I__362 (
            .O(N__2729),
            .I(N__2688));
    LocalMux I__361 (
            .O(N__2726),
            .I(N__2688));
    LocalMux I__360 (
            .O(N__2723),
            .I(N__2688));
    IoSpan4Mux I__359 (
            .O(N__2714),
            .I(N__2688));
    IoInMux I__358 (
            .O(N__2713),
            .I(N__2685));
    IoInMux I__357 (
            .O(N__2712),
            .I(N__2682));
    IoInMux I__356 (
            .O(N__2711),
            .I(N__2679));
    IoInMux I__355 (
            .O(N__2710),
            .I(N__2676));
    IoSpan4Mux I__354 (
            .O(N__2699),
            .I(N__2668));
    IoSpan4Mux I__353 (
            .O(N__2688),
            .I(N__2657));
    LocalMux I__352 (
            .O(N__2685),
            .I(N__2657));
    LocalMux I__351 (
            .O(N__2682),
            .I(N__2657));
    LocalMux I__350 (
            .O(N__2679),
            .I(N__2657));
    LocalMux I__349 (
            .O(N__2676),
            .I(N__2657));
    IoInMux I__348 (
            .O(N__2675),
            .I(N__2654));
    IoInMux I__347 (
            .O(N__2674),
            .I(N__2651));
    IoInMux I__346 (
            .O(N__2673),
            .I(N__2648));
    IoInMux I__345 (
            .O(N__2672),
            .I(N__2645));
    IoInMux I__344 (
            .O(N__2671),
            .I(N__2642));
    Span4Mux_s0_h I__343 (
            .O(N__2668),
            .I(N__2639));
    IoSpan4Mux I__342 (
            .O(N__2657),
            .I(N__2628));
    LocalMux I__341 (
            .O(N__2654),
            .I(N__2628));
    LocalMux I__340 (
            .O(N__2651),
            .I(N__2628));
    LocalMux I__339 (
            .O(N__2648),
            .I(N__2628));
    LocalMux I__338 (
            .O(N__2645),
            .I(N__2628));
    LocalMux I__337 (
            .O(N__2642),
            .I(N__2625));
    Span4Mux_v I__336 (
            .O(N__2639),
            .I(N__2618));
    IoSpan4Mux I__335 (
            .O(N__2628),
            .I(N__2618));
    IoSpan4Mux I__334 (
            .O(N__2625),
            .I(N__2618));
    Span4Mux_s0_h I__333 (
            .O(N__2618),
            .I(N__2614));
    IoInMux I__332 (
            .O(N__2617),
            .I(N__2611));
    Sp12to4 I__331 (
            .O(N__2614),
            .I(N__2606));
    LocalMux I__330 (
            .O(N__2611),
            .I(N__2606));
    Odrv12 I__329 (
            .O(N__2606),
            .I(RnW_c_i_0));
    InMux I__328 (
            .O(N__2603),
            .I(N__2600));
    LocalMux I__327 (
            .O(N__2600),
            .I(N__2597));
    Span4Mux_v I__326 (
            .O(N__2597),
            .I(N__2594));
    Sp12to4 I__325 (
            .O(N__2594),
            .I(N__2591));
    Odrv12 I__324 (
            .O(N__2591),
            .I(D_LM_AMIGA_in_4));
    IoInMux I__323 (
            .O(N__2588),
            .I(N__2585));
    LocalMux I__322 (
            .O(N__2585),
            .I(N__2582));
    IoSpan4Mux I__321 (
            .O(N__2582),
            .I(N__2579));
    IoSpan4Mux I__320 (
            .O(N__2579),
            .I(N__2576));
    Span4Mux_s3_h I__319 (
            .O(N__2576),
            .I(N__2573));
    Sp12to4 I__318 (
            .O(N__2573),
            .I(N__2570));
    Span12Mux_s11_h I__317 (
            .O(N__2570),
            .I(N__2567));
    Odrv12 I__316 (
            .O(N__2567),
            .I(un1_D_LM_AMIGA_4));
    InMux I__315 (
            .O(N__2564),
            .I(N__2561));
    LocalMux I__314 (
            .O(N__2561),
            .I(N__2558));
    Span4Mux_v I__313 (
            .O(N__2558),
            .I(N__2555));
    Sp12to4 I__312 (
            .O(N__2555),
            .I(N__2552));
    Odrv12 I__311 (
            .O(N__2552),
            .I(D_LM_AMIGA_in_5));
    IoInMux I__310 (
            .O(N__2549),
            .I(N__2546));
    LocalMux I__309 (
            .O(N__2546),
            .I(N__2543));
    Span4Mux_s3_h I__308 (
            .O(N__2543),
            .I(N__2540));
    Sp12to4 I__307 (
            .O(N__2540),
            .I(N__2537));
    Span12Mux_v I__306 (
            .O(N__2537),
            .I(N__2534));
    Span12Mux_h I__305 (
            .O(N__2534),
            .I(N__2531));
    Odrv12 I__304 (
            .O(N__2531),
            .I(un1_D_LM_AMIGA_5));
    InMux I__303 (
            .O(N__2528),
            .I(N__2525));
    LocalMux I__302 (
            .O(N__2525),
            .I(N__2522));
    Span12Mux_v I__301 (
            .O(N__2522),
            .I(N__2519));
    Odrv12 I__300 (
            .O(N__2519),
            .I(D_LM_AMIGA_in_6));
    IoInMux I__299 (
            .O(N__2516),
            .I(N__2513));
    LocalMux I__298 (
            .O(N__2513),
            .I(N__2510));
    IoSpan4Mux I__297 (
            .O(N__2510),
            .I(N__2507));
    Span4Mux_s3_h I__296 (
            .O(N__2507),
            .I(N__2504));
    Span4Mux_h I__295 (
            .O(N__2504),
            .I(N__2501));
    Span4Mux_h I__294 (
            .O(N__2501),
            .I(N__2498));
    Sp12to4 I__293 (
            .O(N__2498),
            .I(N__2495));
    Odrv12 I__292 (
            .O(N__2495),
            .I(un1_D_LM_AMIGA_6));
    InMux I__291 (
            .O(N__2492),
            .I(N__2489));
    LocalMux I__290 (
            .O(N__2489),
            .I(N__2486));
    Span4Mux_v I__289 (
            .O(N__2486),
            .I(N__2483));
    Sp12to4 I__288 (
            .O(N__2483),
            .I(N__2480));
    Span12Mux_h I__287 (
            .O(N__2480),
            .I(N__2477));
    Span12Mux_h I__286 (
            .O(N__2477),
            .I(N__2474));
    Odrv12 I__285 (
            .O(N__2474),
            .I(D_UU_040_in_3));
    IoInMux I__284 (
            .O(N__2471),
            .I(N__2468));
    LocalMux I__283 (
            .O(N__2468),
            .I(N__2465));
    IoSpan4Mux I__282 (
            .O(N__2465),
            .I(N__2462));
    IoSpan4Mux I__281 (
            .O(N__2462),
            .I(N__2458));
    InMux I__280 (
            .O(N__2461),
            .I(N__2455));
    Span4Mux_s2_h I__279 (
            .O(N__2458),
            .I(N__2452));
    LocalMux I__278 (
            .O(N__2455),
            .I(N__2449));
    Sp12to4 I__277 (
            .O(N__2452),
            .I(N__2446));
    Span12Mux_s10_v I__276 (
            .O(N__2449),
            .I(N__2443));
    Span12Mux_h I__275 (
            .O(N__2446),
            .I(N__2440));
    Span12Mux_v I__274 (
            .O(N__2443),
            .I(N__2437));
    Span12Mux_h I__273 (
            .O(N__2440),
            .I(N__2434));
    Span12Mux_h I__272 (
            .O(N__2437),
            .I(N__2431));
    Odrv12 I__271 (
            .O(N__2434),
            .I(D_LM_040_in_3));
    Odrv12 I__270 (
            .O(N__2431),
            .I(D_LM_040_in_3));
    IoInMux I__269 (
            .O(N__2426),
            .I(N__2423));
    LocalMux I__268 (
            .O(N__2423),
            .I(N__2420));
    IoSpan4Mux I__267 (
            .O(N__2420),
            .I(N__2417));
    Span4Mux_s3_v I__266 (
            .O(N__2417),
            .I(N__2414));
    Span4Mux_h I__265 (
            .O(N__2414),
            .I(N__2411));
    Odrv4 I__264 (
            .O(N__2411),
            .I(un1_D_UU_040_3));
    InMux I__263 (
            .O(N__2408),
            .I(N__2405));
    LocalMux I__262 (
            .O(N__2405),
            .I(N__2402));
    Span4Mux_v I__261 (
            .O(N__2402),
            .I(N__2399));
    Sp12to4 I__260 (
            .O(N__2399),
            .I(N__2396));
    Odrv12 I__259 (
            .O(N__2396),
            .I(D_LL_AMIGA_in_0));
    IoInMux I__258 (
            .O(N__2393),
            .I(N__2390));
    LocalMux I__257 (
            .O(N__2390),
            .I(N__2387));
    Span12Mux_s9_h I__256 (
            .O(N__2387),
            .I(N__2384));
    Span12Mux_h I__255 (
            .O(N__2384),
            .I(N__2381));
    Odrv12 I__254 (
            .O(N__2381),
            .I(un1_D_LL_AMIGA_0));
    InMux I__253 (
            .O(N__2378),
            .I(N__2375));
    LocalMux I__252 (
            .O(N__2375),
            .I(N__2372));
    Span4Mux_v I__251 (
            .O(N__2372),
            .I(N__2369));
    Sp12to4 I__250 (
            .O(N__2369),
            .I(N__2366));
    Odrv12 I__249 (
            .O(N__2366),
            .I(D_LL_AMIGA_in_1));
    IoInMux I__248 (
            .O(N__2363),
            .I(N__2360));
    LocalMux I__247 (
            .O(N__2360),
            .I(N__2357));
    IoSpan4Mux I__246 (
            .O(N__2357),
            .I(N__2354));
    IoSpan4Mux I__245 (
            .O(N__2354),
            .I(N__2351));
    Span4Mux_s2_h I__244 (
            .O(N__2351),
            .I(N__2348));
    Sp12to4 I__243 (
            .O(N__2348),
            .I(N__2345));
    Span12Mux_s9_h I__242 (
            .O(N__2345),
            .I(N__2342));
    Span12Mux_h I__241 (
            .O(N__2342),
            .I(N__2339));
    Odrv12 I__240 (
            .O(N__2339),
            .I(un1_D_LL_AMIGA_1));
    InMux I__239 (
            .O(N__2336),
            .I(N__2333));
    LocalMux I__238 (
            .O(N__2333),
            .I(N__2330));
    Span12Mux_h I__237 (
            .O(N__2330),
            .I(N__2327));
    Odrv12 I__236 (
            .O(N__2327),
            .I(D_LM_AMIGA_in_3));
    IoInMux I__235 (
            .O(N__2324),
            .I(N__2321));
    LocalMux I__234 (
            .O(N__2321),
            .I(N__2318));
    IoSpan4Mux I__233 (
            .O(N__2318),
            .I(N__2315));
    IoSpan4Mux I__232 (
            .O(N__2315),
            .I(N__2312));
    Span4Mux_s0_h I__231 (
            .O(N__2312),
            .I(N__2309));
    Sp12to4 I__230 (
            .O(N__2309),
            .I(N__2306));
    Span12Mux_h I__229 (
            .O(N__2306),
            .I(N__2303));
    Odrv12 I__228 (
            .O(N__2303),
            .I(un1_D_LM_AMIGA_3));
    InMux I__227 (
            .O(N__2300),
            .I(N__2297));
    LocalMux I__226 (
            .O(N__2297),
            .I(N__2294));
    Span12Mux_h I__225 (
            .O(N__2294),
            .I(N__2291));
    Odrv12 I__224 (
            .O(N__2291),
            .I(A_040_c_1));
    InMux I__223 (
            .O(N__2288),
            .I(N__2285));
    LocalMux I__222 (
            .O(N__2285),
            .I(N__2282));
    Span4Mux_h I__221 (
            .O(N__2282),
            .I(N__2279));
    Span4Mux_v I__220 (
            .O(N__2279),
            .I(N__2276));
    Odrv4 I__219 (
            .O(N__2276),
            .I(A_040_c_0));
    IoInMux I__218 (
            .O(N__2273),
            .I(N__2270));
    LocalMux I__217 (
            .O(N__2270),
            .I(N__2267));
    Span4Mux_s2_v I__216 (
            .O(N__2267),
            .I(N__2264));
    Span4Mux_v I__215 (
            .O(N__2264),
            .I(N__2261));
    Odrv4 I__214 (
            .O(N__2261),
            .I(A_AMIGA_c_0));
    InMux I__213 (
            .O(N__2258),
            .I(N__2255));
    LocalMux I__212 (
            .O(N__2255),
            .I(N__2252));
    Span4Mux_v I__211 (
            .O(N__2252),
            .I(N__2249));
    Sp12to4 I__210 (
            .O(N__2249),
            .I(N__2246));
    Odrv12 I__209 (
            .O(N__2246),
            .I(D_LL_AMIGA_in_2));
    IoInMux I__208 (
            .O(N__2243),
            .I(N__2240));
    LocalMux I__207 (
            .O(N__2240),
            .I(N__2237));
    Span4Mux_s3_h I__206 (
            .O(N__2237),
            .I(N__2234));
    Sp12to4 I__205 (
            .O(N__2234),
            .I(N__2231));
    Span12Mux_s8_v I__204 (
            .O(N__2231),
            .I(N__2228));
    Span12Mux_h I__203 (
            .O(N__2228),
            .I(N__2225));
    Odrv12 I__202 (
            .O(N__2225),
            .I(un1_D_LL_AMIGA_2));
    InMux I__201 (
            .O(N__2222),
            .I(N__2219));
    LocalMux I__200 (
            .O(N__2219),
            .I(N__2216));
    Odrv12 I__199 (
            .O(N__2216),
            .I(D_LM_AMIGA_in_2));
    IoInMux I__198 (
            .O(N__2213),
            .I(N__2210));
    LocalMux I__197 (
            .O(N__2210),
            .I(N__2207));
    Sp12to4 I__196 (
            .O(N__2207),
            .I(N__2204));
    Span12Mux_h I__195 (
            .O(N__2204),
            .I(N__2201));
    Span12Mux_v I__194 (
            .O(N__2201),
            .I(N__2198));
    Odrv12 I__193 (
            .O(N__2198),
            .I(un1_D_LM_AMIGA_2));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .I(N__6959));
    INV \INVU111_CYCLE_SM.CYCLE_STATE_1C  (
            .O(\INVU111_CYCLE_SM.CYCLE_STATE_1C_net ),
            .I(N__6964));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net ),
            .I(N__6967));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net ),
            .I(N__6963));
    INV \INVU111_CYCLE_SM.CYCLE_STATE_0C  (
            .O(\INVU111_CYCLE_SM.CYCLE_STATE_0C_net ),
            .I(N__6966));
    INV \INVU111_CYCLE_SM.A_OUTC  (
            .O(\INVU111_CYCLE_SM.A_OUTC_net ),
            .I(N__6969));
    INV \INVU111_CYCLE_SM.TSnC  (
            .O(\INVU111_CYCLE_SM.TSnC_net ),
            .I(N__5562));
    INV \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C  (
            .O(\INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net ),
            .I(N__6965));
    INV \INVU111_CYCLE_SM.TA_EN_nessC  (
            .O(\INVU111_CYCLE_SM.TA_EN_nessC_net ),
            .I(N__6968));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net ),
            .I(N__6970));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_3  (
            .in0(N__3644),
            .in1(N__2300),
            .in2(_gnd_net_),
            .in3(N__5512),
            .lcout(A_AMIGA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_7  (
            .in0(N__2288),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5513),
            .lcout(A_AMIGA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_5_3_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_5_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_5_3_0  (
            .in0(N__4797),
            .in1(N__2258),
            .in2(_gnd_net_),
            .in3(N__6327),
            .lcout(un1_D_LL_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_5_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_5_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_5_12_5  (
            .in0(N__6316),
            .in1(N__5701),
            .in2(_gnd_net_),
            .in3(N__2222),
            .lcout(un1_D_LM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_5_15_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_5_15_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_5_15_5  (
            .in0(N__6328),
            .in1(N__2927),
            .in2(_gnd_net_),
            .in3(N__2909),
            .lcout(un1_D_UM_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RnW_c_sbtinv_LC_6_11_6.C_ON=1'b0;
    defparam RnW_c_sbtinv_LC_6_11_6.SEQ_MODE=4'b0000;
    defparam RnW_c_sbtinv_LC_6_11_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 RnW_c_sbtinv_LC_6_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4001),
            .lcout(RnW_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_6_13_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_6_13_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_6_13_5  (
            .in0(N__2603),
            .in1(N__6297),
            .in2(_gnd_net_),
            .in3(N__3412),
            .lcout(un1_D_LM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_6_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_6_14_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_6_14_1  (
            .in0(N__2564),
            .in1(N__6299),
            .in2(_gnd_net_),
            .in3(N__5755),
            .lcout(un1_D_LM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_6_17_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_6_17_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_6_17_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_6_17_4  (
            .in0(N__3477),
            .in1(N__6329),
            .in2(_gnd_net_),
            .in3(N__2528),
            .lcout(un1_D_LM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_6_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_6_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_6_20_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_6_20_2  (
            .in0(N__2492),
            .in1(N__6361),
            .in2(_gnd_net_),
            .in3(N__2461),
            .lcout(un1_D_UU_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_7_1_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_7_1_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_7_1_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_7_1_6  (
            .in0(N__2408),
            .in1(N__6326),
            .in2(_gnd_net_),
            .in3(N__2975),
            .lcout(un1_D_LL_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_7_3_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_7_3_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_7_3_2  (
            .in0(N__2378),
            .in1(N__6289),
            .in2(_gnd_net_),
            .in3(N__4568),
            .lcout(un1_D_LL_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_7_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_7_11_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_7_11_0  (
            .in0(N__2336),
            .in1(N__6249),
            .in2(_gnd_net_),
            .in3(N__5933),
            .lcout(un1_D_LM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_7_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_7_15_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_7_15_0  (
            .in0(N__3245),
            .in1(N__6298),
            .in2(_gnd_net_),
            .in3(N__3336),
            .lcout(un1_D_LM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIM3VM1_LC_8_7_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIM3VM1_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIM3VM1_LC_8_7_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIM3VM1_LC_8_7_6  (
            .in0(N__3209),
            .in1(N__6410),
            .in2(_gnd_net_),
            .in3(N__5500),
            .lcout(\U111_CYCLE_SM.FLIP ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_8_12_4.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_8_12_4.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_8_12_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_8_12_4 (
            .in0(N__4702),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_8_19_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_8_19_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_8_19_4  (
            .in0(N__3188),
            .in1(N__6279),
            .in2(_gnd_net_),
            .in3(N__3166),
            .lcout(un1_D_UM_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_8_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_8_20_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_8_20_2  (
            .in0(N__3106),
            .in1(N__6280),
            .in2(_gnd_net_),
            .in3(N__3071),
            .lcout(un1_D_UU_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_9_2_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_9_2_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_9_2_2  (
            .in0(N__3032),
            .in1(N__6269),
            .in2(_gnd_net_),
            .in3(N__5144),
            .lcout(un1_D_LL_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_9_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_9_11_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_9_11_1  (
            .in0(N__2933),
            .in1(N__2968),
            .in2(_gnd_net_),
            .in3(N__5416),
            .lcout(un1_D_UM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_9_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_9_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2955),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net ),
            .ce(N__5231),
            .sr(N__5193));
    defparam \U111_CYCLE_SM.TA_EN_ness_LC_9_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_EN_ness_LC_9_13_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.TA_EN_ness_LC_9_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.TA_EN_ness_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5285),
            .lcout(\U111_CYCLE_SM.TA_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TA_EN_nessC_net ),
            .ce(N__3593),
            .sr(N__3607));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_9_14_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_9_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3416),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net ),
            .ce(N__5232),
            .sr(N__5189));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_9_14_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_9_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3347),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net ),
            .ce(N__5232),
            .sr(N__5189));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_9_14_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_9_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3491),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net ),
            .ce(N__5232),
            .sr(N__5189));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_9_18_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_9_18_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_9_18_5  (
            .in0(N__3581),
            .in1(N__6317),
            .in2(_gnd_net_),
            .in3(N__3530),
            .lcout(un1_D_UU_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_9_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_9_19_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_9_19_2  (
            .in0(N__3490),
            .in1(N__3458),
            .in2(_gnd_net_),
            .in3(N__5485),
            .lcout(un1_D_UU_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_9_19_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_9_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_9_19_5  (
            .in0(N__5484),
            .in1(N__3425),
            .in2(_gnd_net_),
            .in3(N__3402),
            .lcout(un1_D_UU_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_9_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_9_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_9_20_1  (
            .in0(N__5502),
            .in1(N__3356),
            .in2(_gnd_net_),
            .in3(N__3346),
            .lcout(un1_D_UU_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_10_3_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_10_3_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_10_3_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_10_3_7  (
            .in0(N__4423),
            .in1(N__6290),
            .in2(_gnd_net_),
            .in3(N__3284),
            .lcout(un1_D_LL_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_10_7_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_10_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_10_7_5  (
            .in0(N__4190),
            .in1(N__6170),
            .in2(_gnd_net_),
            .in3(N__3719),
            .lcout(un1_D_LM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_10_10_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_10_10_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_10_10_6  (
            .in0(N__6247),
            .in1(N__4499),
            .in2(_gnd_net_),
            .in3(N__3680),
            .lcout(un1_D_LM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TSn_LC_10_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TSn_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TSn_LC_10_11_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U111_CYCLE_SM.TSn_LC_10_11_0  (
            .in0(_gnd_net_),
            .in1(N__4738),
            .in2(_gnd_net_),
            .in3(N__4075),
            .lcout(TSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TSnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A_OUT_LC_10_12_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A_OUT_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.A_OUT_LC_10_12_0 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \U111_CYCLE_SM.A_OUT_LC_10_12_0  (
            .in0(N__3631),
            .in1(N__3617),
            .in2(N__4752),
            .in3(N__5279),
            .lcout(\U111_CYCLE_SM.A_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.A_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_10_12_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_10_12_1 .LUT_INIT=16'b0010010100100000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_10_12_1  (
            .in0(N__5277),
            .in1(N__4668),
            .in2(N__4616),
            .in3(N__4039),
            .lcout(),
            .ltout(\U111_CYCLE_SM.LW_CYCLE_r_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_LC_10_12_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_CYCLE_LC_10_12_2 .LUT_INIT=16'b0000100011001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_LC_10_12_2  (
            .in0(N__5409),
            .in1(N__4742),
            .in2(N__3620),
            .in3(N__5278),
            .lcout(\U111_CYCLE_SM.LW_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.A_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_10_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_10_12_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_0_LC_10_12_3  (
            .in0(N__5276),
            .in1(_gnd_net_),
            .in2(N__4615),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.TS_EN10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_START_RNIIU7U_LC_10_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_RNIIU7U_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_RNIIU7U_LC_10_12_4 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_START_RNIIU7U_LC_10_12_4  (
            .in0(N__5408),
            .in1(N__4605),
            .in2(N__4040),
            .in3(N__5275),
            .lcout(\U111_CYCLE_SM.un1_CYCLE_STATE_1_0 ),
            .ltout(\U111_CYCLE_SM.un1_CYCLE_STATE_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_EN_ness_RNO_LC_10_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_EN_ness_RNO_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_EN_ness_RNO_LC_10_12_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U111_CYCLE_SM.TA_EN_ness_RNO_LC_10_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3611),
            .in3(N__3608),
            .lcout(\U111_CYCLE_SM.un1_CYCLE_STATE_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_LC_10_12_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TS_EN_LC_10_12_6 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \U111_CYCLE_SM.TS_EN_LC_10_12_6  (
            .in0(N__5240),
            .in1(N__4085),
            .in2(N__4079),
            .in3(N__4746),
            .lcout(\U111_CYCLE_SM.TS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.A_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_START_LC_10_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_LC_10_12_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_START_LC_10_12_7  (
            .in0(N__6403),
            .in1(N__4051),
            .in2(N__4753),
            .in3(N__6442),
            .lcout(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.A_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_10_13_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_10_13_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_10_13_4 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_0_LC_10_13_4  (
            .in0(N__5274),
            .in1(N__4669),
            .in2(N__4614),
            .in3(N__4747),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.CYCLE_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_10_13_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_10_13_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_10_13_5  (
            .in0(N__4670),
            .in1(N__5273),
            .in2(_gnd_net_),
            .in3(N__4601),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa ),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_10_13_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_10_13_6 .LUT_INIT=16'b0101000011111111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_10_13_6  (
            .in0(N__3943),
            .in1(_gnd_net_),
            .in2(N__3731),
            .in3(N__4748),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0 ),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_10_13_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_10_13_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3728),
            .in3(N__3725),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_10_14_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_10_14_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_10_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4424),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net ),
            .ce(N__5230),
            .sr(N__5188));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_10_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_10_14_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_10_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4564),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net ),
            .ce(N__5230),
            .sr(N__5188));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_10_14_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_10_14_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_10_14_2  (
            .in0(N__4495),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net ),
            .ce(N__5230),
            .sr(N__5188));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_10_14_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_10_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_10_14_4  (
            .in0(N__4183),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net ),
            .ce(N__5230),
            .sr(N__5188));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_10_15_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_10_15_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_10_15_4  (
            .in0(N__4574),
            .in1(N__5444),
            .in2(_gnd_net_),
            .in3(N__4557),
            .lcout(un1_D_UM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_10_17_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_10_17_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_10_17_7  (
            .in0(N__4488),
            .in1(N__4463),
            .in2(_gnd_net_),
            .in3(N__5476),
            .lcout(un1_D_UU_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_10_18_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_10_18_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_10_18_1  (
            .in0(N__5477),
            .in1(N__4433),
            .in2(_gnd_net_),
            .in3(N__4419),
            .lcout(un1_D_UM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_10_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_10_20_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_10_20_1  (
            .in0(N__6366),
            .in1(N__4352),
            .in2(_gnd_net_),
            .in3(N__4327),
            .lcout(un1_D_UU_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_10_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_10_20_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_10_20_2  (
            .in0(N__4274),
            .in1(N__6365),
            .in2(_gnd_net_),
            .in3(N__4255),
            .lcout(un1_D_UU_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_10_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_10_20_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_10_20_4  (
            .in0(N__4202),
            .in1(N__4171),
            .in2(_gnd_net_),
            .in3(N__5501),
            .lcout(un1_D_UU_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_11_6_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_11_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_11_6_0  (
            .in0(N__6234),
            .in1(N__5360),
            .in2(_gnd_net_),
            .in3(N__4127),
            .lcout(un1_D_LL_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_3  (
            .in0(N__5642),
            .in1(N__6233),
            .in2(_gnd_net_),
            .in3(N__4973),
            .lcout(un1_D_LL_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_11_7_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_11_7_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_11_7_0  (
            .in0(N__5048),
            .in1(N__6232),
            .in2(_gnd_net_),
            .in3(N__4934),
            .lcout(un1_D_LL_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_11_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_11_10_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_11_10_0  (
            .in0(N__6248),
            .in1(N__4892),
            .in2(_gnd_net_),
            .in3(N__4873),
            .lcout(un1_D_UM_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_11_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_11_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_11_11_3  (
            .in0(N__4799),
            .in1(N__4760),
            .in2(_gnd_net_),
            .in3(N__5417),
            .lcout(un1_D_UM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_11_12_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_11_12_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_11_12_0  (
            .in0(N__5346),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net ),
            .ce(N__5233),
            .sr(N__5194));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_11_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_11_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4798),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net ),
            .ce(N__5233),
            .sr(N__5194));
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_13_0 .LUT_INIT=16'b1001000010100000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_13_0  (
            .in0(N__5281),
            .in1(N__4666),
            .in2(N__4754),
            .in3(N__4613),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.CYCLE_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_EN_ness_RNIPNOD_LC_11_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_EN_ness_RNIPNOD_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_EN_ness_RNIPNOD_LC_11_13_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U111_CYCLE_SM.TA_EN_ness_RNIPNOD_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__4679),
            .in2(_gnd_net_),
            .in3(N__4667),
            .lcout(TAn_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_11_13_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_11_13_5 .LUT_INIT=16'b0011001100000010;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_1_LC_11_13_5  (
            .in0(N__5569),
            .in1(N__4612),
            .in2(N__5303),
            .in3(N__5280),
            .lcout(\U111_CYCLE_SM.TS_EN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_11_14_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_11_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5140),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__5234),
            .sr(N__5195));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5705),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__5234),
            .sr(N__5195));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_11_14_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_11_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5047),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__5234),
            .sr(N__5195));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_11_14_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_11_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_11_14_3  (
            .in0(N__5635),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__5234),
            .sr(N__5195));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_11_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_11_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_11_14_5  (
            .in0(N__5774),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__5234),
            .sr(N__5195));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_11_14_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_11_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_11_14_6  (
            .in0(N__5926),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__5234),
            .sr(N__5195));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_11_17_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_11_17_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_11_17_5  (
            .in0(N__5139),
            .in1(N__5087),
            .in2(_gnd_net_),
            .in3(N__5486),
            .lcout(un1_D_UM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_11_18_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_11_18_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_11_18_2  (
            .in0(N__5487),
            .in1(N__5057),
            .in2(_gnd_net_),
            .in3(N__5040),
            .lcout(un1_D_UM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_11_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_11_19_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_11_19_2  (
            .in0(N__6035),
            .in1(N__6368),
            .in2(_gnd_net_),
            .in3(N__5984),
            .lcout(un1_D_UM_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_11_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_11_20_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_11_20_2  (
            .in0(N__5505),
            .in1(N__5942),
            .in2(_gnd_net_),
            .in3(N__5925),
            .lcout(un1_D_UU_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_11_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_11_20_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_11_20_4  (
            .in0(N__6367),
            .in1(N__5870),
            .in2(_gnd_net_),
            .in3(N__5845),
            .lcout(un1_D_UM_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_11_20_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_11_20_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_11_20_5  (
            .in0(N__5786),
            .in1(N__5767),
            .in2(_gnd_net_),
            .in3(N__5506),
            .lcout(un1_D_UU_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_20_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_20_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_20_6  (
            .in0(N__5504),
            .in1(N__5714),
            .in2(_gnd_net_),
            .in3(N__5697),
            .lcout(un1_D_UU_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_11_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_11_20_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_11_20_7  (
            .in0(N__5623),
            .in1(N__5600),
            .in2(_gnd_net_),
            .in3(N__5503),
            .lcout(un1_D_UM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_2.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5570),
            .lcout(GB_BUFFER_CLK40_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_12_12_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_12_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_12_12_1  (
            .in0(N__5440),
            .in1(N__5366),
            .in2(_gnd_net_),
            .in3(N__5353),
            .lcout(un1_D_UM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_12_5.C_ON=1'b0;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_12_5.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6974),
            .lcout(GB_BUFFER_CLK80_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_12_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_12_20_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_12_20_4  (
            .in0(N__6871),
            .in1(N__6362),
            .in2(_gnd_net_),
            .in3(N__6830),
            .lcout(un1_D_UU_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_12_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_12_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_12_20_7  (
            .in0(N__6363),
            .in1(N__6787),
            .in2(_gnd_net_),
            .in3(N__6752),
            .lcout(un1_D_UU_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_13_9_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_13_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_13_9_3  (
            .in0(N__6314),
            .in1(N__6719),
            .in2(_gnd_net_),
            .in3(N__6703),
            .lcout(un1_D_UM_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_13_12_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_13_12_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_13_12_6  (
            .in0(N__6640),
            .in1(N__6315),
            .in2(_gnd_net_),
            .in3(N__6599),
            .lcout(un1_D_UM_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_13_18_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_13_18_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_13_18_4  (
            .in0(N__6566),
            .in1(N__6341),
            .in2(_gnd_net_),
            .in3(N__6521),
            .lcout(un1_D_UM_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_TRANS_LC_13_18_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_13_18_7 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \U111_CYCLE_SM.LW_TRANS_LC_13_18_7  (
            .in0(N__6482),
            .in1(N__6464),
            .in2(_gnd_net_),
            .in3(N__6446),
            .lcout(\U111_CYCLE_SM.LW_TRANS_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_13_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_13_20_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_13_20_7  (
            .in0(N__6386),
            .in1(N__6364),
            .in2(_gnd_net_),
            .in3(N__6085),
            .lcout(un1_D_UU_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_19_17_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_19_17_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_19_17_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_19_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U111_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     May 8 2025 19:59:06

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    DBRn : in std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__12817\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.N_458_cascade_\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a2_0_cascade_\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_442_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_5_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_1_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_1_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_1_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_2_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_433\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_4_i_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_65\ : std_logic;
signal \U712_CHIP_RAM.N_173_cascade_\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_2_3\ : std_logic;
signal \U712_CHIP_RAM.N_301_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_0_1_cascade_\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.LATCH_CLK_6\ : std_logic;
signal \U712_CHIP_RAM.N_396_cascade_\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \U712_CHIP_RAM.N_315\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_336\ : std_logic;
signal \U712_CHIP_RAM.N_372\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_9\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_191_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_191_0\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_0_4\ : std_logic;
signal \U712_CHIP_RAM.N_191\ : std_logic;
signal \U712_CHIP_RAM.N_327\ : std_logic;
signal \U712_CHIP_RAM.N_300\ : std_logic;
signal \U712_CHIP_RAM.N_370\ : std_logic;
signal \U712_CHIP_RAM.N_301\ : std_logic;
signal \U712_CHIP_RAM.N_466_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_299_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.N_399_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_0_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_310\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_385\ : std_logic;
signal \U712_CHIP_RAM.N_182\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_382\ : std_logic;
signal \U712_CHIP_RAM.N_534\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_cascade_\ : std_logic;
signal \U712_REG_SM.N_411_cascade_\ : std_logic;
signal \U712_BYTE_ENABLE.N_446_cascade_\ : std_logic;
signal \N_52_i\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_1\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_2\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_3\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_4\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_5\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_6\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.N_353\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DBENn_7_0_0\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_471\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_429\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_319\ : std_logic;
signal \U712_CHIP_RAM.N_359\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_419_cascade_\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_299\ : std_logic;
signal \U712_CHIP_RAM.N_307\ : std_logic;
signal \U712_CHIP_RAM.N_434\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto7_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_REG_SM.N_322_cascade_\ : std_logic;
signal \U712_REG_SM.N_367_cascade_\ : std_logic;
signal \U712_REG_SM.N_408_cascade_\ : std_logic;
signal \U712_REG_SM.N_367\ : std_logic;
signal \U712_REG_SM.N_410\ : std_logic;
signal \U712_REG_SM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_REG_SM.REGENn_e_1\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \U712_REG_SM.N_322\ : std_logic;
signal \U712_REG_SM.N_131\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLE_5_i_a2_4_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_456\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLE_5_i_a2_5\ : std_logic;
signal \DMA_LATCH_EN_c\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_466\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_REG_SM.N_401_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_324_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_2\ : std_logic;
signal \U712_REG_SM.STATE_COUNTc_0_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_424\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0\ : std_logic;
signal \N_170_i\ : std_logic;
signal \U712_REG_SM.N_325_cascade_\ : std_logic;
signal \U712_REG_SM.N_302\ : std_logic;
signal \U712_REG_SM.N_302_cascade_\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \N_160_i\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_404\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_309_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_309\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1_cascade_\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i_0\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_3\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.START_RSTZ0\ : std_logic;
signal \U712_BYTE_ENABLE.N_443_cascade_\ : std_logic;
signal \N_54_i\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_1\ : std_logic;
signal \U712_CYCLE_TERM.N_452_cascade_\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_BYTE_ENABLE.N_421_cascade_\ : std_logic;
signal \N_168_i\ : std_logic;
signal \U712_CYCLE_TERM.N_326\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \U712_BYTE_ENABLE.N_425\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_402\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.un1_REGENn_0_sqmuxa_0\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \N_166\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \U712_BYTE_ENABLE.N_298_i\ : std_logic;
signal \U712_REG_SM.N_459\ : std_logic;
signal \N_390_i\ : std_logic;
signal \N_389_i\ : std_logic;
signal \A_c_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \N_189\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_2\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \DMA_WRITE_CYCLE\ : std_logic;
signal \RnW_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \DRDDIR_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    TBIn <= \TBIn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    TCIn <= \TCIn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4347\,
            RESETB => \N__5871\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12817\,
            DIN => \N__12816\,
            DOUT => \N__12815\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12817\,
            PADOUT => \N__12816\,
            PADIN => \N__12815\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8787\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12808\,
            DIN => \N__12807\,
            DOUT => \N__12806\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12808\,
            PADOUT => \N__12807\,
            PADIN => \N__12806\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12799\,
            DIN => \N__12798\,
            DOUT => \N__12797\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12799\,
            PADOUT => \N__12798\,
            PADIN => \N__12797\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9288\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12790\,
            DIN => \N__12789\,
            DOUT => \N__12788\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12790\,
            PADOUT => \N__12789\,
            PADIN => \N__12788\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11808\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12781\,
            DIN => \N__12780\,
            DOUT => \N__12779\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12781\,
            PADOUT => \N__12780\,
            PADIN => \N__12779\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12772\,
            DIN => \N__12771\,
            DOUT => \N__12770\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12772\,
            PADOUT => \N__12771\,
            PADIN => \N__12770\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12763\,
            DIN => \N__12762\,
            DOUT => \N__12761\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12763\,
            PADOUT => \N__12762\,
            PADIN => \N__12761\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12754\,
            DIN => \N__12753\,
            DOUT => \N__12752\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12754\,
            PADOUT => \N__12753\,
            PADIN => \N__12752\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12745\,
            DIN => \N__12744\,
            DOUT => \N__12743\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12745\,
            PADOUT => \N__12744\,
            PADIN => \N__12743\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12736\,
            DIN => \N__12735\,
            DOUT => \N__12734\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12736\,
            PADOUT => \N__12735\,
            PADIN => \N__12734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12727\,
            DIN => \N__12726\,
            DOUT => \N__12725\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12727\,
            PADOUT => \N__12726\,
            PADIN => \N__12725\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12718\,
            DIN => \N__12717\,
            DOUT => \N__12716\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12718\,
            PADOUT => \N__12717\,
            PADIN => \N__12716\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6840\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12709\,
            DIN => \N__12708\,
            DOUT => \N__12707\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12709\,
            PADOUT => \N__12708\,
            PADIN => \N__12707\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9903\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12700\,
            DIN => \N__12699\,
            DOUT => \N__12698\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12700\,
            PADOUT => \N__12699\,
            PADIN => \N__12698\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12691\,
            DIN => \N__12690\,
            DOUT => \N__12689\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12691\,
            PADOUT => \N__12690\,
            PADIN => \N__12689\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12682\,
            DIN => \N__12681\,
            DOUT => \N__12680\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12682\,
            PADOUT => \N__12681\,
            PADIN => \N__12680\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12673\,
            DIN => \N__12672\,
            DOUT => \N__12671\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12673\,
            PADOUT => \N__12672\,
            PADIN => \N__12671\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4584\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12664\,
            DIN => \N__12663\,
            DOUT => \N__12662\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12664\,
            PADOUT => \N__12663\,
            PADIN => \N__12662\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12655\,
            DIN => \N__12654\,
            DOUT => \N__12653\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12655\,
            PADOUT => \N__12654\,
            PADIN => \N__12653\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12646\,
            DIN => \N__12645\,
            DOUT => \N__12644\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12646\,
            PADOUT => \N__12645\,
            PADIN => \N__12644\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6678\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12637\,
            DIN => \N__12636\,
            DOUT => \N__12635\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12637\,
            PADOUT => \N__12636\,
            PADIN => \N__12635\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12628\,
            DIN => \N__12627\,
            DOUT => \N__12626\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12628\,
            PADOUT => \N__12627\,
            PADIN => \N__12626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10050\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12619\,
            DIN => \N__12618\,
            DOUT => \N__12617\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12619\,
            PADOUT => \N__12618\,
            PADIN => \N__12617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12610\,
            DIN => \N__12609\,
            DOUT => \N__12608\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12610\,
            PADOUT => \N__12609\,
            PADIN => \N__12608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10326\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12601\,
            DIN => \N__12600\,
            DOUT => \N__12599\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12601\,
            PADOUT => \N__12600\,
            PADIN => \N__12599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8561\,
            DIN0 => OPEN,
            DOUT0 => \N__7869\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12592\,
            DIN => \N__12591\,
            DOUT => \N__12590\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12592\,
            PADOUT => \N__12591\,
            PADIN => \N__12590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12583\,
            DIN => \N__12582\,
            DOUT => \N__12581\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12583\,
            PADOUT => \N__12582\,
            PADIN => \N__12581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12574\,
            DIN => \N__12573\,
            DOUT => \N__12572\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12574\,
            PADOUT => \N__12573\,
            PADIN => \N__12572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12565\,
            DIN => \N__12564\,
            DOUT => \N__12563\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12565\,
            PADOUT => \N__12564\,
            PADIN => \N__12563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12556\,
            DIN => \N__12555\,
            DOUT => \N__12554\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12556\,
            PADOUT => \N__12555\,
            PADIN => \N__12554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12547\,
            DIN => \N__12546\,
            DOUT => \N__12545\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12547\,
            PADOUT => \N__12546\,
            PADIN => \N__12545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6759\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12538\,
            DIN => \N__12537\,
            DOUT => \N__12536\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12538\,
            PADOUT => \N__12537\,
            PADIN => \N__12536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12529\,
            DIN => \N__12528\,
            DOUT => \N__12527\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12529\,
            PADOUT => \N__12528\,
            PADIN => \N__12527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12520\,
            DIN => \N__12519\,
            DOUT => \N__12518\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12520\,
            PADOUT => \N__12519\,
            PADIN => \N__12518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12511\,
            DIN => \N__12510\,
            DOUT => \N__12509\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12511\,
            PADOUT => \N__12510\,
            PADIN => \N__12509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12502\,
            DIN => \N__12501\,
            DOUT => \N__12500\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12502\,
            PADOUT => \N__12501\,
            PADIN => \N__12500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12493\,
            DIN => \N__12492\,
            DOUT => \N__12491\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12493\,
            PADOUT => \N__12492\,
            PADIN => \N__12491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8055\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12484\,
            DIN => \N__12483\,
            DOUT => \N__12482\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12484\,
            PADOUT => \N__12483\,
            PADIN => \N__12482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12475\,
            DIN => \N__12474\,
            DOUT => \N__12473\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12475\,
            PADOUT => \N__12474\,
            PADIN => \N__12473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12466\,
            DIN => \N__12465\,
            DOUT => \N__12464\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12466\,
            PADOUT => \N__12465\,
            PADIN => \N__12464\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8091\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12457\,
            DIN => \N__12456\,
            DOUT => \N__12455\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12457\,
            PADOUT => \N__12456\,
            PADIN => \N__12455\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6720\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12448\,
            DIN => \N__12447\,
            DOUT => \N__12446\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12448\,
            PADOUT => \N__12447\,
            PADIN => \N__12446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12439\,
            DIN => \N__12438\,
            DOUT => \N__12437\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12439\,
            PADOUT => \N__12438\,
            PADIN => \N__12437\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6741\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12430\,
            DIN => \N__12429\,
            DOUT => \N__12428\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12430\,
            PADOUT => \N__12429\,
            PADIN => \N__12428\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6963\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12421\,
            DIN => \N__12420\,
            DOUT => \N__12419\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12421\,
            PADOUT => \N__12420\,
            PADIN => \N__12419\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6627\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12412\,
            DIN => \N__12411\,
            DOUT => \N__12410\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12412\,
            PADOUT => \N__12411\,
            PADIN => \N__12410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12403\,
            DIN => \N__12402\,
            DOUT => \N__12401\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12403\,
            PADOUT => \N__12402\,
            PADIN => \N__12401\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8415\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12394\,
            DIN => \N__12393\,
            DOUT => \N__12392\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12394\,
            PADOUT => \N__12393\,
            PADIN => \N__12392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8562\,
            DIN0 => OPEN,
            DOUT0 => \N__7868\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12385\,
            DIN => \N__12384\,
            DOUT => \N__12383\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12385\,
            PADOUT => \N__12384\,
            PADIN => \N__12383\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9996\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12376\,
            DIN => \N__12375\,
            DOUT => \N__12374\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12376\,
            PADOUT => \N__12375\,
            PADIN => \N__12374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6054\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12367\,
            DIN => \N__12366\,
            DOUT => \N__12365\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12367\,
            PADOUT => \N__12366\,
            PADIN => \N__12365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7134\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12358\,
            DIN => \N__12357\,
            DOUT => \N__12356\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12358\,
            PADOUT => \N__12357\,
            PADIN => \N__12356\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12349\,
            DIN => \N__12348\,
            DOUT => \N__12347\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12349\,
            PADOUT => \N__12348\,
            PADIN => \N__12347\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12340\,
            DIN => \N__12339\,
            DOUT => \N__12338\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12340\,
            PADOUT => \N__12339\,
            PADIN => \N__12338\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5814\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12331\,
            DIN => \N__12330\,
            DOUT => \N__12329\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12331\,
            PADOUT => \N__12330\,
            PADIN => \N__12329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12322\,
            DIN => \N__12321\,
            DOUT => \N__12320\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12322\,
            PADOUT => \N__12321\,
            PADIN => \N__12320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12313\,
            DIN => \N__12312\,
            DOUT => \N__12311\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12313\,
            PADOUT => \N__12312\,
            PADIN => \N__12311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8313\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12304\,
            DIN => \N__12303\,
            DOUT => \N__12302\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12304\,
            PADOUT => \N__12303\,
            PADIN => \N__12302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9888\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12295\,
            DIN => \N__12294\,
            DOUT => \N__12293\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12295\,
            PADOUT => \N__12294\,
            PADIN => \N__12293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12286\,
            DIN => \N__12285\,
            DOUT => \N__12284\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12286\,
            PADOUT => \N__12285\,
            PADIN => \N__12284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8880\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12277\,
            DIN => \N__12276\,
            DOUT => \N__12275\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12277\,
            PADOUT => \N__12276\,
            PADIN => \N__12275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8560\,
            DIN0 => OPEN,
            DOUT0 => \N__7861\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12268\,
            DIN => \N__12267\,
            DOUT => \N__12266\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12268\,
            PADOUT => \N__12267\,
            PADIN => \N__12266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7104\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12259\,
            DIN => \N__12258\,
            DOUT => \N__12257\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12259\,
            PADOUT => \N__12258\,
            PADIN => \N__12257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12250\,
            DIN => \N__12249\,
            DOUT => \N__12248\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12250\,
            PADOUT => \N__12249\,
            PADIN => \N__12248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12241\,
            DIN => \N__12240\,
            DOUT => \N__12239\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12241\,
            PADOUT => \N__12240\,
            PADIN => \N__12239\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4764\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12232\,
            DIN => \N__12231\,
            DOUT => \N__12230\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12232\,
            PADOUT => \N__12231\,
            PADIN => \N__12230\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12223\,
            DIN => \N__12222\,
            DOUT => \N__12221\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12223\,
            PADOUT => \N__12222\,
            PADIN => \N__12221\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12214\,
            DIN => \N__12213\,
            DOUT => \N__12212\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12214\,
            PADOUT => \N__12213\,
            PADIN => \N__12212\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8205\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12205\,
            DIN => \N__12204\,
            DOUT => \N__12203\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12205\,
            PADOUT => \N__12204\,
            PADIN => \N__12203\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12196\,
            DIN => \N__12195\,
            DOUT => \N__12194\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12196\,
            PADOUT => \N__12195\,
            PADIN => \N__12194\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12187\,
            DIN => \N__12186\,
            DOUT => \N__12185\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12187\,
            PADOUT => \N__12186\,
            PADIN => \N__12185\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5838\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12178\,
            DIN => \N__12177\,
            DOUT => \N__12176\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12178\,
            PADOUT => \N__12177\,
            PADIN => \N__12176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9510\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12169\,
            DIN => \N__12168\,
            DOUT => \N__12167\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12169\,
            PADOUT => \N__12168\,
            PADIN => \N__12167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9468\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12160\,
            DIN => \N__12159\,
            DOUT => \N__12158\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12160\,
            PADOUT => \N__12159\,
            PADIN => \N__12158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4395\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12151\,
            DIN => \N__12150\,
            DOUT => \N__12149\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12151\,
            PADOUT => \N__12150\,
            PADIN => \N__12149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12142\,
            DIN => \N__12141\,
            DOUT => \N__12140\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12142\,
            PADOUT => \N__12141\,
            PADIN => \N__12140\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12133\,
            DIN => \N__12132\,
            DOUT => \N__12131\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12133\,
            PADOUT => \N__12132\,
            PADIN => \N__12131\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6915\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12124\,
            DIN => \N__12123\,
            DOUT => \N__12122\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12124\,
            PADOUT => \N__12123\,
            PADIN => \N__12122\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12115\,
            DIN => \N__12114\,
            DOUT => \N__12113\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12115\,
            PADOUT => \N__12114\,
            PADIN => \N__12113\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12106\,
            DIN => \N__12105\,
            DOUT => \N__12104\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12106\,
            PADOUT => \N__12105\,
            PADIN => \N__12104\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4656\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12097\,
            DIN => \N__12096\,
            DOUT => \N__12095\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12097\,
            PADOUT => \N__12096\,
            PADIN => \N__12095\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9645\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12088\,
            DIN => \N__12087\,
            DOUT => \N__12086\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12088\,
            PADOUT => \N__12087\,
            PADIN => \N__12086\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8616\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12079\,
            DIN => \N__12078\,
            DOUT => \N__12077\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12079\,
            PADOUT => \N__12078\,
            PADIN => \N__12077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12070\,
            DIN => \N__12069\,
            DOUT => \N__12068\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12070\,
            PADOUT => \N__12069\,
            PADIN => \N__12068\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8615\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12061\,
            DIN => \N__12060\,
            DOUT => \N__12059\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12061\,
            PADOUT => \N__12060\,
            PADIN => \N__12059\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4362\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12052\,
            DIN => \N__12051\,
            DOUT => \N__12050\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12052\,
            PADOUT => \N__12051\,
            PADIN => \N__12050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6939\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12043\,
            DIN => \N__12042\,
            DOUT => \N__12041\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12043\,
            PADOUT => \N__12042\,
            PADIN => \N__12041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12034\,
            DIN => \N__12033\,
            DOUT => \N__12032\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12034\,
            PADOUT => \N__12033\,
            PADIN => \N__12032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12025\,
            DIN => \N__12024\,
            DOUT => \N__12023\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12025\,
            PADOUT => \N__12024\,
            PADIN => \N__12023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12016\,
            DIN => \N__12015\,
            DOUT => \N__12014\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12016\,
            PADOUT => \N__12015\,
            PADIN => \N__12014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12007\,
            DIN => \N__12006\,
            DOUT => \N__12005\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12007\,
            PADOUT => \N__12006\,
            PADIN => \N__12005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8614\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11998\,
            DIN => \N__11997\,
            DOUT => \N__11996\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11998\,
            PADOUT => \N__11997\,
            PADIN => \N__11996\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7932\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11989\,
            DIN => \N__11988\,
            DOUT => \N__11987\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11989\,
            PADOUT => \N__11988\,
            PADIN => \N__11987\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5457\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11980\,
            DIN => \N__11979\,
            DOUT => \N__11978\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11980\,
            PADOUT => \N__11979\,
            PADIN => \N__11978\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4944\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11971\,
            DIN => \N__11970\,
            DOUT => \N__11969\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11971\,
            PADOUT => \N__11970\,
            PADIN => \N__11969\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2915\ : InMux
    port map (
            O => \N__11952\,
            I => \N__11947\
        );

    \I__2914\ : InMux
    port map (
            O => \N__11951\,
            I => \N__11944\
        );

    \I__2913\ : InMux
    port map (
            O => \N__11950\,
            I => \N__11941\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__11947\,
            I => \N__11938\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__11944\,
            I => \N__11933\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__11941\,
            I => \N__11933\
        );

    \I__2909\ : Span4Mux_v
    port map (
            O => \N__11938\,
            I => \N__11928\
        );

    \I__2908\ : Span4Mux_v
    port map (
            O => \N__11933\,
            I => \N__11928\
        );

    \I__2907\ : Span4Mux_v
    port map (
            O => \N__11928\,
            I => \N__11924\
        );

    \I__2906\ : InMux
    port map (
            O => \N__11927\,
            I => \N__11920\
        );

    \I__2905\ : Span4Mux_h
    port map (
            O => \N__11924\,
            I => \N__11916\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__11923\,
            I => \N__11913\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__11920\,
            I => \N__11910\
        );

    \I__2902\ : InMux
    port map (
            O => \N__11919\,
            I => \N__11907\
        );

    \I__2901\ : Span4Mux_h
    port map (
            O => \N__11916\,
            I => \N__11904\
        );

    \I__2900\ : InMux
    port map (
            O => \N__11913\,
            I => \N__11901\
        );

    \I__2899\ : Sp12to4
    port map (
            O => \N__11910\,
            I => \N__11896\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__11907\,
            I => \N__11896\
        );

    \I__2897\ : Span4Mux_h
    port map (
            O => \N__11904\,
            I => \N__11891\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__11901\,
            I => \N__11891\
        );

    \I__2895\ : Span12Mux_v
    port map (
            O => \N__11896\,
            I => \N__11888\
        );

    \I__2894\ : Span4Mux_h
    port map (
            O => \N__11891\,
            I => \N__11885\
        );

    \I__2893\ : Span12Mux_h
    port map (
            O => \N__11888\,
            I => \N__11882\
        );

    \I__2892\ : Span4Mux_v
    port map (
            O => \N__11885\,
            I => \N__11879\
        );

    \I__2891\ : Odrv12
    port map (
            O => \N__11882\,
            I => \CASUn_c\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__11879\,
            I => \CASUn_c\
        );

    \I__2889\ : InMux
    port map (
            O => \N__11874\,
            I => \N__11869\
        );

    \I__2888\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11865\
        );

    \I__2887\ : InMux
    port map (
            O => \N__11872\,
            I => \N__11862\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__11869\,
            I => \N__11859\
        );

    \I__2885\ : InMux
    port map (
            O => \N__11868\,
            I => \N__11856\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__11865\,
            I => \N__11851\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__11862\,
            I => \N__11851\
        );

    \I__2882\ : Span4Mux_v
    port map (
            O => \N__11859\,
            I => \N__11845\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__11856\,
            I => \N__11845\
        );

    \I__2880\ : Span4Mux_h
    port map (
            O => \N__11851\,
            I => \N__11842\
        );

    \I__2879\ : InMux
    port map (
            O => \N__11850\,
            I => \N__11839\
        );

    \I__2878\ : Span4Mux_v
    port map (
            O => \N__11845\,
            I => \N__11836\
        );

    \I__2877\ : Sp12to4
    port map (
            O => \N__11842\,
            I => \N__11830\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__11839\,
            I => \N__11830\
        );

    \I__2875\ : Span4Mux_v
    port map (
            O => \N__11836\,
            I => \N__11827\
        );

    \I__2874\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11824\
        );

    \I__2873\ : Span12Mux_v
    port map (
            O => \N__11830\,
            I => \N__11819\
        );

    \I__2872\ : Sp12to4
    port map (
            O => \N__11827\,
            I => \N__11819\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__11824\,
            I => \N__11816\
        );

    \I__2870\ : Span12Mux_h
    port map (
            O => \N__11819\,
            I => \N__11811\
        );

    \I__2869\ : Span12Mux_v
    port map (
            O => \N__11816\,
            I => \N__11811\
        );

    \I__2868\ : Odrv12
    port map (
            O => \N__11811\,
            I => \CASLn_c\
        );

    \I__2867\ : IoInMux
    port map (
            O => \N__11808\,
            I => \N__11805\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__11805\,
            I => \N__11802\
        );

    \I__2865\ : Span4Mux_s3_h
    port map (
            O => \N__11802\,
            I => \N__11799\
        );

    \I__2864\ : Span4Mux_v
    port map (
            O => \N__11799\,
            I => \N__11796\
        );

    \I__2863\ : Odrv4
    port map (
            O => \N__11796\,
            I => \DRDDIR_c\
        );

    \I__2862\ : InMux
    port map (
            O => \N__11793\,
            I => \N__11787\
        );

    \I__2861\ : InMux
    port map (
            O => \N__11792\,
            I => \N__11787\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__11787\,
            I => \N__11784\
        );

    \I__2859\ : Span4Mux_h
    port map (
            O => \N__11784\,
            I => \N__11781\
        );

    \I__2858\ : Odrv4
    port map (
            O => \N__11781\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2857\ : InMux
    port map (
            O => \N__11778\,
            I => \N__11774\
        );

    \I__2856\ : InMux
    port map (
            O => \N__11777\,
            I => \N__11771\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__11774\,
            I => \N__11768\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__11771\,
            I => \N__11763\
        );

    \I__2853\ : Span4Mux_v
    port map (
            O => \N__11768\,
            I => \N__11760\
        );

    \I__2852\ : InMux
    port map (
            O => \N__11767\,
            I => \N__11755\
        );

    \I__2851\ : InMux
    port map (
            O => \N__11766\,
            I => \N__11755\
        );

    \I__2850\ : Span4Mux_v
    port map (
            O => \N__11763\,
            I => \N__11752\
        );

    \I__2849\ : Sp12to4
    port map (
            O => \N__11760\,
            I => \N__11747\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__11755\,
            I => \N__11747\
        );

    \I__2847\ : Sp12to4
    port map (
            O => \N__11752\,
            I => \N__11744\
        );

    \I__2846\ : Span12Mux_h
    port map (
            O => \N__11747\,
            I => \N__11741\
        );

    \I__2845\ : Span12Mux_h
    port map (
            O => \N__11744\,
            I => \N__11738\
        );

    \I__2844\ : Odrv12
    port map (
            O => \N__11741\,
            I => \DRA_c_7\
        );

    \I__2843\ : Odrv12
    port map (
            O => \N__11738\,
            I => \DRA_c_7\
        );

    \I__2842\ : InMux
    port map (
            O => \N__11733\,
            I => \N__11727\
        );

    \I__2841\ : InMux
    port map (
            O => \N__11732\,
            I => \N__11724\
        );

    \I__2840\ : InMux
    port map (
            O => \N__11731\,
            I => \N__11721\
        );

    \I__2839\ : InMux
    port map (
            O => \N__11730\,
            I => \N__11718\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__11727\,
            I => \N__11715\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__11724\,
            I => \N__11712\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__11721\,
            I => \N__11707\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__11718\,
            I => \N__11707\
        );

    \I__2834\ : Span4Mux_v
    port map (
            O => \N__11715\,
            I => \N__11702\
        );

    \I__2833\ : Span4Mux_v
    port map (
            O => \N__11712\,
            I => \N__11702\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__11707\,
            I => \N__11699\
        );

    \I__2831\ : Span4Mux_h
    port map (
            O => \N__11702\,
            I => \N__11696\
        );

    \I__2830\ : Span4Mux_h
    port map (
            O => \N__11699\,
            I => \N__11693\
        );

    \I__2829\ : Sp12to4
    port map (
            O => \N__11696\,
            I => \N__11688\
        );

    \I__2828\ : Sp12to4
    port map (
            O => \N__11693\,
            I => \N__11688\
        );

    \I__2827\ : Odrv12
    port map (
            O => \N__11688\,
            I => \DRA_c_8\
        );

    \I__2826\ : InMux
    port map (
            O => \N__11685\,
            I => \N__11682\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__11682\,
            I => \N__11679\
        );

    \I__2824\ : Span4Mux_v
    port map (
            O => \N__11679\,
            I => \N__11676\
        );

    \I__2823\ : Odrv4
    port map (
            O => \N__11676\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2822\ : InMux
    port map (
            O => \N__11673\,
            I => \N__11670\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__11670\,
            I => \N__11664\
        );

    \I__2820\ : InMux
    port map (
            O => \N__11669\,
            I => \N__11661\
        );

    \I__2819\ : InMux
    port map (
            O => \N__11668\,
            I => \N__11658\
        );

    \I__2818\ : InMux
    port map (
            O => \N__11667\,
            I => \N__11655\
        );

    \I__2817\ : Span4Mux_h
    port map (
            O => \N__11664\,
            I => \N__11650\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__11661\,
            I => \N__11650\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__11658\,
            I => \N__11647\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__11655\,
            I => \N__11642\
        );

    \I__2813\ : Sp12to4
    port map (
            O => \N__11650\,
            I => \N__11642\
        );

    \I__2812\ : Span4Mux_h
    port map (
            O => \N__11647\,
            I => \N__11639\
        );

    \I__2811\ : Span12Mux_v
    port map (
            O => \N__11642\,
            I => \N__11636\
        );

    \I__2810\ : Span4Mux_v
    port map (
            O => \N__11639\,
            I => \N__11633\
        );

    \I__2809\ : Span12Mux_h
    port map (
            O => \N__11636\,
            I => \N__11630\
        );

    \I__2808\ : Sp12to4
    port map (
            O => \N__11633\,
            I => \N__11627\
        );

    \I__2807\ : Odrv12
    port map (
            O => \N__11630\,
            I => \DRA_c_3\
        );

    \I__2806\ : Odrv12
    port map (
            O => \N__11627\,
            I => \DRA_c_3\
        );

    \I__2805\ : InMux
    port map (
            O => \N__11622\,
            I => \N__11619\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__11619\,
            I => \N__11615\
        );

    \I__2803\ : InMux
    port map (
            O => \N__11618\,
            I => \N__11612\
        );

    \I__2802\ : Span4Mux_v
    port map (
            O => \N__11615\,
            I => \N__11605\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__11612\,
            I => \N__11605\
        );

    \I__2800\ : InMux
    port map (
            O => \N__11611\,
            I => \N__11602\
        );

    \I__2799\ : InMux
    port map (
            O => \N__11610\,
            I => \N__11599\
        );

    \I__2798\ : Span4Mux_v
    port map (
            O => \N__11605\,
            I => \N__11596\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__11602\,
            I => \N__11593\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__11599\,
            I => \N__11590\
        );

    \I__2795\ : Span4Mux_v
    port map (
            O => \N__11596\,
            I => \N__11587\
        );

    \I__2794\ : Span4Mux_h
    port map (
            O => \N__11593\,
            I => \N__11584\
        );

    \I__2793\ : Span12Mux_v
    port map (
            O => \N__11590\,
            I => \N__11579\
        );

    \I__2792\ : Sp12to4
    port map (
            O => \N__11587\,
            I => \N__11579\
        );

    \I__2791\ : Sp12to4
    port map (
            O => \N__11584\,
            I => \N__11576\
        );

    \I__2790\ : Span12Mux_h
    port map (
            O => \N__11579\,
            I => \N__11573\
        );

    \I__2789\ : Span12Mux_v
    port map (
            O => \N__11576\,
            I => \N__11570\
        );

    \I__2788\ : Odrv12
    port map (
            O => \N__11573\,
            I => \DRA_c_2\
        );

    \I__2787\ : Odrv12
    port map (
            O => \N__11570\,
            I => \DRA_c_2\
        );

    \I__2786\ : InMux
    port map (
            O => \N__11565\,
            I => \N__11562\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__11562\,
            I => \N__11559\
        );

    \I__2784\ : Span4Mux_h
    port map (
            O => \N__11559\,
            I => \N__11556\
        );

    \I__2783\ : Odrv4
    port map (
            O => \N__11556\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__11553\,
            I => \N__11549\
        );

    \I__2781\ : InMux
    port map (
            O => \N__11552\,
            I => \N__11545\
        );

    \I__2780\ : InMux
    port map (
            O => \N__11549\,
            I => \N__11540\
        );

    \I__2779\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11540\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__11545\,
            I => \N__11536\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__11540\,
            I => \N__11525\
        );

    \I__2776\ : InMux
    port map (
            O => \N__11539\,
            I => \N__11522\
        );

    \I__2775\ : Span4Mux_v
    port map (
            O => \N__11536\,
            I => \N__11519\
        );

    \I__2774\ : InMux
    port map (
            O => \N__11535\,
            I => \N__11516\
        );

    \I__2773\ : InMux
    port map (
            O => \N__11534\,
            I => \N__11513\
        );

    \I__2772\ : InMux
    port map (
            O => \N__11533\,
            I => \N__11510\
        );

    \I__2771\ : InMux
    port map (
            O => \N__11532\,
            I => \N__11507\
        );

    \I__2770\ : InMux
    port map (
            O => \N__11531\,
            I => \N__11504\
        );

    \I__2769\ : InMux
    port map (
            O => \N__11530\,
            I => \N__11501\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__11529\,
            I => \N__11497\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__11528\,
            I => \N__11491\
        );

    \I__2766\ : Span4Mux_v
    port map (
            O => \N__11525\,
            I => \N__11487\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__11522\,
            I => \N__11484\
        );

    \I__2764\ : Span4Mux_h
    port map (
            O => \N__11519\,
            I => \N__11481\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__11516\,
            I => \N__11472\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__11513\,
            I => \N__11472\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__11510\,
            I => \N__11472\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__11507\,
            I => \N__11472\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__11504\,
            I => \N__11467\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__11501\,
            I => \N__11464\
        );

    \I__2757\ : InMux
    port map (
            O => \N__11500\,
            I => \N__11455\
        );

    \I__2756\ : InMux
    port map (
            O => \N__11497\,
            I => \N__11455\
        );

    \I__2755\ : InMux
    port map (
            O => \N__11496\,
            I => \N__11455\
        );

    \I__2754\ : InMux
    port map (
            O => \N__11495\,
            I => \N__11455\
        );

    \I__2753\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11452\
        );

    \I__2752\ : InMux
    port map (
            O => \N__11491\,
            I => \N__11447\
        );

    \I__2751\ : InMux
    port map (
            O => \N__11490\,
            I => \N__11447\
        );

    \I__2750\ : Span4Mux_h
    port map (
            O => \N__11487\,
            I => \N__11440\
        );

    \I__2749\ : Span4Mux_v
    port map (
            O => \N__11484\,
            I => \N__11440\
        );

    \I__2748\ : Span4Mux_h
    port map (
            O => \N__11481\,
            I => \N__11435\
        );

    \I__2747\ : Span4Mux_v
    port map (
            O => \N__11472\,
            I => \N__11435\
        );

    \I__2746\ : InMux
    port map (
            O => \N__11471\,
            I => \N__11430\
        );

    \I__2745\ : InMux
    port map (
            O => \N__11470\,
            I => \N__11430\
        );

    \I__2744\ : Span4Mux_h
    port map (
            O => \N__11467\,
            I => \N__11419\
        );

    \I__2743\ : Span4Mux_h
    port map (
            O => \N__11464\,
            I => \N__11419\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__11455\,
            I => \N__11419\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__11452\,
            I => \N__11419\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__11447\,
            I => \N__11419\
        );

    \I__2739\ : InMux
    port map (
            O => \N__11446\,
            I => \N__11414\
        );

    \I__2738\ : InMux
    port map (
            O => \N__11445\,
            I => \N__11414\
        );

    \I__2737\ : Sp12to4
    port map (
            O => \N__11440\,
            I => \N__11409\
        );

    \I__2736\ : Sp12to4
    port map (
            O => \N__11435\,
            I => \N__11409\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__11430\,
            I => \N__11406\
        );

    \I__2734\ : Sp12to4
    port map (
            O => \N__11419\,
            I => \N__11403\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__11414\,
            I => \N__11400\
        );

    \I__2732\ : Span12Mux_h
    port map (
            O => \N__11409\,
            I => \N__11397\
        );

    \I__2731\ : Span12Mux_v
    port map (
            O => \N__11406\,
            I => \N__11394\
        );

    \I__2730\ : Span12Mux_v
    port map (
            O => \N__11403\,
            I => \N__11391\
        );

    \I__2729\ : Span12Mux_h
    port map (
            O => \N__11400\,
            I => \N__11388\
        );

    \I__2728\ : Span12Mux_v
    port map (
            O => \N__11397\,
            I => \N__11383\
        );

    \I__2727\ : Span12Mux_h
    port map (
            O => \N__11394\,
            I => \N__11383\
        );

    \I__2726\ : Span12Mux_h
    port map (
            O => \N__11391\,
            I => \N__11378\
        );

    \I__2725\ : Span12Mux_v
    port map (
            O => \N__11388\,
            I => \N__11378\
        );

    \I__2724\ : Odrv12
    port map (
            O => \N__11383\,
            I => \AGNUS_REV_c\
        );

    \I__2723\ : Odrv12
    port map (
            O => \N__11378\,
            I => \AGNUS_REV_c\
        );

    \I__2722\ : InMux
    port map (
            O => \N__11373\,
            I => \N__11368\
        );

    \I__2721\ : InMux
    port map (
            O => \N__11372\,
            I => \N__11365\
        );

    \I__2720\ : InMux
    port map (
            O => \N__11371\,
            I => \N__11361\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__11368\,
            I => \N__11358\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__11365\,
            I => \N__11355\
        );

    \I__2717\ : InMux
    port map (
            O => \N__11364\,
            I => \N__11352\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__11361\,
            I => \N__11349\
        );

    \I__2715\ : Span4Mux_v
    port map (
            O => \N__11358\,
            I => \N__11346\
        );

    \I__2714\ : Span4Mux_v
    port map (
            O => \N__11355\,
            I => \N__11339\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__11352\,
            I => \N__11339\
        );

    \I__2712\ : Span4Mux_v
    port map (
            O => \N__11349\,
            I => \N__11339\
        );

    \I__2711\ : Sp12to4
    port map (
            O => \N__11346\,
            I => \N__11334\
        );

    \I__2710\ : Sp12to4
    port map (
            O => \N__11339\,
            I => \N__11334\
        );

    \I__2709\ : Span12Mux_h
    port map (
            O => \N__11334\,
            I => \N__11331\
        );

    \I__2708\ : Span12Mux_v
    port map (
            O => \N__11331\,
            I => \N__11328\
        );

    \I__2707\ : Odrv12
    port map (
            O => \N__11328\,
            I => \DRA_c_1\
        );

    \I__2706\ : InMux
    port map (
            O => \N__11325\,
            I => \N__11322\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__11322\,
            I => \N__11318\
        );

    \I__2704\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11315\
        );

    \I__2703\ : Span4Mux_h
    port map (
            O => \N__11318\,
            I => \N__11310\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__11315\,
            I => \N__11310\
        );

    \I__2701\ : Sp12to4
    port map (
            O => \N__11310\,
            I => \N__11307\
        );

    \I__2700\ : Span12Mux_v
    port map (
            O => \N__11307\,
            I => \N__11304\
        );

    \I__2699\ : Span12Mux_h
    port map (
            O => \N__11304\,
            I => \N__11301\
        );

    \I__2698\ : Odrv12
    port map (
            O => \N__11301\,
            I => \DRA_c_0\
        );

    \I__2697\ : InMux
    port map (
            O => \N__11298\,
            I => \N__11295\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__11295\,
            I => \N__11292\
        );

    \I__2695\ : Span4Mux_h
    port map (
            O => \N__11292\,
            I => \N__11289\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__11289\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2693\ : ClkMux
    port map (
            O => \N__11286\,
            I => \N__11268\
        );

    \I__2692\ : ClkMux
    port map (
            O => \N__11285\,
            I => \N__11268\
        );

    \I__2691\ : ClkMux
    port map (
            O => \N__11284\,
            I => \N__11268\
        );

    \I__2690\ : ClkMux
    port map (
            O => \N__11283\,
            I => \N__11268\
        );

    \I__2689\ : ClkMux
    port map (
            O => \N__11282\,
            I => \N__11268\
        );

    \I__2688\ : ClkMux
    port map (
            O => \N__11281\,
            I => \N__11268\
        );

    \I__2687\ : GlobalMux
    port map (
            O => \N__11268\,
            I => \N__11265\
        );

    \I__2686\ : gio2CtrlBuf
    port map (
            O => \N__11265\,
            I => \C3_c_g\
        );

    \I__2685\ : CEMux
    port map (
            O => \N__11262\,
            I => \N__11226\
        );

    \I__2684\ : CEMux
    port map (
            O => \N__11261\,
            I => \N__11226\
        );

    \I__2683\ : CEMux
    port map (
            O => \N__11260\,
            I => \N__11226\
        );

    \I__2682\ : CEMux
    port map (
            O => \N__11259\,
            I => \N__11226\
        );

    \I__2681\ : CEMux
    port map (
            O => \N__11258\,
            I => \N__11226\
        );

    \I__2680\ : CEMux
    port map (
            O => \N__11257\,
            I => \N__11226\
        );

    \I__2679\ : CEMux
    port map (
            O => \N__11256\,
            I => \N__11226\
        );

    \I__2678\ : CEMux
    port map (
            O => \N__11255\,
            I => \N__11226\
        );

    \I__2677\ : CEMux
    port map (
            O => \N__11254\,
            I => \N__11226\
        );

    \I__2676\ : CEMux
    port map (
            O => \N__11253\,
            I => \N__11226\
        );

    \I__2675\ : CEMux
    port map (
            O => \N__11252\,
            I => \N__11226\
        );

    \I__2674\ : CEMux
    port map (
            O => \N__11251\,
            I => \N__11226\
        );

    \I__2673\ : GlobalMux
    port map (
            O => \N__11226\,
            I => \N__11223\
        );

    \I__2672\ : gio2CtrlBuf
    port map (
            O => \N__11223\,
            I => \DBRn_c_i_0_g\
        );

    \I__2671\ : InMux
    port map (
            O => \N__11220\,
            I => \N__11213\
        );

    \I__2670\ : InMux
    port map (
            O => \N__11219\,
            I => \N__11210\
        );

    \I__2669\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11207\
        );

    \I__2668\ : InMux
    port map (
            O => \N__11217\,
            I => \N__11204\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11216\,
            I => \N__11201\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__11213\,
            I => \N__11198\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__11210\,
            I => \N__11181\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__11207\,
            I => \N__11178\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__11204\,
            I => \N__11164\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__11201\,
            I => \N__11151\
        );

    \I__2661\ : Glb2LocalMux
    port map (
            O => \N__11198\,
            I => \N__11064\
        );

    \I__2660\ : SRMux
    port map (
            O => \N__11197\,
            I => \N__11064\
        );

    \I__2659\ : SRMux
    port map (
            O => \N__11196\,
            I => \N__11064\
        );

    \I__2658\ : SRMux
    port map (
            O => \N__11195\,
            I => \N__11064\
        );

    \I__2657\ : SRMux
    port map (
            O => \N__11194\,
            I => \N__11064\
        );

    \I__2656\ : SRMux
    port map (
            O => \N__11193\,
            I => \N__11064\
        );

    \I__2655\ : SRMux
    port map (
            O => \N__11192\,
            I => \N__11064\
        );

    \I__2654\ : SRMux
    port map (
            O => \N__11191\,
            I => \N__11064\
        );

    \I__2653\ : SRMux
    port map (
            O => \N__11190\,
            I => \N__11064\
        );

    \I__2652\ : SRMux
    port map (
            O => \N__11189\,
            I => \N__11064\
        );

    \I__2651\ : SRMux
    port map (
            O => \N__11188\,
            I => \N__11064\
        );

    \I__2650\ : SRMux
    port map (
            O => \N__11187\,
            I => \N__11064\
        );

    \I__2649\ : SRMux
    port map (
            O => \N__11186\,
            I => \N__11064\
        );

    \I__2648\ : SRMux
    port map (
            O => \N__11185\,
            I => \N__11064\
        );

    \I__2647\ : SRMux
    port map (
            O => \N__11184\,
            I => \N__11064\
        );

    \I__2646\ : Glb2LocalMux
    port map (
            O => \N__11181\,
            I => \N__11064\
        );

    \I__2645\ : Glb2LocalMux
    port map (
            O => \N__11178\,
            I => \N__11064\
        );

    \I__2644\ : SRMux
    port map (
            O => \N__11177\,
            I => \N__11064\
        );

    \I__2643\ : SRMux
    port map (
            O => \N__11176\,
            I => \N__11064\
        );

    \I__2642\ : SRMux
    port map (
            O => \N__11175\,
            I => \N__11064\
        );

    \I__2641\ : SRMux
    port map (
            O => \N__11174\,
            I => \N__11064\
        );

    \I__2640\ : SRMux
    port map (
            O => \N__11173\,
            I => \N__11064\
        );

    \I__2639\ : SRMux
    port map (
            O => \N__11172\,
            I => \N__11064\
        );

    \I__2638\ : SRMux
    port map (
            O => \N__11171\,
            I => \N__11064\
        );

    \I__2637\ : SRMux
    port map (
            O => \N__11170\,
            I => \N__11064\
        );

    \I__2636\ : SRMux
    port map (
            O => \N__11169\,
            I => \N__11064\
        );

    \I__2635\ : SRMux
    port map (
            O => \N__11168\,
            I => \N__11064\
        );

    \I__2634\ : SRMux
    port map (
            O => \N__11167\,
            I => \N__11064\
        );

    \I__2633\ : Glb2LocalMux
    port map (
            O => \N__11164\,
            I => \N__11064\
        );

    \I__2632\ : SRMux
    port map (
            O => \N__11163\,
            I => \N__11064\
        );

    \I__2631\ : SRMux
    port map (
            O => \N__11162\,
            I => \N__11064\
        );

    \I__2630\ : SRMux
    port map (
            O => \N__11161\,
            I => \N__11064\
        );

    \I__2629\ : SRMux
    port map (
            O => \N__11160\,
            I => \N__11064\
        );

    \I__2628\ : SRMux
    port map (
            O => \N__11159\,
            I => \N__11064\
        );

    \I__2627\ : SRMux
    port map (
            O => \N__11158\,
            I => \N__11064\
        );

    \I__2626\ : SRMux
    port map (
            O => \N__11157\,
            I => \N__11064\
        );

    \I__2625\ : SRMux
    port map (
            O => \N__11156\,
            I => \N__11064\
        );

    \I__2624\ : SRMux
    port map (
            O => \N__11155\,
            I => \N__11064\
        );

    \I__2623\ : SRMux
    port map (
            O => \N__11154\,
            I => \N__11064\
        );

    \I__2622\ : Glb2LocalMux
    port map (
            O => \N__11151\,
            I => \N__11064\
        );

    \I__2621\ : SRMux
    port map (
            O => \N__11150\,
            I => \N__11064\
        );

    \I__2620\ : SRMux
    port map (
            O => \N__11149\,
            I => \N__11064\
        );

    \I__2619\ : GlobalMux
    port map (
            O => \N__11064\,
            I => \N__11061\
        );

    \I__2618\ : gio2CtrlBuf
    port map (
            O => \N__11061\,
            I => \RESETn_c_i_g\
        );

    \I__2617\ : InMux
    port map (
            O => \N__11058\,
            I => \N__11055\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__11055\,
            I => \N__11052\
        );

    \I__2615\ : Span12Mux_v
    port map (
            O => \N__11052\,
            I => \N__11049\
        );

    \I__2614\ : Span12Mux_h
    port map (
            O => \N__11049\,
            I => \N__11046\
        );

    \I__2613\ : Odrv12
    port map (
            O => \N__11046\,
            I => \RAS1n_c\
        );

    \I__2612\ : InMux
    port map (
            O => \N__11043\,
            I => \N__11039\
        );

    \I__2611\ : InMux
    port map (
            O => \N__11042\,
            I => \N__11036\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__11039\,
            I => \N__11033\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__11036\,
            I => \N__11030\
        );

    \I__2608\ : Span4Mux_v
    port map (
            O => \N__11033\,
            I => \N__11027\
        );

    \I__2607\ : Span12Mux_h
    port map (
            O => \N__11030\,
            I => \N__11024\
        );

    \I__2606\ : Sp12to4
    port map (
            O => \N__11027\,
            I => \N__11021\
        );

    \I__2605\ : Odrv12
    port map (
            O => \N__11024\,
            I => \RAS0n_c\
        );

    \I__2604\ : Odrv12
    port map (
            O => \N__11021\,
            I => \RAS0n_c\
        );

    \I__2603\ : InMux
    port map (
            O => \N__11016\,
            I => \N__11013\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__11013\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2601\ : InMux
    port map (
            O => \N__11010\,
            I => \N__10993\
        );

    \I__2600\ : InMux
    port map (
            O => \N__11009\,
            I => \N__10990\
        );

    \I__2599\ : InMux
    port map (
            O => \N__11008\,
            I => \N__10987\
        );

    \I__2598\ : InMux
    port map (
            O => \N__11007\,
            I => \N__10982\
        );

    \I__2597\ : InMux
    port map (
            O => \N__11006\,
            I => \N__10982\
        );

    \I__2596\ : InMux
    port map (
            O => \N__11005\,
            I => \N__10977\
        );

    \I__2595\ : InMux
    port map (
            O => \N__11004\,
            I => \N__10977\
        );

    \I__2594\ : InMux
    port map (
            O => \N__11003\,
            I => \N__10972\
        );

    \I__2593\ : InMux
    port map (
            O => \N__11002\,
            I => \N__10972\
        );

    \I__2592\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10969\
        );

    \I__2591\ : InMux
    port map (
            O => \N__11000\,
            I => \N__10966\
        );

    \I__2590\ : InMux
    port map (
            O => \N__10999\,
            I => \N__10963\
        );

    \I__2589\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10949\
        );

    \I__2588\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10949\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__10996\,
            I => \N__10944\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__10993\,
            I => \N__10938\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__10990\,
            I => \N__10923\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__10987\,
            I => \N__10923\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__10982\,
            I => \N__10923\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__10977\,
            I => \N__10923\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__10972\,
            I => \N__10923\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__10969\,
            I => \N__10923\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__10966\,
            I => \N__10923\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__10963\,
            I => \N__10920\
        );

    \I__2577\ : InMux
    port map (
            O => \N__10962\,
            I => \N__10917\
        );

    \I__2576\ : InMux
    port map (
            O => \N__10961\,
            I => \N__10914\
        );

    \I__2575\ : InMux
    port map (
            O => \N__10960\,
            I => \N__10909\
        );

    \I__2574\ : InMux
    port map (
            O => \N__10959\,
            I => \N__10909\
        );

    \I__2573\ : InMux
    port map (
            O => \N__10958\,
            I => \N__10902\
        );

    \I__2572\ : InMux
    port map (
            O => \N__10957\,
            I => \N__10902\
        );

    \I__2571\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10902\
        );

    \I__2570\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10897\
        );

    \I__2569\ : InMux
    port map (
            O => \N__10954\,
            I => \N__10897\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__10949\,
            I => \N__10894\
        );

    \I__2567\ : InMux
    port map (
            O => \N__10948\,
            I => \N__10891\
        );

    \I__2566\ : InMux
    port map (
            O => \N__10947\,
            I => \N__10888\
        );

    \I__2565\ : InMux
    port map (
            O => \N__10944\,
            I => \N__10881\
        );

    \I__2564\ : InMux
    port map (
            O => \N__10943\,
            I => \N__10881\
        );

    \I__2563\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10881\
        );

    \I__2562\ : InMux
    port map (
            O => \N__10941\,
            I => \N__10878\
        );

    \I__2561\ : Span4Mux_v
    port map (
            O => \N__10938\,
            I => \N__10870\
        );

    \I__2560\ : Span4Mux_v
    port map (
            O => \N__10923\,
            I => \N__10870\
        );

    \I__2559\ : Span4Mux_v
    port map (
            O => \N__10920\,
            I => \N__10863\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__10917\,
            I => \N__10863\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__10914\,
            I => \N__10863\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__10909\,
            I => \N__10860\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__10902\,
            I => \N__10855\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__10897\,
            I => \N__10855\
        );

    \I__2553\ : Span4Mux_v
    port map (
            O => \N__10894\,
            I => \N__10844\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10891\,
            I => \N__10844\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__10888\,
            I => \N__10844\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__10881\,
            I => \N__10844\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__10878\,
            I => \N__10844\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__10877\,
            I => \N__10841\
        );

    \I__2547\ : InMux
    port map (
            O => \N__10876\,
            I => \N__10835\
        );

    \I__2546\ : InMux
    port map (
            O => \N__10875\,
            I => \N__10835\
        );

    \I__2545\ : Span4Mux_h
    port map (
            O => \N__10870\,
            I => \N__10829\
        );

    \I__2544\ : Span4Mux_v
    port map (
            O => \N__10863\,
            I => \N__10829\
        );

    \I__2543\ : Span4Mux_v
    port map (
            O => \N__10860\,
            I => \N__10822\
        );

    \I__2542\ : Span4Mux_h
    port map (
            O => \N__10855\,
            I => \N__10822\
        );

    \I__2541\ : Span4Mux_v
    port map (
            O => \N__10844\,
            I => \N__10822\
        );

    \I__2540\ : InMux
    port map (
            O => \N__10841\,
            I => \N__10819\
        );

    \I__2539\ : InMux
    port map (
            O => \N__10840\,
            I => \N__10816\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__10835\,
            I => \N__10813\
        );

    \I__2537\ : InMux
    port map (
            O => \N__10834\,
            I => \N__10810\
        );

    \I__2536\ : Sp12to4
    port map (
            O => \N__10829\,
            I => \N__10801\
        );

    \I__2535\ : Sp12to4
    port map (
            O => \N__10822\,
            I => \N__10801\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__10819\,
            I => \N__10801\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__10816\,
            I => \N__10801\
        );

    \I__2532\ : Span12Mux_v
    port map (
            O => \N__10813\,
            I => \N__10796\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__10810\,
            I => \N__10796\
        );

    \I__2530\ : Span12Mux_h
    port map (
            O => \N__10801\,
            I => \N__10793\
        );

    \I__2529\ : Span12Mux_h
    port map (
            O => \N__10796\,
            I => \N__10790\
        );

    \I__2528\ : Odrv12
    port map (
            O => \N__10793\,
            I => \RESETn_c\
        );

    \I__2527\ : Odrv12
    port map (
            O => \N__10790\,
            I => \RESETn_c\
        );

    \I__2526\ : InMux
    port map (
            O => \N__10785\,
            I => \N__10782\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__10782\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__2524\ : InMux
    port map (
            O => \N__10779\,
            I => \N__10776\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__10776\,
            I => \N__10773\
        );

    \I__2522\ : Odrv12
    port map (
            O => \N__10773\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\
        );

    \I__2521\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10767\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__10767\,
            I => \N__10725\
        );

    \I__2519\ : ClkMux
    port map (
            O => \N__10766\,
            I => \N__10623\
        );

    \I__2518\ : ClkMux
    port map (
            O => \N__10765\,
            I => \N__10623\
        );

    \I__2517\ : ClkMux
    port map (
            O => \N__10764\,
            I => \N__10623\
        );

    \I__2516\ : ClkMux
    port map (
            O => \N__10763\,
            I => \N__10623\
        );

    \I__2515\ : ClkMux
    port map (
            O => \N__10762\,
            I => \N__10623\
        );

    \I__2514\ : ClkMux
    port map (
            O => \N__10761\,
            I => \N__10623\
        );

    \I__2513\ : ClkMux
    port map (
            O => \N__10760\,
            I => \N__10623\
        );

    \I__2512\ : ClkMux
    port map (
            O => \N__10759\,
            I => \N__10623\
        );

    \I__2511\ : ClkMux
    port map (
            O => \N__10758\,
            I => \N__10623\
        );

    \I__2510\ : ClkMux
    port map (
            O => \N__10757\,
            I => \N__10623\
        );

    \I__2509\ : ClkMux
    port map (
            O => \N__10756\,
            I => \N__10623\
        );

    \I__2508\ : ClkMux
    port map (
            O => \N__10755\,
            I => \N__10623\
        );

    \I__2507\ : ClkMux
    port map (
            O => \N__10754\,
            I => \N__10623\
        );

    \I__2506\ : ClkMux
    port map (
            O => \N__10753\,
            I => \N__10623\
        );

    \I__2505\ : ClkMux
    port map (
            O => \N__10752\,
            I => \N__10623\
        );

    \I__2504\ : ClkMux
    port map (
            O => \N__10751\,
            I => \N__10623\
        );

    \I__2503\ : ClkMux
    port map (
            O => \N__10750\,
            I => \N__10623\
        );

    \I__2502\ : ClkMux
    port map (
            O => \N__10749\,
            I => \N__10623\
        );

    \I__2501\ : ClkMux
    port map (
            O => \N__10748\,
            I => \N__10623\
        );

    \I__2500\ : ClkMux
    port map (
            O => \N__10747\,
            I => \N__10623\
        );

    \I__2499\ : ClkMux
    port map (
            O => \N__10746\,
            I => \N__10623\
        );

    \I__2498\ : ClkMux
    port map (
            O => \N__10745\,
            I => \N__10623\
        );

    \I__2497\ : ClkMux
    port map (
            O => \N__10744\,
            I => \N__10623\
        );

    \I__2496\ : ClkMux
    port map (
            O => \N__10743\,
            I => \N__10623\
        );

    \I__2495\ : ClkMux
    port map (
            O => \N__10742\,
            I => \N__10623\
        );

    \I__2494\ : ClkMux
    port map (
            O => \N__10741\,
            I => \N__10623\
        );

    \I__2493\ : ClkMux
    port map (
            O => \N__10740\,
            I => \N__10623\
        );

    \I__2492\ : ClkMux
    port map (
            O => \N__10739\,
            I => \N__10623\
        );

    \I__2491\ : ClkMux
    port map (
            O => \N__10738\,
            I => \N__10623\
        );

    \I__2490\ : ClkMux
    port map (
            O => \N__10737\,
            I => \N__10623\
        );

    \I__2489\ : ClkMux
    port map (
            O => \N__10736\,
            I => \N__10623\
        );

    \I__2488\ : ClkMux
    port map (
            O => \N__10735\,
            I => \N__10623\
        );

    \I__2487\ : ClkMux
    port map (
            O => \N__10734\,
            I => \N__10623\
        );

    \I__2486\ : ClkMux
    port map (
            O => \N__10733\,
            I => \N__10623\
        );

    \I__2485\ : ClkMux
    port map (
            O => \N__10732\,
            I => \N__10623\
        );

    \I__2484\ : ClkMux
    port map (
            O => \N__10731\,
            I => \N__10623\
        );

    \I__2483\ : ClkMux
    port map (
            O => \N__10730\,
            I => \N__10623\
        );

    \I__2482\ : ClkMux
    port map (
            O => \N__10729\,
            I => \N__10623\
        );

    \I__2481\ : ClkMux
    port map (
            O => \N__10728\,
            I => \N__10623\
        );

    \I__2480\ : Glb2LocalMux
    port map (
            O => \N__10725\,
            I => \N__10623\
        );

    \I__2479\ : ClkMux
    port map (
            O => \N__10724\,
            I => \N__10623\
        );

    \I__2478\ : ClkMux
    port map (
            O => \N__10723\,
            I => \N__10623\
        );

    \I__2477\ : ClkMux
    port map (
            O => \N__10722\,
            I => \N__10623\
        );

    \I__2476\ : ClkMux
    port map (
            O => \N__10721\,
            I => \N__10623\
        );

    \I__2475\ : ClkMux
    port map (
            O => \N__10720\,
            I => \N__10623\
        );

    \I__2474\ : ClkMux
    port map (
            O => \N__10719\,
            I => \N__10623\
        );

    \I__2473\ : ClkMux
    port map (
            O => \N__10718\,
            I => \N__10623\
        );

    \I__2472\ : GlobalMux
    port map (
            O => \N__10623\,
            I => \CLK80_PLL\
        );

    \I__2471\ : InMux
    port map (
            O => \N__10620\,
            I => \N__10616\
        );

    \I__2470\ : InMux
    port map (
            O => \N__10619\,
            I => \N__10613\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__10616\,
            I => \N__10610\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__10613\,
            I => \N__10607\
        );

    \I__2467\ : Span12Mux_v
    port map (
            O => \N__10610\,
            I => \N__10604\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__10607\,
            I => \N__10601\
        );

    \I__2465\ : Span12Mux_h
    port map (
            O => \N__10604\,
            I => \N__10597\
        );

    \I__2464\ : Span4Mux_v
    port map (
            O => \N__10601\,
            I => \N__10594\
        );

    \I__2463\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10591\
        );

    \I__2462\ : Odrv12
    port map (
            O => \N__10597\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__10594\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__10591\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2459\ : InMux
    port map (
            O => \N__10584\,
            I => \N__10580\
        );

    \I__2458\ : InMux
    port map (
            O => \N__10583\,
            I => \N__10576\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__10580\,
            I => \N__10572\
        );

    \I__2456\ : InMux
    port map (
            O => \N__10579\,
            I => \N__10569\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__10576\,
            I => \N__10566\
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__10575\,
            I => \N__10563\
        );

    \I__2453\ : Span4Mux_v
    port map (
            O => \N__10572\,
            I => \N__10560\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__10569\,
            I => \N__10557\
        );

    \I__2451\ : Span4Mux_v
    port map (
            O => \N__10566\,
            I => \N__10553\
        );

    \I__2450\ : InMux
    port map (
            O => \N__10563\,
            I => \N__10550\
        );

    \I__2449\ : Span4Mux_h
    port map (
            O => \N__10560\,
            I => \N__10545\
        );

    \I__2448\ : Span4Mux_v
    port map (
            O => \N__10557\,
            I => \N__10545\
        );

    \I__2447\ : InMux
    port map (
            O => \N__10556\,
            I => \N__10542\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__10553\,
            I => \N__10539\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__10550\,
            I => \N__10536\
        );

    \I__2444\ : Sp12to4
    port map (
            O => \N__10545\,
            I => \N__10531\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__10542\,
            I => \N__10531\
        );

    \I__2442\ : Sp12to4
    port map (
            O => \N__10539\,
            I => \N__10528\
        );

    \I__2441\ : Sp12to4
    port map (
            O => \N__10536\,
            I => \N__10525\
        );

    \I__2440\ : Span12Mux_h
    port map (
            O => \N__10531\,
            I => \N__10522\
        );

    \I__2439\ : Span12Mux_h
    port map (
            O => \N__10528\,
            I => \N__10517\
        );

    \I__2438\ : Span12Mux_v
    port map (
            O => \N__10525\,
            I => \N__10517\
        );

    \I__2437\ : Span12Mux_v
    port map (
            O => \N__10522\,
            I => \N__10512\
        );

    \I__2436\ : Span12Mux_h
    port map (
            O => \N__10517\,
            I => \N__10512\
        );

    \I__2435\ : Odrv12
    port map (
            O => \N__10512\,
            I => \RnW_c\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10504\
        );

    \I__2433\ : InMux
    port map (
            O => \N__10508\,
            I => \N__10501\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__10507\,
            I => \N__10495\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__10504\,
            I => \N__10492\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__10501\,
            I => \N__10489\
        );

    \I__2429\ : InMux
    port map (
            O => \N__10500\,
            I => \N__10486\
        );

    \I__2428\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10479\
        );

    \I__2427\ : InMux
    port map (
            O => \N__10498\,
            I => \N__10479\
        );

    \I__2426\ : InMux
    port map (
            O => \N__10495\,
            I => \N__10479\
        );

    \I__2425\ : Span4Mux_v
    port map (
            O => \N__10492\,
            I => \N__10471\
        );

    \I__2424\ : Span4Mux_h
    port map (
            O => \N__10489\,
            I => \N__10471\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__10486\,
            I => \N__10471\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__10479\,
            I => \N__10468\
        );

    \I__2421\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10465\
        );

    \I__2420\ : Span4Mux_h
    port map (
            O => \N__10471\,
            I => \N__10460\
        );

    \I__2419\ : Span4Mux_h
    port map (
            O => \N__10468\,
            I => \N__10455\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__10465\,
            I => \N__10455\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10464\,
            I => \N__10450\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10463\,
            I => \N__10450\
        );

    \I__2415\ : Span4Mux_v
    port map (
            O => \N__10460\,
            I => \N__10445\
        );

    \I__2414\ : Span4Mux_h
    port map (
            O => \N__10455\,
            I => \N__10445\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__10450\,
            I => \N__10442\
        );

    \I__2412\ : Span4Mux_v
    port map (
            O => \N__10445\,
            I => \N__10439\
        );

    \I__2411\ : Span12Mux_v
    port map (
            O => \N__10442\,
            I => \N__10436\
        );

    \I__2410\ : Span4Mux_h
    port map (
            O => \N__10439\,
            I => \N__10433\
        );

    \I__2409\ : Span12Mux_h
    port map (
            O => \N__10436\,
            I => \N__10430\
        );

    \I__2408\ : Sp12to4
    port map (
            O => \N__10433\,
            I => \N__10427\
        );

    \I__2407\ : Odrv12
    port map (
            O => \N__10430\,
            I => \SIZ_c_1\
        );

    \I__2406\ : Odrv12
    port map (
            O => \N__10427\,
            I => \SIZ_c_1\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__10422\,
            I => \N__10417\
        );

    \I__2404\ : InMux
    port map (
            O => \N__10421\,
            I => \N__10412\
        );

    \I__2403\ : InMux
    port map (
            O => \N__10420\,
            I => \N__10409\
        );

    \I__2402\ : InMux
    port map (
            O => \N__10417\,
            I => \N__10406\
        );

    \I__2401\ : CascadeMux
    port map (
            O => \N__10416\,
            I => \N__10402\
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__10415\,
            I => \N__10399\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__10412\,
            I => \N__10394\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__10409\,
            I => \N__10391\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__10406\,
            I => \N__10388\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10405\,
            I => \N__10385\
        );

    \I__2395\ : InMux
    port map (
            O => \N__10402\,
            I => \N__10378\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10399\,
            I => \N__10378\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10398\,
            I => \N__10378\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__10397\,
            I => \N__10375\
        );

    \I__2391\ : Span4Mux_v
    port map (
            O => \N__10394\,
            I => \N__10372\
        );

    \I__2390\ : Span4Mux_v
    port map (
            O => \N__10391\,
            I => \N__10365\
        );

    \I__2389\ : Span4Mux_h
    port map (
            O => \N__10388\,
            I => \N__10365\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__10385\,
            I => \N__10365\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__10378\,
            I => \N__10362\
        );

    \I__2386\ : InMux
    port map (
            O => \N__10375\,
            I => \N__10359\
        );

    \I__2385\ : Span4Mux_v
    port map (
            O => \N__10372\,
            I => \N__10356\
        );

    \I__2384\ : Span4Mux_h
    port map (
            O => \N__10365\,
            I => \N__10353\
        );

    \I__2383\ : Span4Mux_h
    port map (
            O => \N__10362\,
            I => \N__10348\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__10359\,
            I => \N__10348\
        );

    \I__2381\ : Span4Mux_v
    port map (
            O => \N__10356\,
            I => \N__10345\
        );

    \I__2380\ : Span4Mux_v
    port map (
            O => \N__10353\,
            I => \N__10340\
        );

    \I__2379\ : Span4Mux_h
    port map (
            O => \N__10348\,
            I => \N__10340\
        );

    \I__2378\ : Span4Mux_h
    port map (
            O => \N__10345\,
            I => \N__10337\
        );

    \I__2377\ : Span4Mux_v
    port map (
            O => \N__10340\,
            I => \N__10334\
        );

    \I__2376\ : Sp12to4
    port map (
            O => \N__10337\,
            I => \N__10329\
        );

    \I__2375\ : Sp12to4
    port map (
            O => \N__10334\,
            I => \N__10329\
        );

    \I__2374\ : Odrv12
    port map (
            O => \N__10329\,
            I => \SIZ_c_0\
        );

    \I__2373\ : IoInMux
    port map (
            O => \N__10326\,
            I => \N__10323\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10323\,
            I => \N__10320\
        );

    \I__2371\ : Span12Mux_s6_v
    port map (
            O => \N__10320\,
            I => \N__10317\
        );

    \I__2370\ : Odrv12
    port map (
            O => \N__10317\,
            I => \N_189\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10314\,
            I => \N__10311\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__10311\,
            I => \N__10308\
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__10308\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10300\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10304\,
            I => \N__10297\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10303\,
            I => \N__10293\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__10300\,
            I => \N__10288\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10297\,
            I => \N__10288\
        );

    \I__2361\ : InMux
    port map (
            O => \N__10296\,
            I => \N__10285\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__10293\,
            I => \N__10282\
        );

    \I__2359\ : Span4Mux_v
    port map (
            O => \N__10288\,
            I => \N__10277\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__10285\,
            I => \N__10277\
        );

    \I__2357\ : Span4Mux_v
    port map (
            O => \N__10282\,
            I => \N__10274\
        );

    \I__2356\ : Span4Mux_h
    port map (
            O => \N__10277\,
            I => \N__10271\
        );

    \I__2355\ : Span4Mux_v
    port map (
            O => \N__10274\,
            I => \N__10268\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__10271\,
            I => \N__10265\
        );

    \I__2353\ : Sp12to4
    port map (
            O => \N__10268\,
            I => \N__10260\
        );

    \I__2352\ : Sp12to4
    port map (
            O => \N__10265\,
            I => \N__10260\
        );

    \I__2351\ : Span12Mux_h
    port map (
            O => \N__10260\,
            I => \N__10257\
        );

    \I__2350\ : Odrv12
    port map (
            O => \N__10257\,
            I => \DRA_c_4\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__10254\,
            I => \N__10251\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10251\,
            I => \N__10248\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__10248\,
            I => \N__10245\
        );

    \I__2346\ : Odrv12
    port map (
            O => \N__10245\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2345\ : InMux
    port map (
            O => \N__10242\,
            I => \N__10235\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10241\,
            I => \N__10235\
        );

    \I__2343\ : InMux
    port map (
            O => \N__10240\,
            I => \N__10232\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__10235\,
            I => \N__10226\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__10232\,
            I => \N__10226\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10223\
        );

    \I__2339\ : Span4Mux_v
    port map (
            O => \N__10226\,
            I => \N__10220\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__10223\,
            I => \N__10217\
        );

    \I__2337\ : Sp12to4
    port map (
            O => \N__10220\,
            I => \N__10212\
        );

    \I__2336\ : Span12Mux_v
    port map (
            O => \N__10217\,
            I => \N__10212\
        );

    \I__2335\ : Span12Mux_h
    port map (
            O => \N__10212\,
            I => \N__10209\
        );

    \I__2334\ : Odrv12
    port map (
            O => \N__10209\,
            I => \DRA_c_6\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10206\,
            I => \N__10203\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__10203\,
            I => \N__10199\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10202\,
            I => \N__10196\
        );

    \I__2330\ : Span4Mux_h
    port map (
            O => \N__10199\,
            I => \N__10189\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10196\,
            I => \N__10189\
        );

    \I__2328\ : InMux
    port map (
            O => \N__10195\,
            I => \N__10186\
        );

    \I__2327\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10183\
        );

    \I__2326\ : Span4Mux_v
    port map (
            O => \N__10189\,
            I => \N__10180\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__10186\,
            I => \N__10175\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__10183\,
            I => \N__10175\
        );

    \I__2323\ : Sp12to4
    port map (
            O => \N__10180\,
            I => \N__10170\
        );

    \I__2322\ : Span12Mux_v
    port map (
            O => \N__10175\,
            I => \N__10170\
        );

    \I__2321\ : Span12Mux_h
    port map (
            O => \N__10170\,
            I => \N__10167\
        );

    \I__2320\ : Odrv12
    port map (
            O => \N__10167\,
            I => \DRA_c_5\
        );

    \I__2319\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10161\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__10161\,
            I => \N__10158\
        );

    \I__2317\ : Span4Mux_v
    port map (
            O => \N__10158\,
            I => \N__10155\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__10155\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2315\ : InMux
    port map (
            O => \N__10152\,
            I => \N__10149\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__10149\,
            I => \N__10144\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10139\
        );

    \I__2312\ : InMux
    port map (
            O => \N__10147\,
            I => \N__10139\
        );

    \I__2311\ : Span4Mux_h
    port map (
            O => \N__10144\,
            I => \N__10134\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__10139\,
            I => \N__10134\
        );

    \I__2309\ : Span4Mux_h
    port map (
            O => \N__10134\,
            I => \N__10130\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10127\
        );

    \I__2307\ : Span4Mux_v
    port map (
            O => \N__10130\,
            I => \N__10124\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__10127\,
            I => \N__10121\
        );

    \I__2305\ : Sp12to4
    port map (
            O => \N__10124\,
            I => \N__10118\
        );

    \I__2304\ : Sp12to4
    port map (
            O => \N__10121\,
            I => \N__10115\
        );

    \I__2303\ : Span12Mux_h
    port map (
            O => \N__10118\,
            I => \N__10112\
        );

    \I__2302\ : Span12Mux_v
    port map (
            O => \N__10115\,
            I => \N__10109\
        );

    \I__2301\ : Span12Mux_v
    port map (
            O => \N__10112\,
            I => \N__10104\
        );

    \I__2300\ : Span12Mux_h
    port map (
            O => \N__10109\,
            I => \N__10104\
        );

    \I__2299\ : Odrv12
    port map (
            O => \N__10104\,
            I => \DRA_c_9\
        );

    \I__2298\ : InMux
    port map (
            O => \N__10101\,
            I => \N__10098\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__10098\,
            I => \N__10095\
        );

    \I__2296\ : Odrv12
    port map (
            O => \N__10095\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2295\ : InMux
    port map (
            O => \N__10092\,
            I => \N__10088\
        );

    \I__2294\ : InMux
    port map (
            O => \N__10091\,
            I => \N__10085\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__10088\,
            I => \N__10082\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__10085\,
            I => \N__10079\
        );

    \I__2291\ : Span4Mux_v
    port map (
            O => \N__10082\,
            I => \N__10073\
        );

    \I__2290\ : Span4Mux_h
    port map (
            O => \N__10079\,
            I => \N__10073\
        );

    \I__2289\ : InMux
    port map (
            O => \N__10078\,
            I => \N__10068\
        );

    \I__2288\ : Span4Mux_h
    port map (
            O => \N__10073\,
            I => \N__10065\
        );

    \I__2287\ : InMux
    port map (
            O => \N__10072\,
            I => \N__10062\
        );

    \I__2286\ : InMux
    port map (
            O => \N__10071\,
            I => \N__10059\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__10068\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__10065\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__10062\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__10059\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2281\ : IoInMux
    port map (
            O => \N__10050\,
            I => \N__10047\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__10047\,
            I => \N__10044\
        );

    \I__2279\ : Span4Mux_s3_v
    port map (
            O => \N__10044\,
            I => \N__10041\
        );

    \I__2278\ : Span4Mux_v
    port map (
            O => \N__10041\,
            I => \N__10038\
        );

    \I__2277\ : Span4Mux_h
    port map (
            O => \N__10038\,
            I => \N__10035\
        );

    \I__2276\ : Odrv4
    port map (
            O => \N__10035\,
            I => \CRCSn_c\
        );

    \I__2275\ : InMux
    port map (
            O => \N__10032\,
            I => \N__10029\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__10029\,
            I => \N__10024\
        );

    \I__2273\ : InMux
    port map (
            O => \N__10028\,
            I => \N__10021\
        );

    \I__2272\ : InMux
    port map (
            O => \N__10027\,
            I => \N__10018\
        );

    \I__2271\ : Span12Mux_h
    port map (
            O => \N__10024\,
            I => \N__10014\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__10021\,
            I => \N__10011\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__10018\,
            I => \N__10008\
        );

    \I__2268\ : InMux
    port map (
            O => \N__10017\,
            I => \N__10005\
        );

    \I__2267\ : Odrv12
    port map (
            O => \N__10014\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__10011\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2265\ : Odrv4
    port map (
            O => \N__10008\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__10005\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2263\ : IoInMux
    port map (
            O => \N__9996\,
            I => \N__9993\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__9993\,
            I => \N__9990\
        );

    \I__2261\ : Span12Mux_s5_h
    port map (
            O => \N__9990\,
            I => \N__9987\
        );

    \I__2260\ : Span12Mux_v
    port map (
            O => \N__9987\,
            I => \N__9984\
        );

    \I__2259\ : Odrv12
    port map (
            O => \N__9984\,
            I => \WEn_c\
        );

    \I__2258\ : InMux
    port map (
            O => \N__9981\,
            I => \N__9978\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__9978\,
            I => \N__9975\
        );

    \I__2256\ : Span4Mux_h
    port map (
            O => \N__9975\,
            I => \N__9972\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__9972\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2254\ : InMux
    port map (
            O => \N__9969\,
            I => \N__9966\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__9966\,
            I => \N__9963\
        );

    \I__2252\ : Odrv12
    port map (
            O => \N__9963\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2251\ : InMux
    port map (
            O => \N__9960\,
            I => \N__9957\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__9957\,
            I => \N__9954\
        );

    \I__2249\ : Span4Mux_h
    port map (
            O => \N__9954\,
            I => \N__9951\
        );

    \I__2248\ : Odrv4
    port map (
            O => \N__9951\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__9948\,
            I => \N__9945\
        );

    \I__2246\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9942\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__9942\,
            I => \N__9939\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__9939\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9936\,
            I => \N__9933\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__9933\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9930\,
            I => \N__9927\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__9927\,
            I => \N__9924\
        );

    \I__2239\ : Odrv4
    port map (
            O => \N__9924\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__9921\,
            I => \N__9917\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9920\,
            I => \N__9912\
        );

    \I__2236\ : InMux
    port map (
            O => \N__9917\,
            I => \N__9912\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__9912\,
            I => \U712_BYTE_ENABLE.N_298_i\
        );

    \I__2234\ : InMux
    port map (
            O => \N__9909\,
            I => \N__9906\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__9906\,
            I => \U712_REG_SM.N_459\
        );

    \I__2232\ : IoInMux
    port map (
            O => \N__9903\,
            I => \N__9900\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9900\,
            I => \N__9897\
        );

    \I__2230\ : Span4Mux_s2_v
    port map (
            O => \N__9897\,
            I => \N__9894\
        );

    \I__2229\ : Span4Mux_v
    port map (
            O => \N__9894\,
            I => \N__9891\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__9891\,
            I => \N_390_i\
        );

    \I__2227\ : IoInMux
    port map (
            O => \N__9888\,
            I => \N__9885\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__9885\,
            I => \N__9882\
        );

    \I__2225\ : Span4Mux_s2_v
    port map (
            O => \N__9882\,
            I => \N__9879\
        );

    \I__2224\ : Span4Mux_v
    port map (
            O => \N__9879\,
            I => \N__9876\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__9876\,
            I => \N_389_i\
        );

    \I__2222\ : InMux
    port map (
            O => \N__9873\,
            I => \N__9860\
        );

    \I__2221\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9860\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9871\,
            I => \N__9860\
        );

    \I__2219\ : InMux
    port map (
            O => \N__9870\,
            I => \N__9855\
        );

    \I__2218\ : InMux
    port map (
            O => \N__9869\,
            I => \N__9855\
        );

    \I__2217\ : InMux
    port map (
            O => \N__9868\,
            I => \N__9851\
        );

    \I__2216\ : InMux
    port map (
            O => \N__9867\,
            I => \N__9848\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__9860\,
            I => \N__9845\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__9855\,
            I => \N__9842\
        );

    \I__2213\ : InMux
    port map (
            O => \N__9854\,
            I => \N__9839\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__9851\,
            I => \N__9836\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__9848\,
            I => \N__9832\
        );

    \I__2210\ : Span4Mux_v
    port map (
            O => \N__9845\,
            I => \N__9827\
        );

    \I__2209\ : Span4Mux_v
    port map (
            O => \N__9842\,
            I => \N__9827\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__9839\,
            I => \N__9824\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__9836\,
            I => \N__9821\
        );

    \I__2206\ : InMux
    port map (
            O => \N__9835\,
            I => \N__9818\
        );

    \I__2205\ : Span12Mux_s10_v
    port map (
            O => \N__9832\,
            I => \N__9807\
        );

    \I__2204\ : Sp12to4
    port map (
            O => \N__9827\,
            I => \N__9807\
        );

    \I__2203\ : Span12Mux_h
    port map (
            O => \N__9824\,
            I => \N__9807\
        );

    \I__2202\ : Sp12to4
    port map (
            O => \N__9821\,
            I => \N__9807\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__9818\,
            I => \N__9807\
        );

    \I__2200\ : Span12Mux_h
    port map (
            O => \N__9807\,
            I => \N__9804\
        );

    \I__2199\ : Odrv12
    port map (
            O => \N__9804\,
            I => \A_c_0\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9801\,
            I => \N__9797\
        );

    \I__2197\ : InMux
    port map (
            O => \N__9800\,
            I => \N__9794\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__9797\,
            I => \N__9786\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__9794\,
            I => \N__9783\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9776\
        );

    \I__2193\ : InMux
    port map (
            O => \N__9792\,
            I => \N__9776\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9791\,
            I => \N__9776\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9790\,
            I => \N__9770\
        );

    \I__2190\ : InMux
    port map (
            O => \N__9789\,
            I => \N__9770\
        );

    \I__2189\ : Span4Mux_v
    port map (
            O => \N__9786\,
            I => \N__9767\
        );

    \I__2188\ : Span4Mux_v
    port map (
            O => \N__9783\,
            I => \N__9764\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__9776\,
            I => \N__9761\
        );

    \I__2186\ : InMux
    port map (
            O => \N__9775\,
            I => \N__9758\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__9770\,
            I => \N__9755\
        );

    \I__2184\ : Span4Mux_v
    port map (
            O => \N__9767\,
            I => \N__9752\
        );

    \I__2183\ : Span4Mux_v
    port map (
            O => \N__9764\,
            I => \N__9747\
        );

    \I__2182\ : Span4Mux_v
    port map (
            O => \N__9761\,
            I => \N__9747\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9758\,
            I => \N__9744\
        );

    \I__2180\ : Span12Mux_v
    port map (
            O => \N__9755\,
            I => \N__9735\
        );

    \I__2179\ : Sp12to4
    port map (
            O => \N__9752\,
            I => \N__9735\
        );

    \I__2178\ : Sp12to4
    port map (
            O => \N__9747\,
            I => \N__9735\
        );

    \I__2177\ : Span12Mux_s7_v
    port map (
            O => \N__9744\,
            I => \N__9735\
        );

    \I__2176\ : Span12Mux_h
    port map (
            O => \N__9735\,
            I => \N__9732\
        );

    \I__2175\ : Odrv12
    port map (
            O => \N__9732\,
            I => \A_c_1\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9729\,
            I => \N__9725\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9721\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9725\,
            I => \N__9717\
        );

    \I__2171\ : InMux
    port map (
            O => \N__9724\,
            I => \N__9714\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9721\,
            I => \N__9711\
        );

    \I__2169\ : InMux
    port map (
            O => \N__9720\,
            I => \N__9708\
        );

    \I__2168\ : Odrv4
    port map (
            O => \N__9717\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9714\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__9711\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9708\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9696\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__9696\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__9693\,
            I => \N__9690\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9690\,
            I => \N__9687\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__9687\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9684\,
            I => \N__9681\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__9681\,
            I => \N__9677\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9680\,
            I => \N__9674\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__9677\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9674\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9669\,
            I => \N__9660\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9660\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9660\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__9660\,
            I => \N__9657\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__9657\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9654\,
            I => \N__9651\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9651\,
            I => \N__9648\
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__9648\,
            I => \U712_REG_SM.N_402\
        );

    \I__2146\ : IoInMux
    port map (
            O => \N__9645\,
            I => \N__9642\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__9642\,
            I => \N__9639\
        );

    \I__2144\ : Span12Mux_s0_v
    port map (
            O => \N__9639\,
            I => \N__9635\
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__9638\,
            I => \N__9632\
        );

    \I__2142\ : Span12Mux_h
    port map (
            O => \N__9635\,
            I => \N__9629\
        );

    \I__2141\ : InMux
    port map (
            O => \N__9632\,
            I => \N__9626\
        );

    \I__2140\ : Odrv12
    port map (
            O => \N__9629\,
            I => \LDSn_c\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__9626\,
            I => \LDSn_c\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9614\
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__9620\,
            I => \N__9610\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__9619\,
            I => \N__9607\
        );

    \I__2135\ : CascadeMux
    port map (
            O => \N__9618\,
            I => \N__9602\
        );

    \I__2134\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9597\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__9614\,
            I => \N__9594\
        );

    \I__2132\ : InMux
    port map (
            O => \N__9613\,
            I => \N__9588\
        );

    \I__2131\ : InMux
    port map (
            O => \N__9610\,
            I => \N__9583\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9607\,
            I => \N__9583\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9606\,
            I => \N__9578\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9605\,
            I => \N__9578\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9574\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9601\,
            I => \N__9569\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9600\,
            I => \N__9569\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9597\,
            I => \N__9564\
        );

    \I__2123\ : Span4Mux_h
    port map (
            O => \N__9594\,
            I => \N__9564\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9557\
        );

    \I__2121\ : InMux
    port map (
            O => \N__9592\,
            I => \N__9557\
        );

    \I__2120\ : InMux
    port map (
            O => \N__9591\,
            I => \N__9557\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__9588\,
            I => \N__9550\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9583\,
            I => \N__9550\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9578\,
            I => \N__9550\
        );

    \I__2116\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9547\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9574\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__9569\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__9564\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__9557\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__9550\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9547\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__9534\,
            I => \N__9530\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9533\,
            I => \N__9524\
        );

    \I__2107\ : InMux
    port map (
            O => \N__9530\,
            I => \N__9524\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9529\,
            I => \N__9521\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__9524\,
            I => \N__9518\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9521\,
            I => \N__9515\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__9518\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\
        );

    \I__2102\ : Odrv4
    port map (
            O => \N__9515\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\
        );

    \I__2101\ : IoInMux
    port map (
            O => \N__9510\,
            I => \N__9507\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__9507\,
            I => \N__9504\
        );

    \I__2099\ : Span4Mux_s2_v
    port map (
            O => \N__9504\,
            I => \N__9501\
        );

    \I__2098\ : Span4Mux_v
    port map (
            O => \N__9501\,
            I => \N__9498\
        );

    \I__2097\ : Span4Mux_v
    port map (
            O => \N__9498\,
            I => \N__9495\
        );

    \I__2096\ : Sp12to4
    port map (
            O => \N__9495\,
            I => \N__9491\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9488\
        );

    \I__2094\ : Odrv12
    port map (
            O => \N__9491\,
            I => \UDSn_c\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__9488\,
            I => \UDSn_c\
        );

    \I__2092\ : IoInMux
    port map (
            O => \N__9483\,
            I => \N__9480\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__9480\,
            I => \N__9477\
        );

    \I__2090\ : Span4Mux_s0_v
    port map (
            O => \N__9477\,
            I => \N__9474\
        );

    \I__2089\ : Span4Mux_v
    port map (
            O => \N__9474\,
            I => \N__9471\
        );

    \I__2088\ : Odrv4
    port map (
            O => \N__9471\,
            I => \RESETn_c_i\
        );

    \I__2087\ : IoInMux
    port map (
            O => \N__9468\,
            I => \N__9465\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9465\,
            I => \N__9462\
        );

    \I__2085\ : Span12Mux_s6_v
    port map (
            O => \N__9462\,
            I => \N__9459\
        );

    \I__2084\ : Odrv12
    port map (
            O => \N__9459\,
            I => \N_166\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9456\,
            I => \N__9443\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9455\,
            I => \N__9425\
        );

    \I__2081\ : InMux
    port map (
            O => \N__9454\,
            I => \N__9425\
        );

    \I__2080\ : InMux
    port map (
            O => \N__9453\,
            I => \N__9425\
        );

    \I__2079\ : InMux
    port map (
            O => \N__9452\,
            I => \N__9425\
        );

    \I__2078\ : InMux
    port map (
            O => \N__9451\,
            I => \N__9425\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9450\,
            I => \N__9425\
        );

    \I__2076\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9420\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9448\,
            I => \N__9420\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__9447\,
            I => \N__9414\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__9446\,
            I => \N__9411\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__9443\,
            I => \N__9403\
        );

    \I__2071\ : InMux
    port map (
            O => \N__9442\,
            I => \N__9400\
        );

    \I__2070\ : InMux
    port map (
            O => \N__9441\,
            I => \N__9391\
        );

    \I__2069\ : InMux
    port map (
            O => \N__9440\,
            I => \N__9391\
        );

    \I__2068\ : InMux
    port map (
            O => \N__9439\,
            I => \N__9391\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9438\,
            I => \N__9391\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__9425\,
            I => \N__9386\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9420\,
            I => \N__9386\
        );

    \I__2064\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9381\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9381\
        );

    \I__2062\ : InMux
    port map (
            O => \N__9417\,
            I => \N__9378\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9375\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9411\,
            I => \N__9372\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__9410\,
            I => \N__9369\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__9409\,
            I => \N__9366\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__9408\,
            I => \N__9363\
        );

    \I__2056\ : CascadeMux
    port map (
            O => \N__9407\,
            I => \N__9360\
        );

    \I__2055\ : InMux
    port map (
            O => \N__9406\,
            I => \N__9357\
        );

    \I__2054\ : Span4Mux_v
    port map (
            O => \N__9403\,
            I => \N__9345\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9400\,
            I => \N__9345\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__9391\,
            I => \N__9345\
        );

    \I__2051\ : Span4Mux_v
    port map (
            O => \N__9386\,
            I => \N__9345\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__9381\,
            I => \N__9345\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9378\,
            I => \N__9339\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9375\,
            I => \N__9339\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9372\,
            I => \N__9336\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9369\,
            I => \N__9333\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9366\,
            I => \N__9330\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9327\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9360\,
            I => \N__9324\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9357\,
            I => \N__9321\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9356\,
            I => \N__9318\
        );

    \I__2040\ : Span4Mux_h
    port map (
            O => \N__9345\,
            I => \N__9315\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9344\,
            I => \N__9312\
        );

    \I__2038\ : Span4Mux_h
    port map (
            O => \N__9339\,
            I => \N__9303\
        );

    \I__2037\ : Span4Mux_h
    port map (
            O => \N__9336\,
            I => \N__9303\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9333\,
            I => \N__9303\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__9330\,
            I => \N__9303\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__9327\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9324\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2032\ : Odrv12
    port map (
            O => \N__9321\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9318\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__9315\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__9312\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__9303\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2027\ : IoInMux
    port map (
            O => \N__9288\,
            I => \N__9285\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__9285\,
            I => \N__9282\
        );

    \I__2025\ : Span4Mux_s2_v
    port map (
            O => \N__9282\,
            I => \N__9279\
        );

    \I__2024\ : Span4Mux_h
    port map (
            O => \N__9279\,
            I => \N__9276\
        );

    \I__2023\ : Sp12to4
    port map (
            O => \N__9276\,
            I => \N__9273\
        );

    \I__2022\ : Span12Mux_s11_v
    port map (
            O => \N__9273\,
            I => \N__9270\
        );

    \I__2021\ : Odrv12
    port map (
            O => \N__9270\,
            I => \CASn_c\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9267\,
            I => \N__9264\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__9264\,
            I => \N__9261\
        );

    \I__2018\ : Span4Mux_v
    port map (
            O => \N__9261\,
            I => \N__9258\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__9258\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9255\,
            I => \N__9252\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9252\,
            I => \N__9249\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__9249\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2013\ : InMux
    port map (
            O => \N__9246\,
            I => \N__9243\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__9243\,
            I => \N__9240\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__9240\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2010\ : InMux
    port map (
            O => \N__9237\,
            I => \N__9229\
        );

    \I__2009\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9229\
        );

    \I__2008\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9223\
        );

    \I__2007\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9223\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__9229\,
            I => \N__9220\
        );

    \I__2005\ : InMux
    port map (
            O => \N__9228\,
            I => \N__9217\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__9223\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__9220\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9217\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__9210\,
            I => \N__9206\
        );

    \I__2000\ : InMux
    port map (
            O => \N__9209\,
            I => \N__9201\
        );

    \I__1999\ : InMux
    port map (
            O => \N__9206\,
            I => \N__9201\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__9201\,
            I => \N__9189\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9200\,
            I => \N__9182\
        );

    \I__1996\ : InMux
    port map (
            O => \N__9199\,
            I => \N__9182\
        );

    \I__1995\ : InMux
    port map (
            O => \N__9198\,
            I => \N__9182\
        );

    \I__1994\ : InMux
    port map (
            O => \N__9197\,
            I => \N__9174\
        );

    \I__1993\ : InMux
    port map (
            O => \N__9196\,
            I => \N__9174\
        );

    \I__1992\ : InMux
    port map (
            O => \N__9195\,
            I => \N__9174\
        );

    \I__1991\ : InMux
    port map (
            O => \N__9194\,
            I => \N__9167\
        );

    \I__1990\ : InMux
    port map (
            O => \N__9193\,
            I => \N__9167\
        );

    \I__1989\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9167\
        );

    \I__1988\ : Span4Mux_v
    port map (
            O => \N__9189\,
            I => \N__9164\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__9182\,
            I => \N__9161\
        );

    \I__1986\ : InMux
    port map (
            O => \N__9181\,
            I => \N__9158\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__9174\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__9167\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__9164\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__9161\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__9158\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__9147\,
            I => \N__9140\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__9146\,
            I => \N__9136\
        );

    \I__1978\ : InMux
    port map (
            O => \N__9145\,
            I => \N__9133\
        );

    \I__1977\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9130\
        );

    \I__1976\ : InMux
    port map (
            O => \N__9143\,
            I => \N__9127\
        );

    \I__1975\ : InMux
    port map (
            O => \N__9140\,
            I => \N__9122\
        );

    \I__1974\ : InMux
    port map (
            O => \N__9139\,
            I => \N__9122\
        );

    \I__1973\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9119\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__9133\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__9130\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__9127\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__9122\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__9119\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1967\ : CascadeMux
    port map (
            O => \N__9108\,
            I => \U712_CYCLE_TERM.N_452_cascade_\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__9105\,
            I => \N__9102\
        );

    \I__1965\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9098\
        );

    \I__1964\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9093\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__9098\,
            I => \N__9090\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9087\
        );

    \I__1961\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9084\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__9093\,
            I => \N__9081\
        );

    \I__1959\ : Span4Mux_v
    port map (
            O => \N__9090\,
            I => \N__9078\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__9087\,
            I => \N__9071\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__9084\,
            I => \N__9071\
        );

    \I__1956\ : Span4Mux_h
    port map (
            O => \N__9081\,
            I => \N__9071\
        );

    \I__1955\ : Sp12to4
    port map (
            O => \N__9078\,
            I => \N__9068\
        );

    \I__1954\ : Sp12to4
    port map (
            O => \N__9071\,
            I => \N__9063\
        );

    \I__1953\ : Span12Mux_h
    port map (
            O => \N__9068\,
            I => \N__9063\
        );

    \I__1952\ : Span12Mux_v
    port map (
            O => \N__9063\,
            I => \N__9060\
        );

    \I__1951\ : Odrv12
    port map (
            O => \N__9060\,
            I => \CLK40_PLL_i\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__9057\,
            I => \N__9052\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__9056\,
            I => \N__9048\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__9055\,
            I => \N__9040\
        );

    \I__1947\ : InMux
    port map (
            O => \N__9052\,
            I => \N__9029\
        );

    \I__1946\ : InMux
    port map (
            O => \N__9051\,
            I => \N__9029\
        );

    \I__1945\ : InMux
    port map (
            O => \N__9048\,
            I => \N__9026\
        );

    \I__1944\ : InMux
    port map (
            O => \N__9047\,
            I => \N__9018\
        );

    \I__1943\ : InMux
    port map (
            O => \N__9046\,
            I => \N__9018\
        );

    \I__1942\ : InMux
    port map (
            O => \N__9045\,
            I => \N__9018\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9044\,
            I => \N__9013\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9043\,
            I => \N__9013\
        );

    \I__1939\ : InMux
    port map (
            O => \N__9040\,
            I => \N__9008\
        );

    \I__1938\ : InMux
    port map (
            O => \N__9039\,
            I => \N__9005\
        );

    \I__1937\ : InMux
    port map (
            O => \N__9038\,
            I => \N__8996\
        );

    \I__1936\ : InMux
    port map (
            O => \N__9037\,
            I => \N__8996\
        );

    \I__1935\ : InMux
    port map (
            O => \N__9036\,
            I => \N__8996\
        );

    \I__1934\ : InMux
    port map (
            O => \N__9035\,
            I => \N__8991\
        );

    \I__1933\ : InMux
    port map (
            O => \N__9034\,
            I => \N__8991\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__9029\,
            I => \N__8987\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__9026\,
            I => \N__8984\
        );

    \I__1930\ : InMux
    port map (
            O => \N__9025\,
            I => \N__8981\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__9018\,
            I => \N__8978\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__9013\,
            I => \N__8975\
        );

    \I__1927\ : InMux
    port map (
            O => \N__9012\,
            I => \N__8970\
        );

    \I__1926\ : InMux
    port map (
            O => \N__9011\,
            I => \N__8970\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__9008\,
            I => \N__8967\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__9005\,
            I => \N__8964\
        );

    \I__1923\ : InMux
    port map (
            O => \N__9004\,
            I => \N__8959\
        );

    \I__1922\ : InMux
    port map (
            O => \N__9003\,
            I => \N__8959\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__8996\,
            I => \N__8954\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__8991\,
            I => \N__8954\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8951\
        );

    \I__1918\ : Span4Mux_v
    port map (
            O => \N__8987\,
            I => \N__8948\
        );

    \I__1917\ : Span4Mux_h
    port map (
            O => \N__8984\,
            I => \N__8945\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__8981\,
            I => \N__8940\
        );

    \I__1915\ : Span4Mux_h
    port map (
            O => \N__8978\,
            I => \N__8940\
        );

    \I__1914\ : Span4Mux_h
    port map (
            O => \N__8975\,
            I => \N__8937\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__8970\,
            I => \N__8931\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__8967\,
            I => \N__8922\
        );

    \I__1911\ : Span4Mux_h
    port map (
            O => \N__8964\,
            I => \N__8922\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__8959\,
            I => \N__8922\
        );

    \I__1909\ : Span4Mux_v
    port map (
            O => \N__8954\,
            I => \N__8922\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8951\,
            I => \N__8919\
        );

    \I__1907\ : Span4Mux_h
    port map (
            O => \N__8948\,
            I => \N__8914\
        );

    \I__1906\ : Span4Mux_v
    port map (
            O => \N__8945\,
            I => \N__8914\
        );

    \I__1905\ : Span4Mux_h
    port map (
            O => \N__8940\,
            I => \N__8911\
        );

    \I__1904\ : Span4Mux_h
    port map (
            O => \N__8937\,
            I => \N__8908\
        );

    \I__1903\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8901\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8935\,
            I => \N__8901\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8934\,
            I => \N__8901\
        );

    \I__1900\ : Span4Mux_h
    port map (
            O => \N__8931\,
            I => \N__8896\
        );

    \I__1899\ : Span4Mux_h
    port map (
            O => \N__8922\,
            I => \N__8896\
        );

    \I__1898\ : Odrv12
    port map (
            O => \N__8919\,
            I => \CPU_CYCLEm\
        );

    \I__1897\ : Odrv4
    port map (
            O => \N__8914\,
            I => \CPU_CYCLEm\
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__8911\,
            I => \CPU_CYCLEm\
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__8908\,
            I => \CPU_CYCLEm\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__8901\,
            I => \CPU_CYCLEm\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__8896\,
            I => \CPU_CYCLEm\
        );

    \I__1892\ : CascadeMux
    port map (
            O => \N__8883\,
            I => \U712_BYTE_ENABLE.N_421_cascade_\
        );

    \I__1891\ : IoInMux
    port map (
            O => \N__8880\,
            I => \N__8877\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__8877\,
            I => \N__8874\
        );

    \I__1889\ : Span4Mux_s3_h
    port map (
            O => \N__8874\,
            I => \N__8871\
        );

    \I__1888\ : Span4Mux_v
    port map (
            O => \N__8871\,
            I => \N__8868\
        );

    \I__1887\ : Sp12to4
    port map (
            O => \N__8868\,
            I => \N__8865\
        );

    \I__1886\ : Span12Mux_h
    port map (
            O => \N__8865\,
            I => \N__8862\
        );

    \I__1885\ : Odrv12
    port map (
            O => \N__8862\,
            I => \N_168_i\
        );

    \I__1884\ : InMux
    port map (
            O => \N__8859\,
            I => \N__8856\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__8856\,
            I => \U712_CYCLE_TERM.N_326\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__8853\,
            I => \N__8850\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8844\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8841\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8848\,
            I => \N__8838\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__8847\,
            I => \N__8835\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8844\,
            I => \N__8830\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8841\,
            I => \N__8830\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8838\,
            I => \N__8827\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8835\,
            I => \N__8824\
        );

    \I__1873\ : Span4Mux_h
    port map (
            O => \N__8830\,
            I => \N__8819\
        );

    \I__1872\ : Span4Mux_v
    port map (
            O => \N__8827\,
            I => \N__8819\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8824\,
            I => \REG_TACK\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__8819\,
            I => \REG_TACK\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8814\,
            I => \N__8807\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8807\
        );

    \I__1867\ : InMux
    port map (
            O => \N__8812\,
            I => \N__8804\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__8807\,
            I => \N__8798\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8804\,
            I => \N__8798\
        );

    \I__1864\ : InMux
    port map (
            O => \N__8803\,
            I => \N__8795\
        );

    \I__1863\ : Span12Mux_v
    port map (
            O => \N__8798\,
            I => \N__8792\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8795\,
            I => \CPU_TACKm\
        );

    \I__1861\ : Odrv12
    port map (
            O => \N__8792\,
            I => \CPU_TACKm\
        );

    \I__1860\ : IoInMux
    port map (
            O => \N__8787\,
            I => \N__8784\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__8784\,
            I => \N__8781\
        );

    \I__1858\ : Span4Mux_s1_v
    port map (
            O => \N__8781\,
            I => \N__8775\
        );

    \I__1857\ : InMux
    port map (
            O => \N__8780\,
            I => \N__8772\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8779\,
            I => \N__8767\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8778\,
            I => \N__8767\
        );

    \I__1854\ : Sp12to4
    port map (
            O => \N__8775\,
            I => \N__8763\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8772\,
            I => \N__8758\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__8767\,
            I => \N__8758\
        );

    \I__1851\ : InMux
    port map (
            O => \N__8766\,
            I => \N__8755\
        );

    \I__1850\ : Span12Mux_h
    port map (
            O => \N__8763\,
            I => \N__8752\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__8758\,
            I => \N__8749\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8755\,
            I => \N__8746\
        );

    \I__1847\ : Span12Mux_v
    port map (
            O => \N__8752\,
            I => \N__8742\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__8749\,
            I => \N__8739\
        );

    \I__1845\ : Span4Mux_v
    port map (
            O => \N__8746\,
            I => \N__8736\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8745\,
            I => \N__8733\
        );

    \I__1843\ : Odrv12
    port map (
            O => \N__8742\,
            I => \DBENn_c\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__8739\,
            I => \DBENn_c\
        );

    \I__1841\ : Odrv4
    port map (
            O => \N__8736\,
            I => \DBENn_c\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8733\,
            I => \DBENn_c\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8724\,
            I => \N__8717\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8723\,
            I => \N__8714\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8722\,
            I => \N__8709\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8721\,
            I => \N__8709\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8705\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__8717\,
            I => \N__8702\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__8714\,
            I => \N__8697\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8709\,
            I => \N__8697\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8694\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8705\,
            I => \N__8691\
        );

    \I__1829\ : Span4Mux_v
    port map (
            O => \N__8702\,
            I => \N__8686\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__8697\,
            I => \N__8686\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8694\,
            I => \N__8683\
        );

    \I__1826\ : Span4Mux_h
    port map (
            O => \N__8691\,
            I => \N__8680\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__8686\,
            I => \DMA_CYCLEm\
        );

    \I__1824\ : Odrv12
    port map (
            O => \N__8683\,
            I => \DMA_CYCLEm\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__8680\,
            I => \DMA_CYCLEm\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__8673\,
            I => \N__8670\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8670\,
            I => \N__8667\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8667\,
            I => \U712_BYTE_ENABLE.N_425\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__8664\,
            I => \N__8660\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8656\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8660\,
            I => \N__8653\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8659\,
            I => \N__8650\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__8656\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8653\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8650\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8643\,
            I => \N__8640\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8640\,
            I => \N__8637\
        );

    \I__1810\ : Span4Mux_h
    port map (
            O => \N__8637\,
            I => \N__8634\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__8634\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8631\,
            I => \N__8628\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8628\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8622\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__8622\,
            I => \N__8619\
        );

    \I__1804\ : Odrv12
    port map (
            O => \N__8619\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\
        );

    \I__1803\ : IoInMux
    port map (
            O => \N__8616\,
            I => \N__8611\
        );

    \I__1802\ : IoInMux
    port map (
            O => \N__8615\,
            I => \N__8608\
        );

    \I__1801\ : IoInMux
    port map (
            O => \N__8614\,
            I => \N__8605\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__8611\,
            I => \N__8602\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8608\,
            I => \N__8599\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8605\,
            I => \N__8596\
        );

    \I__1797\ : Span4Mux_s2_v
    port map (
            O => \N__8602\,
            I => \N__8593\
        );

    \I__1796\ : Span4Mux_s2_v
    port map (
            O => \N__8599\,
            I => \N__8590\
        );

    \I__1795\ : Span4Mux_s3_h
    port map (
            O => \N__8596\,
            I => \N__8587\
        );

    \I__1794\ : Sp12to4
    port map (
            O => \N__8593\,
            I => \N__8582\
        );

    \I__1793\ : Sp12to4
    port map (
            O => \N__8590\,
            I => \N__8582\
        );

    \I__1792\ : Sp12to4
    port map (
            O => \N__8587\,
            I => \N__8579\
        );

    \I__1791\ : Span12Mux_h
    port map (
            O => \N__8582\,
            I => \N__8576\
        );

    \I__1790\ : Span12Mux_v
    port map (
            O => \N__8579\,
            I => \N__8573\
        );

    \I__1789\ : Span12Mux_v
    port map (
            O => \N__8576\,
            I => \N__8570\
        );

    \I__1788\ : Span12Mux_h
    port map (
            O => \N__8573\,
            I => \N__8567\
        );

    \I__1787\ : Odrv12
    port map (
            O => \N__8570\,
            I => \CLK40_PLL_i_i\
        );

    \I__1786\ : Odrv12
    port map (
            O => \N__8567\,
            I => \CLK40_PLL_i_i\
        );

    \I__1785\ : IoInMux
    port map (
            O => \N__8562\,
            I => \N__8557\
        );

    \I__1784\ : IoInMux
    port map (
            O => \N__8561\,
            I => \N__8554\
        );

    \I__1783\ : IoInMux
    port map (
            O => \N__8560\,
            I => \N__8551\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8557\,
            I => \N__8548\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__8554\,
            I => \N__8545\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8551\,
            I => \N__8542\
        );

    \I__1779\ : IoSpan4Mux
    port map (
            O => \N__8548\,
            I => \N__8539\
        );

    \I__1778\ : Span4Mux_s3_v
    port map (
            O => \N__8545\,
            I => \N__8536\
        );

    \I__1777\ : Span4Mux_s3_h
    port map (
            O => \N__8542\,
            I => \N__8533\
        );

    \I__1776\ : Sp12to4
    port map (
            O => \N__8539\,
            I => \N__8530\
        );

    \I__1775\ : Sp12to4
    port map (
            O => \N__8536\,
            I => \N__8527\
        );

    \I__1774\ : Sp12to4
    port map (
            O => \N__8533\,
            I => \N__8524\
        );

    \I__1773\ : Span12Mux_s7_v
    port map (
            O => \N__8530\,
            I => \N__8521\
        );

    \I__1772\ : Span12Mux_h
    port map (
            O => \N__8527\,
            I => \N__8518\
        );

    \I__1771\ : Span12Mux_v
    port map (
            O => \N__8524\,
            I => \N__8515\
        );

    \I__1770\ : Span12Mux_h
    port map (
            O => \N__8521\,
            I => \N__8511\
        );

    \I__1769\ : Span12Mux_v
    port map (
            O => \N__8518\,
            I => \N__8506\
        );

    \I__1768\ : Span12Mux_h
    port map (
            O => \N__8515\,
            I => \N__8506\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8514\,
            I => \N__8503\
        );

    \I__1766\ : Odrv12
    port map (
            O => \N__8511\,
            I => \TACK_EN\
        );

    \I__1765\ : Odrv12
    port map (
            O => \N__8506\,
            I => \TACK_EN\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8503\,
            I => \TACK_EN\
        );

    \I__1763\ : IoInMux
    port map (
            O => \N__8496\,
            I => \N__8493\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__8493\,
            I => \N__8490\
        );

    \I__1761\ : IoSpan4Mux
    port map (
            O => \N__8490\,
            I => \N__8487\
        );

    \I__1760\ : IoSpan4Mux
    port map (
            O => \N__8487\,
            I => \N__8484\
        );

    \I__1759\ : Span4Mux_s3_h
    port map (
            O => \N__8484\,
            I => \N__8481\
        );

    \I__1758\ : Span4Mux_v
    port map (
            O => \N__8481\,
            I => \N__8478\
        );

    \I__1757\ : Span4Mux_v
    port map (
            O => \N__8478\,
            I => \N__8474\
        );

    \I__1756\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8471\
        );

    \I__1755\ : Sp12to4
    port map (
            O => \N__8474\,
            I => \N__8468\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8471\,
            I => \N__8465\
        );

    \I__1753\ : Span12Mux_h
    port map (
            O => \N__8468\,
            I => \N__8460\
        );

    \I__1752\ : Span12Mux_v
    port map (
            O => \N__8465\,
            I => \N__8460\
        );

    \I__1751\ : Span12Mux_h
    port map (
            O => \N__8460\,
            I => \N__8457\
        );

    \I__1750\ : Odrv12
    port map (
            O => \N__8457\,
            I => \C3_c\
        );

    \I__1749\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8451\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8451\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8448\,
            I => \N__8443\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8447\,
            I => \N__8440\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8446\,
            I => \N__8437\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__8443\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8440\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__8437\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8426\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8423\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8426\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8423\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__8418\,
            I => \U712_BYTE_ENABLE.N_443_cascade_\
        );

    \I__1736\ : IoInMux
    port map (
            O => \N__8415\,
            I => \N__8412\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8412\,
            I => \N__8409\
        );

    \I__1734\ : IoSpan4Mux
    port map (
            O => \N__8409\,
            I => \N__8406\
        );

    \I__1733\ : Span4Mux_s2_h
    port map (
            O => \N__8406\,
            I => \N__8403\
        );

    \I__1732\ : Sp12to4
    port map (
            O => \N__8403\,
            I => \N__8400\
        );

    \I__1731\ : Span12Mux_h
    port map (
            O => \N__8400\,
            I => \N__8397\
        );

    \I__1730\ : Span12Mux_v
    port map (
            O => \N__8397\,
            I => \N__8394\
        );

    \I__1729\ : Odrv12
    port map (
            O => \N__8394\,
            I => \N_54_i\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8391\,
            I => \N__8385\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8382\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8379\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__8388\,
            I => \N__8370\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8385\,
            I => \N__8365\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8382\,
            I => \N__8365\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__8379\,
            I => \N__8362\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8378\,
            I => \N__8359\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8356\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8351\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8375\,
            I => \N__8351\
        );

    \I__1717\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8346\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8373\,
            I => \N__8346\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8343\
        );

    \I__1714\ : Span4Mux_v
    port map (
            O => \N__8365\,
            I => \N__8340\
        );

    \I__1713\ : Span4Mux_h
    port map (
            O => \N__8362\,
            I => \N__8337\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__8359\,
            I => \U712_CHIP_RAM.N_309\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8356\,
            I => \U712_CHIP_RAM.N_309\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__8351\,
            I => \U712_CHIP_RAM.N_309\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__8346\,
            I => \U712_CHIP_RAM.N_309\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__8343\,
            I => \U712_CHIP_RAM.N_309\
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__8340\,
            I => \U712_CHIP_RAM.N_309\
        );

    \I__1706\ : Odrv4
    port map (
            O => \N__8337\,
            I => \U712_CHIP_RAM.N_309\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8322\,
            I => \N__8319\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__8319\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__8316\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1_cascade_\
        );

    \I__1702\ : IoInMux
    port map (
            O => \N__8313\,
            I => \N__8310\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8310\,
            I => \N__8307\
        );

    \I__1700\ : Span12Mux_s9_v
    port map (
            O => \N__8307\,
            I => \N__8304\
        );

    \I__1699\ : Odrv12
    port map (
            O => \N__8304\,
            I => \CMA_c_1\
        );

    \I__1698\ : CEMux
    port map (
            O => \N__8301\,
            I => \N__8297\
        );

    \I__1697\ : CEMux
    port map (
            O => \N__8300\,
            I => \N__8294\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__8297\,
            I => \N__8287\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8294\,
            I => \N__8284\
        );

    \I__1694\ : CEMux
    port map (
            O => \N__8293\,
            I => \N__8281\
        );

    \I__1693\ : CEMux
    port map (
            O => \N__8292\,
            I => \N__8278\
        );

    \I__1692\ : CEMux
    port map (
            O => \N__8291\,
            I => \N__8275\
        );

    \I__1691\ : CEMux
    port map (
            O => \N__8290\,
            I => \N__8272\
        );

    \I__1690\ : Span4Mux_v
    port map (
            O => \N__8287\,
            I => \N__8265\
        );

    \I__1689\ : Span4Mux_h
    port map (
            O => \N__8284\,
            I => \N__8265\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8281\,
            I => \N__8265\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__8278\,
            I => \N__8260\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8275\,
            I => \N__8260\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8272\,
            I => \N__8257\
        );

    \I__1684\ : Span4Mux_h
    port map (
            O => \N__8265\,
            I => \N__8254\
        );

    \I__1683\ : Span4Mux_v
    port map (
            O => \N__8260\,
            I => \N__8251\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__8257\,
            I => \N__8248\
        );

    \I__1681\ : Odrv4
    port map (
            O => \N__8254\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__8251\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__8248\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__1678\ : InMux
    port map (
            O => \N__8241\,
            I => \N__8238\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__8238\,
            I => \N__8235\
        );

    \I__1676\ : Span12Mux_v
    port map (
            O => \N__8235\,
            I => \N__8232\
        );

    \I__1675\ : Span12Mux_h
    port map (
            O => \N__8232\,
            I => \N__8229\
        );

    \I__1674\ : Odrv12
    port map (
            O => \N__8229\,
            I => \A_c_15\
        );

    \I__1673\ : InMux
    port map (
            O => \N__8226\,
            I => \N__8222\
        );

    \I__1672\ : InMux
    port map (
            O => \N__8225\,
            I => \N__8219\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__8222\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8219\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__8214\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\
        );

    \I__1668\ : InMux
    port map (
            O => \N__8211\,
            I => \N__8208\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__8208\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1666\ : IoInMux
    port map (
            O => \N__8205\,
            I => \N__8202\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__8202\,
            I => \N__8199\
        );

    \I__1664\ : IoSpan4Mux
    port map (
            O => \N__8199\,
            I => \N__8196\
        );

    \I__1663\ : IoSpan4Mux
    port map (
            O => \N__8196\,
            I => \N__8192\
        );

    \I__1662\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8189\
        );

    \I__1661\ : Span4Mux_s2_v
    port map (
            O => \N__8192\,
            I => \N__8186\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__8189\,
            I => \N__8183\
        );

    \I__1659\ : Sp12to4
    port map (
            O => \N__8186\,
            I => \N__8180\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__8183\,
            I => \N__8177\
        );

    \I__1657\ : Span12Mux_s8_v
    port map (
            O => \N__8180\,
            I => \N__8174\
        );

    \I__1656\ : Sp12to4
    port map (
            O => \N__8177\,
            I => \N__8171\
        );

    \I__1655\ : Span12Mux_v
    port map (
            O => \N__8174\,
            I => \N__8166\
        );

    \I__1654\ : Span12Mux_h
    port map (
            O => \N__8171\,
            I => \N__8166\
        );

    \I__1653\ : Odrv12
    port map (
            O => \N__8166\,
            I => \A_c_10\
        );

    \I__1652\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8159\
        );

    \I__1651\ : InMux
    port map (
            O => \N__8162\,
            I => \N__8156\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__8159\,
            I => \N__8153\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__8156\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__8153\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__8148\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\
        );

    \I__1646\ : InMux
    port map (
            O => \N__8145\,
            I => \N__8142\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__8142\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__1644\ : InMux
    port map (
            O => \N__8139\,
            I => \N__8136\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__8136\,
            I => \N__8133\
        );

    \I__1642\ : Span12Mux_v
    port map (
            O => \N__8133\,
            I => \N__8130\
        );

    \I__1641\ : Span12Mux_h
    port map (
            O => \N__8130\,
            I => \N__8127\
        );

    \I__1640\ : Odrv12
    port map (
            O => \N__8127\,
            I => \A_c_13\
        );

    \I__1639\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8120\
        );

    \I__1638\ : InMux
    port map (
            O => \N__8123\,
            I => \N__8117\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__8120\,
            I => \N__8114\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__8117\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\
        );

    \I__1635\ : Odrv4
    port map (
            O => \N__8114\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__8109\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\
        );

    \I__1633\ : InMux
    port map (
            O => \N__8106\,
            I => \N__8103\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__8103\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1631\ : InMux
    port map (
            O => \N__8100\,
            I => \N__8094\
        );

    \I__1630\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8094\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__8094\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__1628\ : IoInMux
    port map (
            O => \N__8091\,
            I => \N__8088\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__8088\,
            I => \N__8085\
        );

    \I__1626\ : IoSpan4Mux
    port map (
            O => \N__8085\,
            I => \N__8082\
        );

    \I__1625\ : IoSpan4Mux
    port map (
            O => \N__8082\,
            I => \N__8079\
        );

    \I__1624\ : Span4Mux_s1_v
    port map (
            O => \N__8079\,
            I => \N__8076\
        );

    \I__1623\ : Sp12to4
    port map (
            O => \N__8076\,
            I => \N__8073\
        );

    \I__1622\ : Span12Mux_s9_v
    port map (
            O => \N__8073\,
            I => \N__8070\
        );

    \I__1621\ : Odrv12
    port map (
            O => \N__8070\,
            I => \ASn_c\
        );

    \I__1620\ : CEMux
    port map (
            O => \N__8067\,
            I => \N__8064\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__8064\,
            I => \N__8061\
        );

    \I__1618\ : Span4Mux_h
    port map (
            O => \N__8061\,
            I => \N__8058\
        );

    \I__1617\ : Odrv4
    port map (
            O => \N__8058\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0\
        );

    \I__1616\ : IoInMux
    port map (
            O => \N__8055\,
            I => \N__8052\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__8052\,
            I => \N__8049\
        );

    \I__1614\ : Span4Mux_s3_v
    port map (
            O => \N__8049\,
            I => \N__8046\
        );

    \I__1613\ : Span4Mux_h
    port map (
            O => \N__8046\,
            I => \N__8043\
        );

    \I__1612\ : Span4Mux_h
    port map (
            O => \N__8043\,
            I => \N__8040\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__8040\,
            I => \RASn_c\
        );

    \I__1610\ : InMux
    port map (
            O => \N__8037\,
            I => \N__8034\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__8034\,
            I => \N__8031\
        );

    \I__1608\ : Odrv12
    port map (
            O => \N__8031\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1607\ : InMux
    port map (
            O => \N__8028\,
            I => \N__8025\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__8025\,
            I => \N__8022\
        );

    \I__1605\ : Odrv12
    port map (
            O => \N__8022\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__1604\ : InMux
    port map (
            O => \N__8019\,
            I => \N__8016\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__8016\,
            I => \N__8013\
        );

    \I__1602\ : Span4Mux_h
    port map (
            O => \N__8013\,
            I => \N__8007\
        );

    \I__1601\ : InMux
    port map (
            O => \N__8012\,
            I => \N__8004\
        );

    \I__1600\ : InMux
    port map (
            O => \N__8011\,
            I => \N__8001\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8010\,
            I => \N__7998\
        );

    \I__1598\ : Span4Mux_v
    port map (
            O => \N__8007\,
            I => \N__7991\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__8004\,
            I => \N__7991\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__8001\,
            I => \N__7986\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7998\,
            I => \N__7986\
        );

    \I__1594\ : InMux
    port map (
            O => \N__7997\,
            I => \N__7983\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7996\,
            I => \N__7980\
        );

    \I__1592\ : Odrv4
    port map (
            O => \N__7991\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1591\ : Odrv12
    port map (
            O => \N__7986\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__7983\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7980\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__7971\,
            I => \U712_CHIP_RAM.N_309_cascade_\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__7968\,
            I => \U712_REG_SM.N_325_cascade_\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7962\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7962\,
            I => \U712_REG_SM.N_302\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__7959\,
            I => \U712_REG_SM.N_302_cascade_\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7956\,
            I => \N__7953\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7953\,
            I => \N__7950\
        );

    \I__1581\ : Span4Mux_v
    port map (
            O => \N__7950\,
            I => \N__7945\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7949\,
            I => \N__7942\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7948\,
            I => \N__7939\
        );

    \I__1578\ : Odrv4
    port map (
            O => \N__7945\,
            I => \REG_CYCLEm\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7942\,
            I => \REG_CYCLEm\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__7939\,
            I => \REG_CYCLEm\
        );

    \I__1575\ : IoInMux
    port map (
            O => \N__7932\,
            I => \N__7929\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__7929\,
            I => \N__7926\
        );

    \I__1573\ : IoSpan4Mux
    port map (
            O => \N__7926\,
            I => \N__7923\
        );

    \I__1572\ : IoSpan4Mux
    port map (
            O => \N__7923\,
            I => \N__7920\
        );

    \I__1571\ : Sp12to4
    port map (
            O => \N__7920\,
            I => \N__7917\
        );

    \I__1570\ : Span12Mux_v
    port map (
            O => \N__7917\,
            I => \N__7914\
        );

    \I__1569\ : Odrv12
    port map (
            O => \N__7914\,
            I => \N_160_i\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__7911\,
            I => \N__7906\
        );

    \I__1567\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7898\
        );

    \I__1566\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7898\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7906\,
            I => \N__7895\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7905\,
            I => \N__7892\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7904\,
            I => \N__7887\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7903\,
            I => \N__7887\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7898\,
            I => \N__7884\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__7895\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7892\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7887\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1557\ : Odrv12
    port map (
            O => \N__7884\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7872\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7872\,
            I => \U712_REG_SM.N_404\
        );

    \I__1554\ : IoInMux
    port map (
            O => \N__7869\,
            I => \N__7865\
        );

    \I__1553\ : IoInMux
    port map (
            O => \N__7868\,
            I => \N__7862\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7865\,
            I => \N__7858\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7862\,
            I => \N__7855\
        );

    \I__1550\ : IoInMux
    port map (
            O => \N__7861\,
            I => \N__7852\
        );

    \I__1549\ : Span4Mux_s3_v
    port map (
            O => \N__7858\,
            I => \N__7849\
        );

    \I__1548\ : Span4Mux_s1_v
    port map (
            O => \N__7855\,
            I => \N__7846\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7852\,
            I => \N__7843\
        );

    \I__1546\ : Span4Mux_v
    port map (
            O => \N__7849\,
            I => \N__7840\
        );

    \I__1545\ : Span4Mux_v
    port map (
            O => \N__7846\,
            I => \N__7837\
        );

    \I__1544\ : Span4Mux_s2_h
    port map (
            O => \N__7843\,
            I => \N__7834\
        );

    \I__1543\ : Span4Mux_h
    port map (
            O => \N__7840\,
            I => \N__7831\
        );

    \I__1542\ : Sp12to4
    port map (
            O => \N__7837\,
            I => \N__7828\
        );

    \I__1541\ : Sp12to4
    port map (
            O => \N__7834\,
            I => \N__7825\
        );

    \I__1540\ : Sp12to4
    port map (
            O => \N__7831\,
            I => \N__7822\
        );

    \I__1539\ : Span12Mux_h
    port map (
            O => \N__7828\,
            I => \N__7819\
        );

    \I__1538\ : Span12Mux_v
    port map (
            O => \N__7825\,
            I => \N__7816\
        );

    \I__1537\ : Span12Mux_v
    port map (
            O => \N__7822\,
            I => \N__7812\
        );

    \I__1536\ : Span12Mux_v
    port map (
            O => \N__7819\,
            I => \N__7807\
        );

    \I__1535\ : Span12Mux_h
    port map (
            O => \N__7816\,
            I => \N__7807\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7815\,
            I => \N__7804\
        );

    \I__1533\ : Odrv12
    port map (
            O => \N__7812\,
            I => \TACK_OUTn\
        );

    \I__1532\ : Odrv12
    port map (
            O => \N__7807\,
            I => \TACK_OUTn\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__7804\,
            I => \TACK_OUTn\
        );

    \I__1530\ : InMux
    port map (
            O => \N__7797\,
            I => \N__7793\
        );

    \I__1529\ : IoInMux
    port map (
            O => \N__7796\,
            I => \N__7790\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7793\,
            I => \N__7787\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7790\,
            I => \N__7784\
        );

    \I__1526\ : Sp12to4
    port map (
            O => \N__7787\,
            I => \N__7781\
        );

    \I__1525\ : IoSpan4Mux
    port map (
            O => \N__7784\,
            I => \N__7778\
        );

    \I__1524\ : Span12Mux_v
    port map (
            O => \N__7781\,
            I => \N__7775\
        );

    \I__1523\ : IoSpan4Mux
    port map (
            O => \N__7778\,
            I => \N__7772\
        );

    \I__1522\ : Span12Mux_h
    port map (
            O => \N__7775\,
            I => \N__7769\
        );

    \I__1521\ : IoSpan4Mux
    port map (
            O => \N__7772\,
            I => \N__7766\
        );

    \I__1520\ : Odrv12
    port map (
            O => \N__7769\,
            I => \C1_c\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__7766\,
            I => \C1_c\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7758\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__7758\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7755\,
            I => \N__7750\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7754\,
            I => \N__7747\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7734\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7750\,
            I => \N__7731\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__7747\,
            I => \N__7727\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7720\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7745\,
            I => \N__7720\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7744\,
            I => \N__7720\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7743\,
            I => \N__7714\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7742\,
            I => \N__7714\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7711\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7740\,
            I => \N__7702\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7739\,
            I => \N__7702\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__7738\,
            I => \N__7699\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7737\,
            I => \N__7688\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7734\,
            I => \N__7685\
        );

    \I__1500\ : Span4Mux_h
    port map (
            O => \N__7731\,
            I => \N__7682\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7730\,
            I => \N__7679\
        );

    \I__1498\ : Span4Mux_h
    port map (
            O => \N__7727\,
            I => \N__7674\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7720\,
            I => \N__7674\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7719\,
            I => \N__7671\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7714\,
            I => \N__7666\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7711\,
            I => \N__7666\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7661\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7709\,
            I => \N__7661\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7708\,
            I => \N__7656\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7707\,
            I => \N__7656\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7702\,
            I => \N__7653\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7699\,
            I => \N__7648\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7698\,
            I => \N__7648\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7697\,
            I => \N__7645\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7696\,
            I => \N__7640\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7695\,
            I => \N__7640\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7694\,
            I => \N__7633\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7693\,
            I => \N__7633\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7692\,
            I => \N__7633\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7691\,
            I => \N__7630\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7688\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1478\ : Odrv4
    port map (
            O => \N__7685\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__7682\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7679\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1475\ : Odrv4
    port map (
            O => \N__7674\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7671\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1473\ : Odrv12
    port map (
            O => \N__7666\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__7661\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7656\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1470\ : Odrv4
    port map (
            O => \N__7653\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7648\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7645\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__7640\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7633\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7630\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7599\,
            I => \N__7587\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7598\,
            I => \N__7584\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7597\,
            I => \N__7575\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7596\,
            I => \N__7572\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7595\,
            I => \N__7569\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7594\,
            I => \N__7562\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7593\,
            I => \N__7562\
        );

    \I__1457\ : InMux
    port map (
            O => \N__7592\,
            I => \N__7562\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7591\,
            I => \N__7557\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7590\,
            I => \N__7557\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7587\,
            I => \N__7553\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7584\,
            I => \N__7550\
        );

    \I__1452\ : CascadeMux
    port map (
            O => \N__7583\,
            I => \N__7542\
        );

    \I__1451\ : CascadeMux
    port map (
            O => \N__7582\,
            I => \N__7537\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7581\,
            I => \N__7534\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7580\,
            I => \N__7527\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7579\,
            I => \N__7527\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7578\,
            I => \N__7527\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7575\,
            I => \N__7524\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7572\,
            I => \N__7517\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__7569\,
            I => \N__7517\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7562\,
            I => \N__7517\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__7557\,
            I => \N__7514\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7556\,
            I => \N__7511\
        );

    \I__1440\ : Span4Mux_h
    port map (
            O => \N__7553\,
            I => \N__7508\
        );

    \I__1439\ : Span12Mux_v
    port map (
            O => \N__7550\,
            I => \N__7505\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7549\,
            I => \N__7500\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7548\,
            I => \N__7500\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7547\,
            I => \N__7495\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7546\,
            I => \N__7495\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7490\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7542\,
            I => \N__7490\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7541\,
            I => \N__7483\
        );

    \I__1431\ : InMux
    port map (
            O => \N__7540\,
            I => \N__7483\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7537\,
            I => \N__7483\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7534\,
            I => \N__7478\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__7527\,
            I => \N__7478\
        );

    \I__1427\ : Span4Mux_h
    port map (
            O => \N__7524\,
            I => \N__7471\
        );

    \I__1426\ : Span4Mux_v
    port map (
            O => \N__7517\,
            I => \N__7471\
        );

    \I__1425\ : Span4Mux_h
    port map (
            O => \N__7514\,
            I => \N__7471\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__7511\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__7508\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1422\ : Odrv12
    port map (
            O => \N__7505\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7500\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7495\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__7490\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__7483\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1417\ : Odrv4
    port map (
            O => \N__7478\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1416\ : Odrv4
    port map (
            O => \N__7471\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__7452\,
            I => \N__7447\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__7451\,
            I => \N__7444\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__7450\,
            I => \N__7440\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7447\,
            I => \N__7435\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7444\,
            I => \N__7432\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__7443\,
            I => \N__7429\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7440\,
            I => \N__7426\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7439\,
            I => \N__7420\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7438\,
            I => \N__7420\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7435\,
            I => \N__7415\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7432\,
            I => \N__7415\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7429\,
            I => \N__7412\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7426\,
            I => \N__7409\
        );

    \I__1402\ : InMux
    port map (
            O => \N__7425\,
            I => \N__7405\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7420\,
            I => \N__7402\
        );

    \I__1400\ : Span4Mux_h
    port map (
            O => \N__7415\,
            I => \N__7397\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7412\,
            I => \N__7397\
        );

    \I__1398\ : Span4Mux_h
    port map (
            O => \N__7409\,
            I => \N__7394\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7408\,
            I => \N__7391\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7405\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1395\ : Odrv4
    port map (
            O => \N__7402\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__7397\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__7394\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7391\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7380\,
            I => \N__7375\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7379\,
            I => \N__7372\
        );

    \I__1389\ : InMux
    port map (
            O => \N__7378\,
            I => \N__7368\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__7375\,
            I => \N__7364\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7372\,
            I => \N__7361\
        );

    \I__1386\ : InMux
    port map (
            O => \N__7371\,
            I => \N__7358\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7368\,
            I => \N__7355\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7367\,
            I => \N__7352\
        );

    \I__1383\ : Odrv4
    port map (
            O => \N__7364\,
            I => \U712_CHIP_RAM.N_466\
        );

    \I__1382\ : Odrv4
    port map (
            O => \N__7361\,
            I => \U712_CHIP_RAM.N_466\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__7358\,
            I => \U712_CHIP_RAM.N_466\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__7355\,
            I => \U712_CHIP_RAM.N_466\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__7352\,
            I => \U712_CHIP_RAM.N_466\
        );

    \I__1378\ : CEMux
    port map (
            O => \N__7341\,
            I => \N__7338\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7338\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7335\,
            I => \N__7332\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__7332\,
            I => \N__7329\
        );

    \I__1374\ : Span4Mux_v
    port map (
            O => \N__7329\,
            I => \N__7326\
        );

    \I__1373\ : Sp12to4
    port map (
            O => \N__7326\,
            I => \N__7323\
        );

    \I__1372\ : Span12Mux_h
    port map (
            O => \N__7323\,
            I => \N__7320\
        );

    \I__1371\ : Span12Mux_v
    port map (
            O => \N__7320\,
            I => \N__7317\
        );

    \I__1370\ : Odrv12
    port map (
            O => \N__7317\,
            I => \REGSPACEn_c\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7314\,
            I => \N__7310\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7313\,
            I => \N__7307\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7310\,
            I => \N__7304\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__7307\,
            I => \N__7301\
        );

    \I__1365\ : Span4Mux_v
    port map (
            O => \N__7304\,
            I => \N__7298\
        );

    \I__1364\ : Span4Mux_v
    port map (
            O => \N__7301\,
            I => \N__7295\
        );

    \I__1363\ : Sp12to4
    port map (
            O => \N__7298\,
            I => \N__7290\
        );

    \I__1362\ : Sp12to4
    port map (
            O => \N__7295\,
            I => \N__7290\
        );

    \I__1361\ : Span12Mux_h
    port map (
            O => \N__7290\,
            I => \N__7287\
        );

    \I__1360\ : Span12Mux_v
    port map (
            O => \N__7287\,
            I => \N__7284\
        );

    \I__1359\ : Odrv12
    port map (
            O => \N__7284\,
            I => \TSn_c\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__7281\,
            I => \U712_REG_SM.N_401_cascade_\
        );

    \I__1357\ : InMux
    port map (
            O => \N__7278\,
            I => \N__7271\
        );

    \I__1356\ : InMux
    port map (
            O => \N__7277\,
            I => \N__7271\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7276\,
            I => \N__7267\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7271\,
            I => \N__7264\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7270\,
            I => \N__7261\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__7267\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1351\ : Odrv4
    port map (
            O => \N__7264\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__7261\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7254\,
            I => \N__7250\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7253\,
            I => \N__7247\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__7250\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7247\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__7242\,
            I => \N__7238\
        );

    \I__1344\ : InMux
    port map (
            O => \N__7241\,
            I => \N__7233\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7230\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7237\,
            I => \N__7227\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7236\,
            I => \N__7224\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__7233\,
            I => \N__7221\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__7230\,
            I => \N__7216\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__7227\,
            I => \N__7216\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__7224\,
            I => \N__7212\
        );

    \I__1336\ : Span4Mux_h
    port map (
            O => \N__7221\,
            I => \N__7209\
        );

    \I__1335\ : Span4Mux_h
    port map (
            O => \N__7216\,
            I => \N__7206\
        );

    \I__1334\ : InMux
    port map (
            O => \N__7215\,
            I => \N__7203\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__7212\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1332\ : Odrv4
    port map (
            O => \N__7209\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1331\ : Odrv4
    port map (
            O => \N__7206\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__7203\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__7194\,
            I => \U712_REG_SM.N_324_cascade_\
        );

    \I__1328\ : InMux
    port map (
            O => \N__7191\,
            I => \N__7188\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__7188\,
            I => \N__7184\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7187\,
            I => \N__7179\
        );

    \I__1325\ : Span4Mux_v
    port map (
            O => \N__7184\,
            I => \N__7176\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7183\,
            I => \N__7171\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7182\,
            I => \N__7171\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__7179\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__7176\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__7171\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1319\ : InMux
    port map (
            O => \N__7164\,
            I => \N__7161\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__7161\,
            I => \U712_REG_SM.STATE_COUNTc_0_0\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7158\,
            I => \N__7154\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7157\,
            I => \N__7151\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__7154\,
            I => \U712_BYTE_ENABLE.N_424\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__7151\,
            I => \U712_BYTE_ENABLE.N_424\
        );

    \I__1313\ : InMux
    port map (
            O => \N__7146\,
            I => \N__7142\
        );

    \I__1312\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7139\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7142\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__7139\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0\
        );

    \I__1309\ : IoInMux
    port map (
            O => \N__7134\,
            I => \N__7131\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__7131\,
            I => \N__7128\
        );

    \I__1307\ : IoSpan4Mux
    port map (
            O => \N__7128\,
            I => \N__7125\
        );

    \I__1306\ : IoSpan4Mux
    port map (
            O => \N__7125\,
            I => \N__7122\
        );

    \I__1305\ : Sp12to4
    port map (
            O => \N__7122\,
            I => \N__7119\
        );

    \I__1304\ : Span12Mux_s7_v
    port map (
            O => \N__7119\,
            I => \N__7116\
        );

    \I__1303\ : Span12Mux_h
    port map (
            O => \N__7116\,
            I => \N__7113\
        );

    \I__1302\ : Odrv12
    port map (
            O => \N__7113\,
            I => \N_170_i\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7110\,
            I => \N__7107\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__7107\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1299\ : IoInMux
    port map (
            O => \N__7104\,
            I => \N__7101\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__7101\,
            I => \N__7098\
        );

    \I__1297\ : Span12Mux_s6_v
    port map (
            O => \N__7098\,
            I => \N__7095\
        );

    \I__1296\ : Odrv12
    port map (
            O => \N__7095\,
            I => \CMA_c_2\
        );

    \I__1295\ : InMux
    port map (
            O => \N__7092\,
            I => \N__7089\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__7089\,
            I => \N__7086\
        );

    \I__1293\ : Span4Mux_v
    port map (
            O => \N__7086\,
            I => \N__7083\
        );

    \I__1292\ : Span4Mux_h
    port map (
            O => \N__7083\,
            I => \N__7080\
        );

    \I__1291\ : Sp12to4
    port map (
            O => \N__7080\,
            I => \N__7077\
        );

    \I__1290\ : Odrv12
    port map (
            O => \N__7077\,
            I => \A_c_7\
        );

    \I__1289\ : InMux
    port map (
            O => \N__7074\,
            I => \N__7070\
        );

    \I__1288\ : InMux
    port map (
            O => \N__7073\,
            I => \N__7067\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__7070\,
            I => \N__7064\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__7067\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\
        );

    \I__1285\ : Odrv4
    port map (
            O => \N__7064\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\
        );

    \I__1284\ : InMux
    port map (
            O => \N__7059\,
            I => \N__7056\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__7056\,
            I => \N__7053\
        );

    \I__1282\ : Span12Mux_h
    port map (
            O => \N__7053\,
            I => \N__7050\
        );

    \I__1281\ : Span12Mux_v
    port map (
            O => \N__7050\,
            I => \N__7047\
        );

    \I__1280\ : Odrv12
    port map (
            O => \N__7047\,
            I => \A_c_2\
        );

    \I__1279\ : InMux
    port map (
            O => \N__7044\,
            I => \N__7040\
        );

    \I__1278\ : InMux
    port map (
            O => \N__7043\,
            I => \N__7037\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__7040\,
            I => \N__7034\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__7037\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__7034\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\
        );

    \I__1274\ : InMux
    port map (
            O => \N__7029\,
            I => \N__7026\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__7026\,
            I => \N__7023\
        );

    \I__1272\ : Span4Mux_v
    port map (
            O => \N__7023\,
            I => \N__7020\
        );

    \I__1271\ : Sp12to4
    port map (
            O => \N__7020\,
            I => \N__7017\
        );

    \I__1270\ : Span12Mux_h
    port map (
            O => \N__7017\,
            I => \N__7014\
        );

    \I__1269\ : Odrv12
    port map (
            O => \N__7014\,
            I => \A_c_8\
        );

    \I__1268\ : InMux
    port map (
            O => \N__7011\,
            I => \N__7008\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__7008\,
            I => \N__6997\
        );

    \I__1266\ : InMux
    port map (
            O => \N__7007\,
            I => \N__6994\
        );

    \I__1265\ : InMux
    port map (
            O => \N__7006\,
            I => \N__6987\
        );

    \I__1264\ : InMux
    port map (
            O => \N__7005\,
            I => \N__6987\
        );

    \I__1263\ : InMux
    port map (
            O => \N__7004\,
            I => \N__6987\
        );

    \I__1262\ : InMux
    port map (
            O => \N__7003\,
            I => \N__6984\
        );

    \I__1261\ : InMux
    port map (
            O => \N__7002\,
            I => \N__6977\
        );

    \I__1260\ : InMux
    port map (
            O => \N__7001\,
            I => \N__6977\
        );

    \I__1259\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6977\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__6997\,
            I => \N__6974\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6994\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__6987\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__6984\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6977\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__6974\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__1252\ : IoInMux
    port map (
            O => \N__6963\,
            I => \N__6960\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__6960\,
            I => \N__6957\
        );

    \I__1250\ : IoSpan4Mux
    port map (
            O => \N__6957\,
            I => \N__6954\
        );

    \I__1249\ : Span4Mux_s2_h
    port map (
            O => \N__6954\,
            I => \N__6951\
        );

    \I__1248\ : Sp12to4
    port map (
            O => \N__6951\,
            I => \N__6948\
        );

    \I__1247\ : Span12Mux_s11_h
    port map (
            O => \N__6948\,
            I => \N__6945\
        );

    \I__1246\ : Span12Mux_v
    port map (
            O => \N__6945\,
            I => \N__6942\
        );

    \I__1245\ : Odrv12
    port map (
            O => \N__6942\,
            I => \CMA_c_4\
        );

    \I__1244\ : IoInMux
    port map (
            O => \N__6939\,
            I => \N__6936\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__6936\,
            I => \N__6933\
        );

    \I__1242\ : IoSpan4Mux
    port map (
            O => \N__6933\,
            I => \N__6930\
        );

    \I__1241\ : Span4Mux_s3_h
    port map (
            O => \N__6930\,
            I => \N__6927\
        );

    \I__1240\ : Sp12to4
    port map (
            O => \N__6927\,
            I => \N__6924\
        );

    \I__1239\ : Span12Mux_h
    port map (
            O => \N__6924\,
            I => \N__6921\
        );

    \I__1238\ : Span12Mux_v
    port map (
            O => \N__6921\,
            I => \N__6918\
        );

    \I__1237\ : Odrv12
    port map (
            O => \N__6918\,
            I => \CMA_c_3\
        );

    \I__1236\ : IoInMux
    port map (
            O => \N__6915\,
            I => \N__6912\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6912\,
            I => \N__6909\
        );

    \I__1234\ : Span12Mux_s7_h
    port map (
            O => \N__6909\,
            I => \N__6906\
        );

    \I__1233\ : Span12Mux_v
    port map (
            O => \N__6906\,
            I => \N__6903\
        );

    \I__1232\ : Odrv12
    port map (
            O => \N__6903\,
            I => \CMA_c_6\
        );

    \I__1231\ : CascadeMux
    port map (
            O => \N__6900\,
            I => \N__6895\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__6899\,
            I => \N__6889\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__6898\,
            I => \N__6886\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6895\,
            I => \N__6883\
        );

    \I__1227\ : CascadeMux
    port map (
            O => \N__6894\,
            I => \N__6880\
        );

    \I__1226\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6870\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6892\,
            I => \N__6870\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6889\,
            I => \N__6870\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6886\,
            I => \N__6870\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__6883\,
            I => \N__6867\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6864\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6879\,
            I => \N__6861\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6870\,
            I => \N__6858\
        );

    \I__1218\ : Span4Mux_h
    port map (
            O => \N__6867\,
            I => \N__6855\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__6864\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__6861\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1215\ : Odrv4
    port map (
            O => \N__6858\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__6855\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6843\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6843\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1211\ : IoInMux
    port map (
            O => \N__6840\,
            I => \N__6837\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6837\,
            I => \N__6834\
        );

    \I__1209\ : IoSpan4Mux
    port map (
            O => \N__6834\,
            I => \N__6831\
        );

    \I__1208\ : IoSpan4Mux
    port map (
            O => \N__6831\,
            I => \N__6828\
        );

    \I__1207\ : Span4Mux_s3_h
    port map (
            O => \N__6828\,
            I => \N__6825\
        );

    \I__1206\ : Sp12to4
    port map (
            O => \N__6825\,
            I => \N__6822\
        );

    \I__1205\ : Span12Mux_h
    port map (
            O => \N__6822\,
            I => \N__6819\
        );

    \I__1204\ : Odrv12
    port map (
            O => \N__6819\,
            I => \CMA_c_7\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6816\,
            I => \N__6812\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6815\,
            I => \N__6809\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6812\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_5\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6809\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_5\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6804\,
            I => \N__6800\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6803\,
            I => \N__6797\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6800\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_4\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__6797\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_4\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__6792\,
            I => \N__6788\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6785\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6782\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6785\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_3\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__6782\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_3\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6773\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6770\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6773\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_7\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__6770\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_7\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6762\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6762\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_5_i_a2_5\
        );

    \I__1184\ : IoInMux
    port map (
            O => \N__6759\,
            I => \N__6756\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6756\,
            I => \N__6753\
        );

    \I__1182\ : IoSpan4Mux
    port map (
            O => \N__6753\,
            I => \N__6750\
        );

    \I__1181\ : Span4Mux_s3_v
    port map (
            O => \N__6750\,
            I => \N__6747\
        );

    \I__1180\ : Span4Mux_v
    port map (
            O => \N__6747\,
            I => \N__6744\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__6744\,
            I => \DMA_LATCH_EN_c\
        );

    \I__1178\ : IoInMux
    port map (
            O => \N__6741\,
            I => \N__6738\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6738\,
            I => \N__6735\
        );

    \I__1176\ : Span4Mux_s3_v
    port map (
            O => \N__6735\,
            I => \N__6732\
        );

    \I__1175\ : Span4Mux_h
    port map (
            O => \N__6732\,
            I => \N__6729\
        );

    \I__1174\ : Sp12to4
    port map (
            O => \N__6729\,
            I => \N__6726\
        );

    \I__1173\ : Span12Mux_v
    port map (
            O => \N__6726\,
            I => \N__6723\
        );

    \I__1172\ : Odrv12
    port map (
            O => \N__6723\,
            I => \CMA_c_10\
        );

    \I__1171\ : IoInMux
    port map (
            O => \N__6720\,
            I => \N__6716\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6713\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6716\,
            I => \N__6710\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6713\,
            I => \N__6707\
        );

    \I__1167\ : Span12Mux_s4_v
    port map (
            O => \N__6710\,
            I => \N__6704\
        );

    \I__1166\ : Span4Mux_v
    port map (
            O => \N__6707\,
            I => \N__6701\
        );

    \I__1165\ : Span12Mux_h
    port map (
            O => \N__6704\,
            I => \N__6698\
        );

    \I__1164\ : Span4Mux_h
    port map (
            O => \N__6701\,
            I => \N__6695\
        );

    \I__1163\ : Span12Mux_v
    port map (
            O => \N__6698\,
            I => \N__6692\
        );

    \I__1162\ : Sp12to4
    port map (
            O => \N__6695\,
            I => \N__6689\
        );

    \I__1161\ : Odrv12
    port map (
            O => \N__6692\,
            I => \A_c_9\
        );

    \I__1160\ : Odrv12
    port map (
            O => \N__6689\,
            I => \A_c_9\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__6684\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__6681\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_\
        );

    \I__1157\ : IoInMux
    port map (
            O => \N__6678\,
            I => \N__6675\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6675\,
            I => \N__6672\
        );

    \I__1155\ : Span4Mux_s3_v
    port map (
            O => \N__6672\,
            I => \N__6669\
        );

    \I__1154\ : Sp12to4
    port map (
            O => \N__6669\,
            I => \N__6666\
        );

    \I__1153\ : Span12Mux_h
    port map (
            O => \N__6666\,
            I => \N__6663\
        );

    \I__1152\ : Odrv12
    port map (
            O => \N__6663\,
            I => \CMA_c_0\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__6660\,
            I => \U712_REG_SM.N_408_cascade_\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6657\,
            I => \N__6654\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6654\,
            I => \U712_REG_SM.N_367\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6648\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6648\,
            I => \U712_REG_SM.N_410\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6645\,
            I => \N__6641\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6644\,
            I => \N__6638\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6641\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6638\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6633\,
            I => \N__6630\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__6630\,
            I => \U712_REG_SM.REGENn_e_1\
        );

    \I__1140\ : IoInMux
    port map (
            O => \N__6627\,
            I => \N__6624\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6624\,
            I => \N__6621\
        );

    \I__1138\ : Span4Mux_s0_v
    port map (
            O => \N__6621\,
            I => \N__6618\
        );

    \I__1137\ : Sp12to4
    port map (
            O => \N__6618\,
            I => \N__6615\
        );

    \I__1136\ : Span12Mux_s7_h
    port map (
            O => \N__6615\,
            I => \N__6612\
        );

    \I__1135\ : Span12Mux_v
    port map (
            O => \N__6612\,
            I => \N__6607\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6611\,
            I => \N__6604\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6601\
        );

    \I__1132\ : Odrv12
    port map (
            O => \N__6607\,
            I => \REGENn_c\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6604\,
            I => \REGENn_c\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__6601\,
            I => \REGENn_c\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6588\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6593\,
            I => \N__6588\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__6588\,
            I => \U712_REG_SM.N_322\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6585\,
            I => \N__6582\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6582\,
            I => \U712_REG_SM.N_131\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6579\,
            I => \N__6576\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6576\,
            I => \N__6573\
        );

    \I__1122\ : Span4Mux_v
    port map (
            O => \N__6573\,
            I => \N__6568\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6563\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6563\
        );

    \I__1119\ : Odrv4
    port map (
            O => \N__6568\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6563\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__6558\,
            I => \N__6554\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6557\,
            I => \N__6548\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6548\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6553\,
            I => \N__6545\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__6548\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_1\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6545\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_1\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6540\,
            I => \N__6536\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6539\,
            I => \N__6533\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6536\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_6\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6533\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_6\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6528\,
            I => \N__6524\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6527\,
            I => \N__6521\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6524\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_2\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6521\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_2\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6516\,
            I => \N__6510\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6515\,
            I => \N__6507\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6514\,
            I => \N__6502\
        );

    \I__1100\ : InMux
    port map (
            O => \N__6513\,
            I => \N__6502\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6510\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__6507\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__6502\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__6495\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_5_i_a2_4_cascade_\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__6492\,
            I => \N__6489\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6489\,
            I => \N__6486\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6486\,
            I => \N__6483\
        );

    \I__1092\ : Span4Mux_h
    port map (
            O => \N__6483\,
            I => \N__6480\
        );

    \I__1091\ : Odrv4
    port map (
            O => \N__6480\,
            I => \U712_CHIP_RAM.N_456\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__6477\,
            I => \U712_CHIP_RAM.N_419_cascade_\
        );

    \I__1089\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6471\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__6471\,
            I => \N__6468\
        );

    \I__1087\ : Span4Mux_v
    port map (
            O => \N__6468\,
            I => \N__6465\
        );

    \I__1086\ : Span4Mux_h
    port map (
            O => \N__6465\,
            I => \N__6462\
        );

    \I__1085\ : Sp12to4
    port map (
            O => \N__6462\,
            I => \N__6459\
        );

    \I__1084\ : Odrv12
    port map (
            O => \N__6459\,
            I => \RAMSPACEn_c\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__6456\,
            I => \N__6453\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6453\,
            I => \N__6450\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__6450\,
            I => \N__6445\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6449\,
            I => \N__6442\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6448\,
            I => \N__6438\
        );

    \I__1078\ : Span4Mux_v
    port map (
            O => \N__6445\,
            I => \N__6435\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__6442\,
            I => \N__6432\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6441\,
            I => \N__6429\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6438\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1074\ : Odrv4
    port map (
            O => \N__6435\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1073\ : Odrv4
    port map (
            O => \N__6432\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__6429\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__6420\,
            I => \N__6415\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6419\,
            I => \N__6411\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__6418\,
            I => \N__6408\
        );

    \I__1068\ : InMux
    port map (
            O => \N__6415\,
            I => \N__6405\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__6414\,
            I => \N__6401\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6411\,
            I => \N__6398\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6408\,
            I => \N__6394\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__6405\,
            I => \N__6391\
        );

    \I__1063\ : CascadeMux
    port map (
            O => \N__6404\,
            I => \N__6386\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6401\,
            I => \N__6380\
        );

    \I__1061\ : Span4Mux_v
    port map (
            O => \N__6398\,
            I => \N__6372\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6369\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6394\,
            I => \N__6364\
        );

    \I__1058\ : Span4Mux_v
    port map (
            O => \N__6391\,
            I => \N__6364\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6359\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6389\,
            I => \N__6359\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6386\,
            I => \N__6352\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6352\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6384\,
            I => \N__6352\
        );

    \I__1052\ : InMux
    port map (
            O => \N__6383\,
            I => \N__6349\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6380\,
            I => \N__6346\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6379\,
            I => \N__6343\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6378\,
            I => \N__6338\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6377\,
            I => \N__6338\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6376\,
            I => \N__6333\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6375\,
            I => \N__6333\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__6372\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__6369\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1043\ : Odrv4
    port map (
            O => \N__6364\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6359\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__6352\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6349\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1039\ : Odrv4
    port map (
            O => \N__6346\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6343\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6338\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6333\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6308\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6305\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6308\,
            I => \U712_CHIP_RAM.N_299\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6305\,
            I => \U712_CHIP_RAM.N_299\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6300\,
            I => \N__6297\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6297\,
            I => \N__6293\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__6296\,
            I => \N__6290\
        );

    \I__1028\ : Span4Mux_h
    port map (
            O => \N__6293\,
            I => \N__6287\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6290\,
            I => \N__6284\
        );

    \I__1026\ : Odrv4
    port map (
            O => \N__6287\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__6284\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6279\,
            I => \N__6276\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__6276\,
            I => \U712_CHIP_RAM.N_434\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6273\,
            I => \N__6270\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__6270\,
            I => \N__6266\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6263\
        );

    \I__1019\ : Span4Mux_h
    port map (
            O => \N__6266\,
            I => \N__6260\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__6263\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1017\ : Odrv4
    port map (
            O => \N__6260\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6255\,
            I => \N__6252\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6252\,
            I => \U712_CHIP_RAM.REFRESH5lto7_0\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6246\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__6246\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__1012\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6238\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6242\,
            I => \N__6233\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6233\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6238\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6233\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__6228\,
            I => \U712_REG_SM.N_322_cascade_\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__6225\,
            I => \U712_REG_SM.N_367_cascade_\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__6222\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6219\,
            I => \N__6216\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6216\,
            I => \N__6212\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6215\,
            I => \N__6209\
        );

    \I__1001\ : Span4Mux_v
    port map (
            O => \N__6212\,
            I => \N__6204\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__6209\,
            I => \N__6204\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__6204\,
            I => \U712_CHIP_RAM.N_429\
        );

    \I__998\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6198\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__6198\,
            I => \N__6195\
        );

    \I__996\ : Odrv4
    port map (
            O => \N__6195\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__6192\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_cascade_\
        );

    \I__994\ : InMux
    port map (
            O => \N__6189\,
            I => \N__6186\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__6186\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__992\ : InMux
    port map (
            O => \N__6183\,
            I => \N__6179\
        );

    \I__991\ : InMux
    port map (
            O => \N__6182\,
            I => \N__6176\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__6179\,
            I => \U712_CHIP_RAM.N_319\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__6176\,
            I => \U712_CHIP_RAM.N_319\
        );

    \I__988\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6168\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__6168\,
            I => \N__6165\
        );

    \I__986\ : Odrv12
    port map (
            O => \N__6165\,
            I => \U712_CHIP_RAM.N_359\
        );

    \I__985\ : InMux
    port map (
            O => \N__6162\,
            I => \N__6158\
        );

    \I__984\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6155\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__6158\,
            I => \N__6151\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__6155\,
            I => \N__6148\
        );

    \I__981\ : InMux
    port map (
            O => \N__6154\,
            I => \N__6145\
        );

    \I__980\ : Span4Mux_v
    port map (
            O => \N__6151\,
            I => \N__6142\
        );

    \I__979\ : Span4Mux_h
    port map (
            O => \N__6148\,
            I => \N__6137\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__6145\,
            I => \N__6137\
        );

    \I__977\ : Sp12to4
    port map (
            O => \N__6142\,
            I => \N__6134\
        );

    \I__976\ : Span4Mux_v
    port map (
            O => \N__6137\,
            I => \N__6131\
        );

    \I__975\ : Span12Mux_h
    port map (
            O => \N__6134\,
            I => \N__6128\
        );

    \I__974\ : Span4Mux_h
    port map (
            O => \N__6131\,
            I => \N__6125\
        );

    \I__973\ : Span12Mux_v
    port map (
            O => \N__6128\,
            I => \N__6122\
        );

    \I__972\ : Sp12to4
    port map (
            O => \N__6125\,
            I => \N__6119\
        );

    \I__971\ : Odrv12
    port map (
            O => \N__6122\,
            I => \AWEn_c\
        );

    \I__970\ : Odrv12
    port map (
            O => \N__6119\,
            I => \AWEn_c\
        );

    \I__969\ : InMux
    port map (
            O => \N__6114\,
            I => \N__6110\
        );

    \I__968\ : InMux
    port map (
            O => \N__6113\,
            I => \N__6107\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__6110\,
            I => \N__6104\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__6107\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__965\ : Odrv4
    port map (
            O => \N__6104\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__964\ : InMux
    port map (
            O => \N__6099\,
            I => \N__6096\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__6096\,
            I => \N__6093\
        );

    \I__962\ : Span4Mux_h
    port map (
            O => \N__6093\,
            I => \N__6089\
        );

    \I__961\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6086\
        );

    \I__960\ : Odrv4
    port map (
            O => \N__6089\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0_a2_0\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__6086\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0_a2_0\
        );

    \I__958\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6077\
        );

    \I__957\ : InMux
    port map (
            O => \N__6080\,
            I => \N__6074\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__6077\,
            I => \N__6071\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__6074\,
            I => \N__6068\
        );

    \I__954\ : Span4Mux_v
    port map (
            O => \N__6071\,
            I => \N__6062\
        );

    \I__953\ : Span4Mux_v
    port map (
            O => \N__6068\,
            I => \N__6062\
        );

    \I__952\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6059\
        );

    \I__951\ : Odrv4
    port map (
            O => \N__6062\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__6059\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__949\ : IoInMux
    port map (
            O => \N__6054\,
            I => \N__6051\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__6051\,
            I => \N__6048\
        );

    \I__947\ : IoSpan4Mux
    port map (
            O => \N__6048\,
            I => \N__6045\
        );

    \I__946\ : Span4Mux_s0_v
    port map (
            O => \N__6045\,
            I => \N__6042\
        );

    \I__945\ : Sp12to4
    port map (
            O => \N__6042\,
            I => \N__6039\
        );

    \I__944\ : Span12Mux_v
    port map (
            O => \N__6039\,
            I => \N__6035\
        );

    \I__943\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6032\
        );

    \I__942\ : Odrv12
    port map (
            O => \N__6035\,
            I => \DBDIR_c\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__6032\,
            I => \DBDIR_c\
        );

    \I__940\ : InMux
    port map (
            O => \N__6027\,
            I => \N__6024\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__6024\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i\
        );

    \I__938\ : InMux
    port map (
            O => \N__6021\,
            I => \N__6018\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__6018\,
            I => \N__6015\
        );

    \I__936\ : Span12Mux_v
    port map (
            O => \N__6015\,
            I => \N__6012\
        );

    \I__935\ : Span12Mux_h
    port map (
            O => \N__6012\,
            I => \N__6009\
        );

    \I__934\ : Odrv12
    port map (
            O => \N__6009\,
            I => \A_c_12\
        );

    \I__933\ : InMux
    port map (
            O => \N__6006\,
            I => \N__6003\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__6003\,
            I => \N__6000\
        );

    \I__931\ : Span4Mux_h
    port map (
            O => \N__6000\,
            I => \N__5997\
        );

    \I__930\ : Span4Mux_v
    port map (
            O => \N__5997\,
            I => \N__5994\
        );

    \I__929\ : Sp12to4
    port map (
            O => \N__5994\,
            I => \N__5991\
        );

    \I__928\ : Odrv12
    port map (
            O => \N__5991\,
            I => \A_c_5\
        );

    \I__927\ : InMux
    port map (
            O => \N__5988\,
            I => \N__5982\
        );

    \I__926\ : InMux
    port map (
            O => \N__5987\,
            I => \N__5982\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__5982\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\
        );

    \I__924\ : InMux
    port map (
            O => \N__5979\,
            I => \N__5975\
        );

    \I__923\ : InMux
    port map (
            O => \N__5978\,
            I => \N__5971\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__5975\,
            I => \N__5968\
        );

    \I__921\ : InMux
    port map (
            O => \N__5974\,
            I => \N__5965\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__5971\,
            I => \U712_CHIP_RAM.N_471\
        );

    \I__919\ : Odrv4
    port map (
            O => \N__5968\,
            I => \U712_CHIP_RAM.N_471\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5965\,
            I => \U712_CHIP_RAM.N_471\
        );

    \I__917\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5955\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5955\,
            I => \N__5952\
        );

    \I__915\ : Span12Mux_v
    port map (
            O => \N__5952\,
            I => \N__5949\
        );

    \I__914\ : Span12Mux_h
    port map (
            O => \N__5949\,
            I => \N__5946\
        );

    \I__913\ : Odrv12
    port map (
            O => \N__5946\,
            I => \A_c_3\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__5943\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\
        );

    \I__911\ : InMux
    port map (
            O => \N__5940\,
            I => \N__5937\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__5937\,
            I => \N__5934\
        );

    \I__909\ : Span12Mux_v
    port map (
            O => \N__5934\,
            I => \N__5931\
        );

    \I__908\ : Span12Mux_h
    port map (
            O => \N__5931\,
            I => \N__5928\
        );

    \I__907\ : Odrv12
    port map (
            O => \N__5928\,
            I => \A_c_4\
        );

    \I__906\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5921\
        );

    \I__905\ : InMux
    port map (
            O => \N__5924\,
            I => \N__5918\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5921\,
            I => \N__5915\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5918\,
            I => \N__5912\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__5915\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\
        );

    \I__901\ : Odrv4
    port map (
            O => \N__5912\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\
        );

    \I__900\ : InMux
    port map (
            O => \N__5907\,
            I => \N__5904\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__5904\,
            I => \N__5901\
        );

    \I__898\ : Span4Mux_v
    port map (
            O => \N__5901\,
            I => \N__5898\
        );

    \I__897\ : Sp12to4
    port map (
            O => \N__5898\,
            I => \N__5895\
        );

    \I__896\ : Span12Mux_h
    port map (
            O => \N__5895\,
            I => \N__5892\
        );

    \I__895\ : Odrv12
    port map (
            O => \N__5892\,
            I => \A_c_6\
        );

    \I__894\ : SRMux
    port map (
            O => \N__5889\,
            I => \N__5885\
        );

    \I__893\ : SRMux
    port map (
            O => \N__5888\,
            I => \N__5882\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5885\,
            I => \N__5879\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__5882\,
            I => \N__5876\
        );

    \I__890\ : Odrv4
    port map (
            O => \N__5879\,
            I => \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\
        );

    \I__889\ : Odrv4
    port map (
            O => \N__5876\,
            I => \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\
        );

    \I__888\ : IoInMux
    port map (
            O => \N__5871\,
            I => \N__5867\
        );

    \I__887\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5864\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5867\,
            I => \N__5861\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5864\,
            I => \N__5858\
        );

    \I__884\ : IoSpan4Mux
    port map (
            O => \N__5861\,
            I => \N__5855\
        );

    \I__883\ : Span4Mux_v
    port map (
            O => \N__5858\,
            I => \N__5852\
        );

    \I__882\ : Span4Mux_s3_v
    port map (
            O => \N__5855\,
            I => \N__5849\
        );

    \I__881\ : Span4Mux_v
    port map (
            O => \N__5852\,
            I => \N__5846\
        );

    \I__880\ : Span4Mux_v
    port map (
            O => \N__5849\,
            I => \N__5843\
        );

    \I__879\ : Odrv4
    port map (
            O => \N__5846\,
            I => \CONSTANT_ONE_NET\
        );

    \I__878\ : Odrv4
    port map (
            O => \N__5843\,
            I => \CONSTANT_ONE_NET\
        );

    \I__877\ : IoInMux
    port map (
            O => \N__5838\,
            I => \N__5835\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5835\,
            I => \N__5832\
        );

    \I__875\ : IoSpan4Mux
    port map (
            O => \N__5832\,
            I => \N__5829\
        );

    \I__874\ : Span4Mux_s0_v
    port map (
            O => \N__5829\,
            I => \N__5826\
        );

    \I__873\ : Sp12to4
    port map (
            O => \N__5826\,
            I => \N__5823\
        );

    \I__872\ : Span12Mux_h
    port map (
            O => \N__5823\,
            I => \N__5820\
        );

    \I__871\ : Span12Mux_v
    port map (
            O => \N__5820\,
            I => \N__5817\
        );

    \I__870\ : Odrv12
    port map (
            O => \N__5817\,
            I => \CMA_c_5\
        );

    \I__869\ : IoInMux
    port map (
            O => \N__5814\,
            I => \N__5811\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5811\,
            I => \N__5808\
        );

    \I__867\ : IoSpan4Mux
    port map (
            O => \N__5808\,
            I => \N__5805\
        );

    \I__866\ : Span4Mux_s2_v
    port map (
            O => \N__5805\,
            I => \N__5801\
        );

    \I__865\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5798\
        );

    \I__864\ : Sp12to4
    port map (
            O => \N__5801\,
            I => \N__5795\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5798\,
            I => \N__5792\
        );

    \I__862\ : Span12Mux_s8_v
    port map (
            O => \N__5795\,
            I => \N__5789\
        );

    \I__861\ : Span4Mux_v
    port map (
            O => \N__5792\,
            I => \N__5786\
        );

    \I__860\ : Span12Mux_v
    port map (
            O => \N__5789\,
            I => \N__5783\
        );

    \I__859\ : Sp12to4
    port map (
            O => \N__5786\,
            I => \N__5780\
        );

    \I__858\ : Span12Mux_h
    port map (
            O => \N__5783\,
            I => \N__5777\
        );

    \I__857\ : Span12Mux_h
    port map (
            O => \N__5780\,
            I => \N__5774\
        );

    \I__856\ : Odrv12
    port map (
            O => \N__5777\,
            I => \A_c_11\
        );

    \I__855\ : Odrv12
    port map (
            O => \N__5774\,
            I => \A_c_11\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__5769\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\
        );

    \I__853\ : InMux
    port map (
            O => \N__5766\,
            I => \N__5763\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5763\,
            I => \N__5760\
        );

    \I__851\ : Span4Mux_v
    port map (
            O => \N__5760\,
            I => \N__5757\
        );

    \I__850\ : Span4Mux_v
    port map (
            O => \N__5757\,
            I => \N__5754\
        );

    \I__849\ : Span4Mux_v
    port map (
            O => \N__5754\,
            I => \N__5751\
        );

    \I__848\ : Sp12to4
    port map (
            O => \N__5751\,
            I => \N__5748\
        );

    \I__847\ : Span12Mux_h
    port map (
            O => \N__5748\,
            I => \N__5745\
        );

    \I__846\ : Odrv12
    port map (
            O => \N__5745\,
            I => \A_c_17\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__5742\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\
        );

    \I__844\ : InMux
    port map (
            O => \N__5739\,
            I => \N__5735\
        );

    \I__843\ : InMux
    port map (
            O => \N__5738\,
            I => \N__5732\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5735\,
            I => \N__5729\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5732\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__5729\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__839\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5721\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5721\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\
        );

    \I__837\ : InMux
    port map (
            O => \N__5718\,
            I => \N__5715\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__5715\,
            I => \N__5712\
        );

    \I__835\ : Span12Mux_v
    port map (
            O => \N__5712\,
            I => \N__5709\
        );

    \I__834\ : Span12Mux_h
    port map (
            O => \N__5709\,
            I => \N__5706\
        );

    \I__833\ : Odrv12
    port map (
            O => \N__5706\,
            I => \A_c_14\
        );

    \I__832\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5700\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5700\,
            I => \U712_CHIP_RAM.N_353\
        );

    \I__830\ : InMux
    port map (
            O => \N__5697\,
            I => \N__5694\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__5694\,
            I => \N__5691\
        );

    \I__828\ : Span12Mux_v
    port map (
            O => \N__5691\,
            I => \N__5688\
        );

    \I__827\ : Span12Mux_h
    port map (
            O => \N__5688\,
            I => \N__5685\
        );

    \I__826\ : Odrv12
    port map (
            O => \N__5685\,
            I => \A_c_20\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__5682\,
            I => \N__5679\
        );

    \I__824\ : InMux
    port map (
            O => \N__5679\,
            I => \N__5675\
        );

    \I__823\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5672\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5675\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5672\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__5667\,
            I => \N__5664\
        );

    \I__819\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5661\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5661\,
            I => \U712_CHIP_RAM.DBENn_7_0_0\
        );

    \I__817\ : InMux
    port map (
            O => \N__5658\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_1\
        );

    \I__816\ : InMux
    port map (
            O => \N__5655\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_2\
        );

    \I__815\ : InMux
    port map (
            O => \N__5652\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_3\
        );

    \I__814\ : InMux
    port map (
            O => \N__5649\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_4\
        );

    \I__813\ : InMux
    port map (
            O => \N__5646\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_5\
        );

    \I__812\ : InMux
    port map (
            O => \N__5643\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_6\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__5640\,
            I => \N__5631\
        );

    \I__810\ : InMux
    port map (
            O => \N__5639\,
            I => \N__5624\
        );

    \I__809\ : InMux
    port map (
            O => \N__5638\,
            I => \N__5624\
        );

    \I__808\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5624\
        );

    \I__807\ : InMux
    port map (
            O => \N__5636\,
            I => \N__5621\
        );

    \I__806\ : InMux
    port map (
            O => \N__5635\,
            I => \N__5618\
        );

    \I__805\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5613\
        );

    \I__804\ : InMux
    port map (
            O => \N__5631\,
            I => \N__5613\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5624\,
            I => \N__5606\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5621\,
            I => \N__5606\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5618\,
            I => \N__5606\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__5613\,
            I => \N__5600\
        );

    \I__799\ : Span4Mux_v
    port map (
            O => \N__5606\,
            I => \N__5597\
        );

    \I__798\ : InMux
    port map (
            O => \N__5605\,
            I => \N__5588\
        );

    \I__797\ : InMux
    port map (
            O => \N__5604\,
            I => \N__5583\
        );

    \I__796\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5583\
        );

    \I__795\ : Span4Mux_h
    port map (
            O => \N__5600\,
            I => \N__5578\
        );

    \I__794\ : Span4Mux_h
    port map (
            O => \N__5597\,
            I => \N__5578\
        );

    \I__793\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5575\
        );

    \I__792\ : InMux
    port map (
            O => \N__5595\,
            I => \N__5566\
        );

    \I__791\ : InMux
    port map (
            O => \N__5594\,
            I => \N__5566\
        );

    \I__790\ : InMux
    port map (
            O => \N__5593\,
            I => \N__5566\
        );

    \I__789\ : InMux
    port map (
            O => \N__5592\,
            I => \N__5566\
        );

    \I__788\ : InMux
    port map (
            O => \N__5591\,
            I => \N__5563\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5588\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5583\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__785\ : Odrv4
    port map (
            O => \N__5578\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__5575\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5566\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5563\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__781\ : InMux
    port map (
            O => \N__5550\,
            I => \N__5547\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5547\,
            I => \N__5544\
        );

    \I__779\ : Odrv12
    port map (
            O => \N__5544\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_0\
        );

    \I__778\ : CascadeMux
    port map (
            O => \N__5541\,
            I => \N__5537\
        );

    \I__777\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5531\
        );

    \I__776\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5528\
        );

    \I__775\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5525\
        );

    \I__774\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5520\
        );

    \I__773\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5520\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5531\,
            I => \N__5517\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5528\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5525\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5520\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__768\ : Odrv4
    port map (
            O => \N__5517\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__767\ : InMux
    port map (
            O => \N__5508\,
            I => \N__5505\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5505\,
            I => \N__5502\
        );

    \I__765\ : Odrv12
    port map (
            O => \N__5502\,
            I => \U712_CHIP_RAM.N_382\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__5499\,
            I => \N__5494\
        );

    \I__763\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5490\
        );

    \I__762\ : InMux
    port map (
            O => \N__5497\,
            I => \N__5487\
        );

    \I__761\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5482\
        );

    \I__760\ : InMux
    port map (
            O => \N__5493\,
            I => \N__5482\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5490\,
            I => \N__5474\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5487\,
            I => \N__5474\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__5482\,
            I => \N__5474\
        );

    \I__756\ : InMux
    port map (
            O => \N__5481\,
            I => \N__5471\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__5474\,
            I => \U712_CHIP_RAM.N_534\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5471\,
            I => \U712_CHIP_RAM.N_534\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__5466\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_cascade_\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__5463\,
            I => \U712_REG_SM.N_411_cascade_\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__5460\,
            I => \U712_BYTE_ENABLE.N_446_cascade_\
        );

    \I__750\ : IoInMux
    port map (
            O => \N__5457\,
            I => \N__5454\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__5454\,
            I => \N__5451\
        );

    \I__748\ : IoSpan4Mux
    port map (
            O => \N__5451\,
            I => \N__5448\
        );

    \I__747\ : Span4Mux_s3_v
    port map (
            O => \N__5448\,
            I => \N__5445\
        );

    \I__746\ : Sp12to4
    port map (
            O => \N__5445\,
            I => \N__5442\
        );

    \I__745\ : Span12Mux_s11_v
    port map (
            O => \N__5442\,
            I => \N__5439\
        );

    \I__744\ : Odrv12
    port map (
            O => \N__5439\,
            I => \N_52_i\
        );

    \I__743\ : InMux
    port map (
            O => \N__5436\,
            I => \N__5433\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__5433\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__5430\,
            I => \U712_CHIP_RAM.N_399_cascade_\
        );

    \I__740\ : InMux
    port map (
            O => \N__5427\,
            I => \N__5424\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5424\,
            I => \N__5420\
        );

    \I__738\ : InMux
    port map (
            O => \N__5423\,
            I => \N__5417\
        );

    \I__737\ : Span4Mux_h
    port map (
            O => \N__5420\,
            I => \N__5414\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__5417\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__5414\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__734\ : InMux
    port map (
            O => \N__5409\,
            I => \N__5406\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5406\,
            I => \N__5402\
        );

    \I__732\ : InMux
    port map (
            O => \N__5405\,
            I => \N__5399\
        );

    \I__731\ : Span4Mux_h
    port map (
            O => \N__5402\,
            I => \N__5396\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__5399\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__729\ : Odrv4
    port map (
            O => \N__5396\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__5391\,
            I => \N__5388\
        );

    \I__727\ : InMux
    port map (
            O => \N__5388\,
            I => \N__5385\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5385\,
            I => \N__5381\
        );

    \I__725\ : InMux
    port map (
            O => \N__5384\,
            I => \N__5378\
        );

    \I__724\ : Span4Mux_h
    port map (
            O => \N__5381\,
            I => \N__5375\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__5378\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__5375\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__721\ : InMux
    port map (
            O => \N__5370\,
            I => \N__5367\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5367\,
            I => \N__5363\
        );

    \I__719\ : InMux
    port map (
            O => \N__5366\,
            I => \N__5360\
        );

    \I__718\ : Span4Mux_v
    port map (
            O => \N__5363\,
            I => \N__5357\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5360\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__716\ : Odrv4
    port map (
            O => \N__5357\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__715\ : InMux
    port map (
            O => \N__5352\,
            I => \N__5349\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__5349\,
            I => \N__5346\
        );

    \I__713\ : Span4Mux_v
    port map (
            O => \N__5346\,
            I => \N__5343\
        );

    \I__712\ : Odrv4
    port map (
            O => \N__5343\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_0_3\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__5340\,
            I => \N__5337\
        );

    \I__710\ : InMux
    port map (
            O => \N__5337\,
            I => \N__5334\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__5334\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__708\ : InMux
    port map (
            O => \N__5331\,
            I => \N__5328\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__5328\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1\
        );

    \I__706\ : InMux
    port map (
            O => \N__5325\,
            I => \N__5322\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5322\,
            I => \N__5318\
        );

    \I__704\ : InMux
    port map (
            O => \N__5321\,
            I => \N__5315\
        );

    \I__703\ : Span4Mux_v
    port map (
            O => \N__5318\,
            I => \N__5312\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5315\,
            I => \N__5309\
        );

    \I__701\ : Odrv4
    port map (
            O => \N__5312\,
            I => \U712_CHIP_RAM.N_310\
        );

    \I__700\ : Odrv4
    port map (
            O => \N__5309\,
            I => \U712_CHIP_RAM.N_310\
        );

    \I__699\ : InMux
    port map (
            O => \N__5304\,
            I => \N__5301\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5301\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0\
        );

    \I__697\ : CEMux
    port map (
            O => \N__5298\,
            I => \N__5294\
        );

    \I__696\ : CEMux
    port map (
            O => \N__5297\,
            I => \N__5291\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__5294\,
            I => \N__5286\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__5291\,
            I => \N__5286\
        );

    \I__693\ : Span4Mux_v
    port map (
            O => \N__5286\,
            I => \N__5283\
        );

    \I__692\ : Odrv4
    port map (
            O => \N__5283\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__5280\,
            I => \N__5273\
        );

    \I__690\ : CascadeMux
    port map (
            O => \N__5279\,
            I => \N__5268\
        );

    \I__689\ : CascadeMux
    port map (
            O => \N__5278\,
            I => \N__5265\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__5277\,
            I => \N__5261\
        );

    \I__687\ : CascadeMux
    port map (
            O => \N__5276\,
            I => \N__5258\
        );

    \I__686\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5254\
        );

    \I__685\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5251\
        );

    \I__684\ : InMux
    port map (
            O => \N__5271\,
            I => \N__5247\
        );

    \I__683\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5242\
        );

    \I__682\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5242\
        );

    \I__681\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5239\
        );

    \I__680\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5234\
        );

    \I__679\ : InMux
    port map (
            O => \N__5258\,
            I => \N__5234\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__5257\,
            I => \N__5226\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5254\,
            I => \N__5219\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__5251\,
            I => \N__5219\
        );

    \I__675\ : InMux
    port map (
            O => \N__5250\,
            I => \N__5216\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__5247\,
            I => \N__5209\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__5242\,
            I => \N__5209\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__5239\,
            I => \N__5209\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__5234\,
            I => \N__5206\
        );

    \I__670\ : InMux
    port map (
            O => \N__5233\,
            I => \N__5201\
        );

    \I__669\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5201\
        );

    \I__668\ : InMux
    port map (
            O => \N__5231\,
            I => \N__5198\
        );

    \I__667\ : InMux
    port map (
            O => \N__5230\,
            I => \N__5195\
        );

    \I__666\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5186\
        );

    \I__665\ : InMux
    port map (
            O => \N__5226\,
            I => \N__5186\
        );

    \I__664\ : InMux
    port map (
            O => \N__5225\,
            I => \N__5186\
        );

    \I__663\ : InMux
    port map (
            O => \N__5224\,
            I => \N__5186\
        );

    \I__662\ : Odrv4
    port map (
            O => \N__5219\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5216\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__5209\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__659\ : Odrv12
    port map (
            O => \N__5206\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__5201\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__5198\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__5195\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__5186\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__654\ : InMux
    port map (
            O => \N__5169\,
            I => \N__5166\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__5166\,
            I => \N__5163\
        );

    \I__652\ : Odrv4
    port map (
            O => \N__5163\,
            I => \U712_CHIP_RAM.N_385\
        );

    \I__651\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5146\
        );

    \I__650\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5146\
        );

    \I__649\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5146\
        );

    \I__648\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5141\
        );

    \I__647\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5141\
        );

    \I__646\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5134\
        );

    \I__645\ : InMux
    port map (
            O => \N__5154\,
            I => \N__5134\
        );

    \I__644\ : InMux
    port map (
            O => \N__5153\,
            I => \N__5134\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__5146\,
            I => \U712_CHIP_RAM.N_182\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__5141\,
            I => \U712_CHIP_RAM.N_182\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__5134\,
            I => \U712_CHIP_RAM.N_182\
        );

    \I__640\ : InMux
    port map (
            O => \N__5127\,
            I => \N__5123\
        );

    \I__639\ : InMux
    port map (
            O => \N__5126\,
            I => \N__5120\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__5123\,
            I => \N__5115\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__5120\,
            I => \N__5115\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__5115\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__635\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5108\
        );

    \I__634\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5105\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__5108\,
            I => \N__5102\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__5105\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__5102\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__630\ : InMux
    port map (
            O => \N__5097\,
            I => \N__5094\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__5094\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_0_4\
        );

    \I__628\ : InMux
    port map (
            O => \N__5091\,
            I => \N__5084\
        );

    \I__627\ : InMux
    port map (
            O => \N__5090\,
            I => \N__5084\
        );

    \I__626\ : InMux
    port map (
            O => \N__5089\,
            I => \N__5081\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__5084\,
            I => \U712_CHIP_RAM.N_191\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__5081\,
            I => \U712_CHIP_RAM.N_191\
        );

    \I__623\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5072\
        );

    \I__622\ : InMux
    port map (
            O => \N__5075\,
            I => \N__5069\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__5072\,
            I => \U712_CHIP_RAM.N_327\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__5069\,
            I => \U712_CHIP_RAM.N_327\
        );

    \I__619\ : InMux
    port map (
            O => \N__5064\,
            I => \N__5059\
        );

    \I__618\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5054\
        );

    \I__617\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5054\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__5059\,
            I => \U712_CHIP_RAM.N_300\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__5054\,
            I => \U712_CHIP_RAM.N_300\
        );

    \I__614\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5046\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__5046\,
            I => \U712_CHIP_RAM.N_370\
        );

    \I__612\ : CascadeMux
    port map (
            O => \N__5043\,
            I => \N__5034\
        );

    \I__611\ : InMux
    port map (
            O => \N__5042\,
            I => \N__5031\
        );

    \I__610\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5028\
        );

    \I__609\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5025\
        );

    \I__608\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5022\
        );

    \I__607\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5017\
        );

    \I__606\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5017\
        );

    \I__605\ : InMux
    port map (
            O => \N__5034\,
            I => \N__5014\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__5031\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__5028\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5025\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__5022\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__5017\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__5014\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__5001\,
            I => \U712_CHIP_RAM.N_466_cascade_\
        );

    \I__597\ : CascadeMux
    port map (
            O => \N__4998\,
            I => \U712_CHIP_RAM.N_299_cascade_\
        );

    \I__596\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4991\
        );

    \I__595\ : InMux
    port map (
            O => \N__4994\,
            I => \N__4988\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__4991\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4988\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\
        );

    \I__592\ : InMux
    port map (
            O => \N__4983\,
            I => \N__4980\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4980\,
            I => \N__4977\
        );

    \I__590\ : Span12Mux_h
    port map (
            O => \N__4977\,
            I => \N__4974\
        );

    \I__589\ : Span12Mux_v
    port map (
            O => \N__4974\,
            I => \N__4971\
        );

    \I__588\ : Odrv12
    port map (
            O => \N__4971\,
            I => \A_c_16\
        );

    \I__587\ : InMux
    port map (
            O => \N__4968\,
            I => \N__4965\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4965\,
            I => \U712_CHIP_RAM.CMA_5_i_0_9\
        );

    \I__585\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4959\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4959\,
            I => \N__4956\
        );

    \I__583\ : Span4Mux_h
    port map (
            O => \N__4956\,
            I => \N__4953\
        );

    \I__582\ : Sp12to4
    port map (
            O => \N__4953\,
            I => \N__4950\
        );

    \I__581\ : Span12Mux_v
    port map (
            O => \N__4950\,
            I => \N__4947\
        );

    \I__580\ : Odrv12
    port map (
            O => \N__4947\,
            I => \A_c_19\
        );

    \I__579\ : IoInMux
    port map (
            O => \N__4944\,
            I => \N__4941\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4941\,
            I => \N__4938\
        );

    \I__577\ : Span12Mux_s7_h
    port map (
            O => \N__4938\,
            I => \N__4935\
        );

    \I__576\ : Span12Mux_h
    port map (
            O => \N__4935\,
            I => \N__4932\
        );

    \I__575\ : Odrv12
    port map (
            O => \N__4932\,
            I => \CMA_c_9\
        );

    \I__574\ : SRMux
    port map (
            O => \N__4929\,
            I => \N__4926\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4926\,
            I => \N__4922\
        );

    \I__572\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4919\
        );

    \I__571\ : Span4Mux_v
    port map (
            O => \N__4922\,
            I => \N__4916\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4919\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__4916\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__568\ : InMux
    port map (
            O => \N__4911\,
            I => \N__4906\
        );

    \I__567\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4903\
        );

    \I__566\ : InMux
    port map (
            O => \N__4909\,
            I => \N__4899\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__4906\,
            I => \N__4896\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4903\,
            I => \N__4893\
        );

    \I__563\ : InMux
    port map (
            O => \N__4902\,
            I => \N__4890\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4899\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__561\ : Odrv4
    port map (
            O => \N__4896\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__560\ : Odrv4
    port map (
            O => \N__4893\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4890\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__4881\,
            I => \N__4878\
        );

    \I__557\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4875\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4875\,
            I => \N__4870\
        );

    \I__555\ : InMux
    port map (
            O => \N__4874\,
            I => \N__4867\
        );

    \I__554\ : InMux
    port map (
            O => \N__4873\,
            I => \N__4863\
        );

    \I__553\ : Span4Mux_h
    port map (
            O => \N__4870\,
            I => \N__4860\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__4867\,
            I => \N__4857\
        );

    \I__551\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4854\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4863\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__549\ : Odrv4
    port map (
            O => \N__4860\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__548\ : Odrv12
    port map (
            O => \N__4857\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4854\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__546\ : InMux
    port map (
            O => \N__4845\,
            I => \N__4842\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__4842\,
            I => \N__4839\
        );

    \I__544\ : Odrv4
    port map (
            O => \N__4839\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_2\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__4836\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_\
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__4833\,
            I => \N__4830\
        );

    \I__541\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4827\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4827\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_1\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__4824\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_3_cascade_\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__4821\,
            I => \U712_CHIP_RAM.N_191_cascade_\
        );

    \I__537\ : CEMux
    port map (
            O => \N__4818\,
            I => \N__4815\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4815\,
            I => \U712_CHIP_RAM.N_191_0\
        );

    \I__535\ : InMux
    port map (
            O => \N__4812\,
            I => \N__4809\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__4809\,
            I => \N__4806\
        );

    \I__533\ : Span12Mux_h
    port map (
            O => \N__4806\,
            I => \N__4803\
        );

    \I__532\ : Span12Mux_v
    port map (
            O => \N__4803\,
            I => \N__4800\
        );

    \I__531\ : Odrv12
    port map (
            O => \N__4800\,
            I => \A_c_18\
        );

    \I__530\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4794\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__4794\,
            I => \N__4790\
        );

    \I__528\ : InMux
    port map (
            O => \N__4793\,
            I => \N__4787\
        );

    \I__527\ : Odrv4
    port map (
            O => \N__4790\,
            I => \U712_CHIP_RAM.N_315\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4787\,
            I => \U712_CHIP_RAM.N_315\
        );

    \I__525\ : CascadeMux
    port map (
            O => \N__4782\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_\
        );

    \I__524\ : InMux
    port map (
            O => \N__4779\,
            I => \N__4776\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4776\,
            I => \U712_CHIP_RAM.N_336\
        );

    \I__522\ : InMux
    port map (
            O => \N__4773\,
            I => \N__4770\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4770\,
            I => \N__4767\
        );

    \I__520\ : Odrv4
    port map (
            O => \N__4767\,
            I => \U712_CHIP_RAM.N_372\
        );

    \I__519\ : IoInMux
    port map (
            O => \N__4764\,
            I => \N__4761\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4761\,
            I => \N__4758\
        );

    \I__517\ : IoSpan4Mux
    port map (
            O => \N__4758\,
            I => \N__4755\
        );

    \I__516\ : Span4Mux_s0_h
    port map (
            O => \N__4755\,
            I => \N__4752\
        );

    \I__515\ : Sp12to4
    port map (
            O => \N__4752\,
            I => \N__4749\
        );

    \I__514\ : Span12Mux_h
    port map (
            O => \N__4749\,
            I => \N__4746\
        );

    \I__513\ : Span12Mux_v
    port map (
            O => \N__4746\,
            I => \N__4743\
        );

    \I__512\ : Odrv12
    port map (
            O => \N__4743\,
            I => \CMA_c_8\
        );

    \I__511\ : InMux
    port map (
            O => \N__4740\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__510\ : InMux
    port map (
            O => \N__4737\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__509\ : InMux
    port map (
            O => \N__4734\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__508\ : CascadeMux
    port map (
            O => \N__4731\,
            I => \N__4728\
        );

    \I__507\ : InMux
    port map (
            O => \N__4728\,
            I => \N__4724\
        );

    \I__506\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4719\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4724\,
            I => \N__4716\
        );

    \I__504\ : InMux
    port map (
            O => \N__4723\,
            I => \N__4711\
        );

    \I__503\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4711\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4719\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__501\ : Odrv4
    port map (
            O => \N__4716\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4711\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__499\ : InMux
    port map (
            O => \N__4704\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__498\ : InMux
    port map (
            O => \N__4701\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__497\ : InMux
    port map (
            O => \N__4698\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__496\ : InMux
    port map (
            O => \N__4695\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__495\ : InMux
    port map (
            O => \N__4692\,
            I => \N__4687\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__4691\,
            I => \N__4683\
        );

    \I__493\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4680\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__4687\,
            I => \N__4677\
        );

    \I__491\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4672\
        );

    \I__490\ : InMux
    port map (
            O => \N__4683\,
            I => \N__4672\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4680\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__488\ : Odrv12
    port map (
            O => \N__4677\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4672\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__486\ : InMux
    port map (
            O => \N__4665\,
            I => \N__4662\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__4662\,
            I => \U712_CHIP_RAM.LATCH_CLK_6\
        );

    \I__484\ : CascadeMux
    port map (
            O => \N__4659\,
            I => \U712_CHIP_RAM.N_396_cascade_\
        );

    \I__483\ : IoInMux
    port map (
            O => \N__4656\,
            I => \N__4653\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4653\,
            I => \N__4650\
        );

    \I__481\ : Span12Mux_s1_v
    port map (
            O => \N__4650\,
            I => \N__4647\
        );

    \I__480\ : Span12Mux_v
    port map (
            O => \N__4647\,
            I => \N__4643\
        );

    \I__479\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4640\
        );

    \I__478\ : Odrv12
    port map (
            O => \N__4643\,
            I => \LATCH_CLK_c\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4640\,
            I => \LATCH_CLK_c\
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__4635\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_2_0_cascade_\
        );

    \I__475\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4629\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4629\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_2_3\
        );

    \I__473\ : CascadeMux
    port map (
            O => \N__4626\,
            I => \U712_CHIP_RAM.N_301_cascade_\
        );

    \I__472\ : CascadeMux
    port map (
            O => \N__4623\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_0_1_cascade_\
        );

    \I__471\ : CascadeMux
    port map (
            O => \N__4620\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_1_5_cascade_\
        );

    \I__470\ : InMux
    port map (
            O => \N__4617\,
            I => \N__4614\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4614\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_1_4\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__4611\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_2_2_cascade_\
        );

    \I__467\ : InMux
    port map (
            O => \N__4608\,
            I => \N__4602\
        );

    \I__466\ : InMux
    port map (
            O => \N__4607\,
            I => \N__4602\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4602\,
            I => \U712_CHIP_RAM.N_433\
        );

    \I__464\ : CascadeMux
    port map (
            O => \N__4599\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_4_i_2_cascade_\
        );

    \I__463\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4593\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4593\,
            I => \N__4590\
        );

    \I__461\ : Odrv4
    port map (
            O => \N__4590\,
            I => \U712_CHIP_RAM.N_65\
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__4587\,
            I => \U712_CHIP_RAM.N_173_cascade_\
        );

    \I__459\ : IoInMux
    port map (
            O => \N__4584\,
            I => \N__4581\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4581\,
            I => \N__4578\
        );

    \I__457\ : Span12Mux_s8_v
    port map (
            O => \N__4578\,
            I => \N__4575\
        );

    \I__456\ : Odrv12
    port map (
            O => \N__4575\,
            I => \VBENn_c\
        );

    \I__455\ : InMux
    port map (
            O => \N__4572\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__454\ : InMux
    port map (
            O => \N__4569\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__453\ : InMux
    port map (
            O => \N__4566\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__452\ : ClkMux
    port map (
            O => \N__4563\,
            I => \N__4539\
        );

    \I__451\ : ClkMux
    port map (
            O => \N__4562\,
            I => \N__4539\
        );

    \I__450\ : ClkMux
    port map (
            O => \N__4561\,
            I => \N__4539\
        );

    \I__449\ : ClkMux
    port map (
            O => \N__4560\,
            I => \N__4539\
        );

    \I__448\ : ClkMux
    port map (
            O => \N__4559\,
            I => \N__4539\
        );

    \I__447\ : ClkMux
    port map (
            O => \N__4558\,
            I => \N__4539\
        );

    \I__446\ : ClkMux
    port map (
            O => \N__4557\,
            I => \N__4539\
        );

    \I__445\ : ClkMux
    port map (
            O => \N__4556\,
            I => \N__4539\
        );

    \I__444\ : GlobalMux
    port map (
            O => \N__4539\,
            I => \N__4536\
        );

    \I__443\ : gio2CtrlBuf
    port map (
            O => \N__4536\,
            I => \C1_c_g\
        );

    \I__442\ : InMux
    port map (
            O => \N__4533\,
            I => \N__4529\
        );

    \I__441\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4526\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4529\,
            I => \N__4523\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4526\,
            I => \N__4520\
        );

    \I__438\ : Span4Mux_v
    port map (
            O => \N__4523\,
            I => \N__4517\
        );

    \I__437\ : Span4Mux_v
    port map (
            O => \N__4520\,
            I => \N__4514\
        );

    \I__436\ : Span4Mux_h
    port map (
            O => \N__4517\,
            I => \N__4511\
        );

    \I__435\ : Sp12to4
    port map (
            O => \N__4514\,
            I => \N__4508\
        );

    \I__434\ : Sp12to4
    port map (
            O => \N__4511\,
            I => \N__4503\
        );

    \I__433\ : Span12Mux_h
    port map (
            O => \N__4508\,
            I => \N__4503\
        );

    \I__432\ : Odrv12
    port map (
            O => \N__4503\,
            I => \DBRn_c\
        );

    \I__431\ : InMux
    port map (
            O => \N__4500\,
            I => \N__4497\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__4497\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__429\ : InMux
    port map (
            O => \N__4494\,
            I => \N__4491\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__4491\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_1_1\
        );

    \I__427\ : CascadeMux
    port map (
            O => \N__4488\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_1_0_cascade_\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__4485\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1_cascade_\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__4482\,
            I => \U712_CHIP_RAM.N_442_cascade_\
        );

    \I__424\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4473\
        );

    \I__423\ : InMux
    port map (
            O => \N__4478\,
            I => \N__4473\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4473\,
            I => \U712_CHIP_RAM.CLK_EN_5_0\
        );

    \I__421\ : InMux
    port map (
            O => \N__4470\,
            I => \N__4467\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__4467\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__419\ : InMux
    port map (
            O => \N__4464\,
            I => \bfn_7_13_0_\
        );

    \I__418\ : InMux
    port map (
            O => \N__4461\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__417\ : InMux
    port map (
            O => \N__4458\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__416\ : InMux
    port map (
            O => \N__4455\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__415\ : InMux
    port map (
            O => \N__4452\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__4449\,
            I => \N__4446\
        );

    \I__413\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4443\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__4443\,
            I => \N__4439\
        );

    \I__411\ : InMux
    port map (
            O => \N__4442\,
            I => \N__4436\
        );

    \I__410\ : Span4Mux_h
    port map (
            O => \N__4439\,
            I => \N__4433\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__4436\,
            I => \N__4430\
        );

    \I__408\ : Span4Mux_v
    port map (
            O => \N__4433\,
            I => \N__4427\
        );

    \I__407\ : Span4Mux_h
    port map (
            O => \N__4430\,
            I => \N__4424\
        );

    \I__406\ : Odrv4
    port map (
            O => \N__4427\,
            I => \DBRn_c_i\
        );

    \I__405\ : Odrv4
    port map (
            O => \N__4424\,
            I => \DBRn_c_i\
        );

    \I__404\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4416\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__4416\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\
        );

    \I__402\ : CascadeMux
    port map (
            O => \N__4413\,
            I => \U712_CHIP_RAM.N_458_cascade_\
        );

    \I__401\ : CascadeMux
    port map (
            O => \N__4410\,
            I => \N__4407\
        );

    \I__400\ : InMux
    port map (
            O => \N__4407\,
            I => \N__4401\
        );

    \I__399\ : InMux
    port map (
            O => \N__4406\,
            I => \N__4401\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__4401\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\
        );

    \I__397\ : CascadeMux
    port map (
            O => \N__4398\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a2_0_cascade_\
        );

    \I__396\ : IoInMux
    port map (
            O => \N__4395\,
            I => \N__4392\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4392\,
            I => \N__4389\
        );

    \I__394\ : Span12Mux_s2_h
    port map (
            O => \N__4389\,
            I => \N__4386\
        );

    \I__393\ : Span12Mux_h
    port map (
            O => \N__4386\,
            I => \N__4383\
        );

    \I__392\ : Span12Mux_v
    port map (
            O => \N__4383\,
            I => \N__4379\
        );

    \I__391\ : InMux
    port map (
            O => \N__4382\,
            I => \N__4376\
        );

    \I__390\ : Odrv12
    port map (
            O => \N__4379\,
            I => \CLK_EN_c\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__4376\,
            I => \CLK_EN_c\
        );

    \I__388\ : IoInMux
    port map (
            O => \N__4371\,
            I => \N__4368\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__4368\,
            I => \N__4365\
        );

    \I__386\ : Odrv12
    port map (
            O => \N__4365\,
            I => \DBRn_c_i_0\
        );

    \I__385\ : IoInMux
    port map (
            O => \N__4362\,
            I => \N__4359\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__4359\,
            I => \N__4356\
        );

    \I__383\ : Span4Mux_s3_v
    port map (
            O => \N__4356\,
            I => \N__4353\
        );

    \I__382\ : Span4Mux_h
    port map (
            O => \N__4353\,
            I => \N__4350\
        );

    \I__381\ : Odrv4
    port map (
            O => \N__4350\,
            I => \CLK80_PLL_i_i\
        );

    \I__380\ : IoInMux
    port map (
            O => \N__4347\,
            I => \N__4344\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__378\ : IoSpan4Mux
    port map (
            O => \N__4341\,
            I => \N__4338\
        );

    \I__377\ : Span4Mux_s2_v
    port map (
            O => \N__4338\,
            I => \N__4335\
        );

    \I__376\ : Sp12to4
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__375\ : Span12Mux_v
    port map (
            O => \N__4332\,
            I => \N__4329\
        );

    \I__374\ : Odrv12
    port map (
            O => \N__4329\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__4559\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__4561\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__4562\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__4557\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__4556\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__4558\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            I => \N__4563\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_12_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7796\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9483\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4371\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8496\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__4442\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11220\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_3_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10770\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4533\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__10152\,
            in1 => \N__11552\,
            in2 => \N__4449\,
            in3 => \N__5738\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            ce => 'H',
            sr => \N__11195\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010001000"
        )
    port map (
            in0 => \N__5272\,
            in1 => \N__7754\,
            in2 => \N__6420\,
            in3 => \N__7598\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_5_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__10958\,
            in1 => \_gnd_net_\,
            in2 => \N__4410\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10753\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6081\,
            in1 => \N__4419\,
            in2 => \_gnd_net_\,
            in3 => \N__4406\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_458_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__10956\,
            in1 => \N__8708\,
            in2 => \N__4413\,
            in3 => \N__7425\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10753\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_4_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10957\,
            in2 => \_gnd_net_\,
            in3 => \N__8625\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10753\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7740\,
            in1 => \N__7599\,
            in2 => \N__6418\,
            in3 => \N__5604\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000110011011100"
        )
    port map (
            in0 => \N__5038\,
            in1 => \N__4382\,
            in2 => \N__4398\,
            in3 => \N__4479\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10758\,
            ce => 'H',
            sr => \N__11173\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIN5DI_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5232\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5536\,
            lcout => \U712_CHIP_RAM.CLK_EN_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8934\,
            in1 => \N__7739\,
            in2 => \_gnd_net_\,
            in3 => \N__5233\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4793\,
            in1 => \N__5603\,
            in2 => \N__4485\,
            in3 => \N__5037\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_442_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__8935\,
            in1 => \_gnd_net_\,
            in2 => \N__4482\,
            in3 => \N__4478\,
            lcout => \U712_CHIP_RAM.N_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__8936\,
            in1 => \N__7011\,
            in2 => \_gnd_net_\,
            in3 => \N__6219\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10758\,
            ce => 'H',
            sr => \N__11173\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4470\,
            in2 => \_gnd_net_\,
            in3 => \N__4464\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__4560\,
            ce => 'H',
            sr => \N__4929\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5366\,
            in2 => \_gnd_net_\,
            in3 => \N__4461\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__4560\,
            ce => 'H',
            sr => \N__4929\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5405\,
            in2 => \_gnd_net_\,
            in3 => \N__4458\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__4560\,
            ce => 'H',
            sr => \N__4929\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5423\,
            in2 => \_gnd_net_\,
            in3 => \N__4455\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__4560\,
            ce => 'H',
            sr => \N__4929\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5384\,
            in2 => \_gnd_net_\,
            in3 => \N__4452\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__4560\,
            ce => 'H',
            sr => \N__4929\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5111\,
            in2 => \_gnd_net_\,
            in3 => \N__4572\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__4560\,
            ce => 'H',
            sr => \N__4929\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5127\,
            in2 => \_gnd_net_\,
            in3 => \N__4569\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__4560\,
            ce => 'H',
            sr => \N__4929\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6269\,
            in2 => \_gnd_net_\,
            in3 => \N__4566\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4560\,
            ce => 'H',
            sr => \N__4929\
        );

    \DBR_SYNC_0_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4532\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10765\,
            ce => 'H',
            sr => \N__11160\
        );

    \DBR_SYNC_1_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4500\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10765\,
            ce => 'H',
            sr => \N__11160\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNIK9021_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__10071\,
            in1 => \N__7996\,
            in2 => \N__9409\,
            in3 => \N__10017\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_2_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__5264\,
            in1 => \N__4692\,
            in2 => \N__5640\,
            in3 => \N__4874\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__6419\,
            in1 => \N__4910\,
            in2 => \N__4731\,
            in3 => \N__5634\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMDsr_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__4608\,
            in1 => \N__4494\,
            in2 => \N__4488\,
            in3 => \N__5325\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMDsr_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__8011\,
            in1 => \N__5090\,
            in2 => \N__4620\,
            in3 => \N__4617\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10738\,
            ce => 'H',
            sr => \N__11188\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__7595\,
            in1 => \N__4607\,
            in2 => \N__5280\,
            in3 => \N__7753\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMDsr_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__5091\,
            in1 => \N__4632\,
            in2 => \N__4611\,
            in3 => \N__10078\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10738\,
            ce => 'H',
            sr => \N__11188\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5637\,
            in1 => \N__7745\,
            in2 => \N__5278\,
            in3 => \N__7592\,
            lcout => \U712_CHIP_RAM.N_433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110110011101"
        )
    port map (
            in0 => \N__5639\,
            in1 => \N__7746\,
            in2 => \N__5279\,
            in3 => \N__6312\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_4_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__7594\,
            in1 => \N__5042\,
            in2 => \N__4599\,
            in3 => \N__5064\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_173_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__4596\,
            in1 => \N__11010\,
            in2 => \N__4587\,
            in3 => \N__8803\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10743\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__9025\,
            in1 => \N__7956\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__5638\,
            in1 => \N__7744\,
            in2 => \_gnd_net_\,
            in3 => \N__5040\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMDsr_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110111"
        )
    port map (
            in0 => \N__7593\,
            in1 => \N__5169\,
            in2 => \N__4635\,
            in3 => \N__5321\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNILL5O1_0_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__6378\,
            in1 => \N__7590\,
            in2 => \N__5257\,
            in3 => \N__7697\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIC9HD1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__5593\,
            in1 => \N__7691\,
            in2 => \_gnd_net_\,
            in3 => \N__7408\,
            lcout => \U712_CHIP_RAM.N_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4866\,
            in1 => \N__4902\,
            in2 => \N__4691\,
            in3 => \N__4722\,
            lcout => \U712_CHIP_RAM.N_301\,
            ltout => \U712_CHIP_RAM.N_301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__5592\,
            in1 => \_gnd_net_\,
            in2 => \N__4626\,
            in3 => \N__5224\,
            lcout => \U712_CHIP_RAM.N_534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4686\,
            in1 => \N__4723\,
            in2 => \_gnd_net_\,
            in3 => \N__5594\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__5595\,
            in1 => \N__5229\,
            in2 => \_gnd_net_\,
            in3 => \N__5039\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMDsr_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__4773\,
            in1 => \N__7591\,
            in2 => \N__4623\,
            in3 => \N__5076\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5225\,
            in2 => \_gnd_net_\,
            in3 => \N__6377\,
            lcout => \U712_CHIP_RAM.N_300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6397\,
            in2 => \_gnd_net_\,
            in3 => \N__8720\,
            lcout => \U712_CHIP_RAM.LATCH_CLK_6\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5158\,
            in1 => \N__5250\,
            in2 => \_gnd_net_\,
            in3 => \N__4740\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__10754\,
            ce => \N__5297\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7730\,
            in2 => \_gnd_net_\,
            in3 => \N__4737\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5159\,
            in1 => \N__5605\,
            in2 => \_gnd_net_\,
            in3 => \N__4734\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__10754\,
            ce => \N__5297\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5153\,
            in1 => \N__4727\,
            in2 => \_gnd_net_\,
            in3 => \N__4704\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__10754\,
            ce => \N__5297\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5160\,
            in1 => \N__4909\,
            in2 => \_gnd_net_\,
            in3 => \N__4701\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__10754\,
            ce => \N__5297\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5154\,
            in1 => \N__4873\,
            in2 => \_gnd_net_\,
            in3 => \N__4698\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__10754\,
            ce => \N__5297\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__4690\,
            in1 => \N__5155\,
            in2 => \_gnd_net_\,
            in3 => \N__4695\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10754\,
            ce => \N__5297\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4797\,
            in1 => \N__5498\,
            in2 => \N__7738\,
            in3 => \N__7545\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_396_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__11006\,
            in1 => \N__4665\,
            in2 => \N__4659\,
            in3 => \N__4646\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5534\,
            in2 => \_gnd_net_\,
            in3 => \N__6379\,
            lcout => \U712_CHIP_RAM.N_315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__6154\,
            in1 => \N__10556\,
            in2 => \_gnd_net_\,
            in3 => \N__7439\,
            lcout => \U712_CHIP_RAM.N_336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIU7TF5_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__7438\,
            in1 => \N__6099\,
            in2 => \N__6456\,
            in3 => \N__5979\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__5535\,
            in1 => \N__11007\,
            in2 => \N__4782\,
            in3 => \N__4779\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100110101011"
        )
    port map (
            in0 => \N__6383\,
            in1 => \N__5231\,
            in2 => \N__7583\,
            in3 => \N__7698\,
            lcout => \U712_CHIP_RAM.N_372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11008\,
            in2 => \_gnd_net_\,
            in3 => \N__5436\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10762\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__11009\,
            in1 => \N__6067\,
            in2 => \_gnd_net_\,
            in3 => \N__7215\,
            lcout => \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__8012\,
            in1 => \N__9406\,
            in2 => \_gnd_net_\,
            in3 => \N__10028\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8389\,
            in1 => \N__8037\,
            in2 => \N__6900\,
            in3 => \N__5724\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10731\,
            ce => \N__8293\,
            sr => \N__11189\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__4968\,
            in1 => \N__4962\,
            in2 => \N__9056\,
            in3 => \N__8028\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10731\,
            ce => \N__8293\,
            sr => \N__11189\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIDBLK1_3_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__7997\,
            in1 => \N__4925\,
            in2 => \N__9410\,
            in3 => \N__10072\,
            lcout => \U712_CHIP_RAM.un1_CMA25_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7742\,
            in2 => \_gnd_net_\,
            in3 => \N__7379\,
            lcout => \U712_CHIP_RAM.DBENn_7_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_0_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__5508\,
            in1 => \N__4911\,
            in2 => \N__4881\,
            in3 => \N__4845\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111001011111010"
        )
    port map (
            in0 => \N__7596\,
            in1 => \N__7743\,
            in2 => \N__4836\,
            in3 => \N__5271\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10734\,
            ce => \N__4818\,
            sr => \N__11184\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI1DB24_2_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__6182\,
            in1 => \N__7741\,
            in2 => \N__4833\,
            in3 => \N__5063\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI2MHHA_2_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__5550\,
            in1 => \N__5049\,
            in2 => \N__4824\,
            in3 => \N__5041\,
            lcout => \U712_CHIP_RAM.N_191\,
            ltout => \U712_CHIP_RAM.N_191_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_0_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11219\,
            in1 => \_gnd_net_\,
            in2 => \N__4821\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_191_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4812\,
            in1 => \N__4995\,
            in2 => \_gnd_net_\,
            in3 => \N__7003\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10739\,
            ce => 'H',
            sr => \N__11174\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__5097\,
            in1 => \N__5089\,
            in2 => \N__9408\,
            in3 => \N__5352\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10739\,
            ce => 'H',
            sr => \N__11174\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI7FAQ2_3_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__5635\,
            in1 => \N__5075\,
            in2 => \_gnd_net_\,
            in3 => \N__5062\,
            lcout => \U712_CHIP_RAM.N_370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__6183\,
            in1 => \N__10954\,
            in2 => \N__7443\,
            in3 => \N__5978\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5591\,
            in1 => \N__6375\,
            in2 => \N__5043\,
            in3 => \N__5230\,
            lcout => \U712_CHIP_RAM.N_466\,
            ltout => \U712_CHIP_RAM.N_466_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__7692\,
            in1 => \_gnd_net_\,
            in2 => \N__5001\,
            in3 => \N__7578\,
            lcout => \U712_CHIP_RAM.N_471\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5540\,
            in2 => \_gnd_net_\,
            in3 => \N__6376\,
            lcout => \U712_CHIP_RAM.N_299\,
            ltout => \U712_CHIP_RAM.N_299_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7693\,
            in1 => \N__7579\,
            in2 => \N__4998\,
            in3 => \N__5481\,
            lcout => \U712_CHIP_RAM.N_429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4994\,
            in1 => \N__4983\,
            in2 => \_gnd_net_\,
            in3 => \N__9356\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7694\,
            in1 => \N__7580\,
            in2 => \_gnd_net_\,
            in3 => \N__7371\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__10955\,
            in1 => \N__5497\,
            in2 => \N__5430\,
            in3 => \N__6300\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__5427\,
            in1 => \N__5409\,
            in2 => \N__5391\,
            in3 => \N__5370\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011000100"
        )
    port map (
            in0 => \N__6243\,
            in1 => \N__7547\,
            in2 => \N__5277\,
            in3 => \N__7708\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__11000\,
            in1 => \N__5156\,
            in2 => \N__5340\,
            in3 => \N__5331\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10748\,
            ce => \N__5298\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7707\,
            in2 => \_gnd_net_\,
            in3 => \N__6385\,
            lcout => \U712_CHIP_RAM.N_310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001011011110"
        )
    port map (
            in0 => \N__5870\,
            in1 => \N__5157\,
            in2 => \N__6404\,
            in3 => \N__5304\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10748\,
            ce => \N__5298\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111111101"
        )
    port map (
            in0 => \N__5636\,
            in1 => \N__6384\,
            in2 => \N__5276\,
            in3 => \N__7546\,
            lcout => \U712_CHIP_RAM.N_385\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__11002\,
            in1 => \N__6279\,
            in2 => \N__6296\,
            in3 => \N__5493\,
            lcout => \U712_CHIP_RAM.N_182\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5126\,
            in2 => \_gnd_net_\,
            in3 => \N__5112\,
            lcout => \U712_CHIP_RAM.REFRESH5lto7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010101010101"
        )
    port map (
            in0 => \N__11003\,
            in1 => \N__5596\,
            in2 => \N__7582\,
            in3 => \N__7695\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_0_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010110001"
        )
    port map (
            in0 => \N__7540\,
            in1 => \N__7696\,
            in2 => \N__5541\,
            in3 => \N__6389\,
            lcout => \U712_CHIP_RAM.N_382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6390\,
            in1 => \N__7541\,
            in2 => \N__5499\,
            in3 => \N__7737\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11001\,
            in2 => \N__5466\,
            in3 => \N__7556\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10755\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__7905\,
            in1 => \N__7191\,
            in2 => \N__9210\,
            in3 => \N__7236\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__11005\,
            in1 => \N__9209\,
            in2 => \N__5463\,
            in3 => \N__9621\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__11872\,
            in1 => \N__8766\,
            in2 => \_gnd_net_\,
            in3 => \N__8724\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_52_i_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__7146\,
            in1 => \N__7158\,
            in2 => \N__5460\,
            in3 => \N__9800\,
            lcout => \N_52_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__11004\,
            in1 => \N__11873\,
            in2 => \_gnd_net_\,
            in3 => \N__11927\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6513\,
            in2 => \N__6558\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBR_COUNT_2_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6527\,
            in2 => \_gnd_net_\,
            in3 => \N__5658\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_1\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_2\,
            clk => \N__10763\,
            ce => 'H',
            sr => \N__5888\
        );

    \U712_CHIP_RAM.DBR_COUNT_3_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6791\,
            in2 => \_gnd_net_\,
            in3 => \N__5655\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_2\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_3\,
            clk => \N__10763\,
            ce => 'H',
            sr => \N__5888\
        );

    \U712_CHIP_RAM.DBR_COUNT_4_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6804\,
            in2 => \_gnd_net_\,
            in3 => \N__5652\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_3\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_4\,
            clk => \N__10763\,
            ce => 'H',
            sr => \N__5888\
        );

    \U712_CHIP_RAM.DBR_COUNT_5_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6816\,
            in2 => \_gnd_net_\,
            in3 => \N__5649\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_4\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_5\,
            clk => \N__10763\,
            ce => 'H',
            sr => \N__5888\
        );

    \U712_CHIP_RAM.DBR_COUNT_6_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6540\,
            in2 => \_gnd_net_\,
            in3 => \N__5646\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_5\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_6\,
            clk => \N__10763\,
            ce => 'H',
            sr => \N__5888\
        );

    \U712_CHIP_RAM.DBR_COUNT_7_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6777\,
            in2 => \_gnd_net_\,
            in3 => \N__5643\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10763\,
            ce => 'H',
            sr => \N__5888\
        );

    \U712_CHIP_RAM.DBR_COUNT_1_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__6514\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6557\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10763\,
            ce => 'H',
            sr => \N__5888\
        );

    \U712_CHIP_RAM.DBR_COUNT_0_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6516\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10766\,
            ce => 'H',
            sr => \N__5889\
        );

    \CONSTANT_ONE_LUT4_LC_10_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__5703\,
            in1 => \N__8390\,
            in2 => \N__9447\,
            in3 => \N__6171\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10722\,
            ce => \N__8290\,
            sr => \N__11190\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5804\,
            in1 => \N__5924\,
            in2 => \_gnd_net_\,
            in3 => \N__9439\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9440\,
            in1 => \N__9038\,
            in2 => \N__5769\,
            in3 => \N__9267\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9438\,
            in1 => \N__5678\,
            in2 => \_gnd_net_\,
            in3 => \N__5766\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9037\,
            in1 => \N__9441\,
            in2 => \N__5742\,
            in3 => \N__5739\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5718\,
            in1 => \N__9036\,
            in2 => \_gnd_net_\,
            in3 => \N__9960\,
            lcout => \U712_CHIP_RAM.N_353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__5697\,
            in1 => \N__11531\,
            in2 => \N__5682\,
            in3 => \N__7007\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10732\,
            ce => 'H',
            sr => \N__11175\
        );

    \U712_CHIP_RAM.DBENn_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011101110"
        )
    port map (
            in0 => \N__8745\,
            in1 => \N__6201\,
            in2 => \N__5667\,
            in3 => \N__9969\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10732\,
            ce => 'H',
            sr => \N__11175\
        );

    \U712_CHIP_RAM.DBDIR_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__6162\,
            in1 => \N__6038\,
            in2 => \_gnd_net_\,
            in3 => \N__6114\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10732\,
            ce => 'H',
            sr => \N__11175\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI3LH42_3_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11218\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6027\,
            lcout => \U712_CHIP_RAM.un1_CMA25_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6021\,
            in1 => \N__5987\,
            in2 => \_gnd_net_\,
            in3 => \N__9344\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5988\,
            in1 => \N__6006\,
            in2 => \_gnd_net_\,
            in3 => \N__7001\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10735\,
            ce => 'H',
            sr => \N__11168\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIU7TF5_0_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6449\,
            in1 => \N__6092\,
            in2 => \N__7450\,
            in3 => \N__5974\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5958\,
            in2 => \N__5943\,
            in3 => \N__8162\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10735\,
            ce => 'H',
            sr => \N__11168\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5925\,
            in1 => \N__5940\,
            in2 => \_gnd_net_\,
            in3 => \N__7000\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10735\,
            ce => 'H',
            sr => \N__11168\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7002\,
            in1 => \N__5907\,
            in2 => \_gnd_net_\,
            in3 => \N__8123\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10735\,
            ce => 'H',
            sr => \N__11168\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7719\,
            in1 => \N__7367\,
            in2 => \N__7451\,
            in3 => \N__7581\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6222\,
            in3 => \N__6215\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6192\,
            in3 => \N__11217\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9004\,
            in1 => \N__6189\,
            in2 => \N__9407\,
            in3 => \N__10101\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__6241\,
            in1 => \N__6571\,
            in2 => \_gnd_net_\,
            in3 => \N__6441\,
            lcout => \U712_CHIP_RAM.N_319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9003\,
            in1 => \N__7074\,
            in2 => \_gnd_net_\,
            in3 => \N__9930\,
            lcout => \U712_CHIP_RAM.N_359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011000000"
        )
    port map (
            in0 => \N__6161\,
            in1 => \N__10600\,
            in2 => \N__10877\,
            in3 => \N__6113\,
            lcout => \DMA_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10740\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIFGNH_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6572\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6242\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__7241\,
            in1 => \N__10943\,
            in2 => \N__6492\,
            in3 => \N__6080\,
            lcout => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10744\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8990\,
            in2 => \_gnd_net_\,
            in3 => \N__6448\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_419_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__7313\,
            in1 => \N__10942\,
            in2 => \N__6477\,
            in3 => \N__6474\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10744\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010000100000"
        )
    port map (
            in0 => \N__7709\,
            in1 => \N__7548\,
            in2 => \N__6414\,
            in3 => \N__6311\,
            lcout => \U712_CHIP_RAM.N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__7549\,
            in1 => \N__7710\,
            in2 => \_gnd_net_\,
            in3 => \N__7378\,
            lcout => \U712_CHIP_RAM.N_434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__6273\,
            in1 => \N__6255\,
            in2 => \N__10996\,
            in3 => \N__6249\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10744\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7182\,
            in2 => \_gnd_net_\,
            in3 => \N__9139\,
            lcout => \U712_REG_SM.N_322\,
            ltout => \U712_REG_SM.N_322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9237\,
            in1 => \N__7277\,
            in2 => \N__6228\,
            in3 => \N__7903\,
            lcout => \U712_REG_SM.N_410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__9605\,
            in1 => \N__9236\,
            in2 => \_gnd_net_\,
            in3 => \N__9198\,
            lcout => \U712_REG_SM.N_367\,
            ltout => \U712_REG_SM.N_367_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6644\,
            in2 => \N__6225\,
            in3 => \N__7904\,
            lcout => \U712_REG_SM.N_131\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_RNO_0_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000100010"
        )
    port map (
            in0 => \N__9199\,
            in1 => \N__7278\,
            in2 => \N__9147\,
            in3 => \N__6610\,
            lcout => \U712_REG_SM.REGENn_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9606\,
            in1 => \N__7183\,
            in2 => \N__7242\,
            in3 => \N__9200\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_408_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011100100"
        )
    port map (
            in0 => \N__10948\,
            in1 => \N__7948\,
            in2 => \N__6660\,
            in3 => \N__6657\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10749\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001101"
        )
    port map (
            in0 => \N__6594\,
            in1 => \N__6651\,
            in2 => \N__7911\,
            in3 => \N__7965\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10756\,
            ce => 'H',
            sr => \N__11156\
        );

    \U712_REG_SM.WRITE_CYCLE_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__10579\,
            in1 => \N__6645\,
            in2 => \_gnd_net_\,
            in3 => \N__8446\,
            lcout => \U712_REG_SM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10756\,
            ce => 'H',
            sr => \N__11156\
        );

    \U712_REG_SM.REGENn_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010011010100010"
        )
    port map (
            in0 => \N__6611\,
            in1 => \N__6633\,
            in2 => \N__9618\,
            in3 => \N__7254\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10756\,
            ce => 'H',
            sr => \N__11156\
        );

    \U712_REG_SM.REG_TACK_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__6593\,
            in1 => \N__7875\,
            in2 => \N__8847\,
            in3 => \N__6585\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10756\,
            ce => 'H',
            sr => \N__11156\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6579\,
            in1 => \N__6553\,
            in2 => \_gnd_net_\,
            in3 => \N__6539\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_5_i_a2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6528\,
            in1 => \N__6515\,
            in2 => \N__6495\,
            in3 => \N__6765\,
            lcout => \U712_CHIP_RAM.N_456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__10463\,
            in1 => \N__9868\,
            in2 => \_gnd_net_\,
            in3 => \N__9011\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6815\,
            in1 => \N__6803\,
            in2 => \N__6792\,
            in3 => \N__6776\,
            lcout => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_5_i_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__9012\,
            in1 => \N__10464\,
            in2 => \_gnd_net_\,
            in3 => \N__10421\,
            lcout => \U712_BYTE_ENABLE.N_424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9835\,
            in1 => \N__10405\,
            in2 => \N__10575\,
            in3 => \N__10500\,
            lcout => \U712_REG_SM.N_402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__11868\,
            in1 => \N__11919\,
            in2 => \_gnd_net_\,
            in3 => \N__10619\,
            lcout => \DMA_LATCH_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__8391\,
            in1 => \N__10092\,
            in2 => \_gnd_net_\,
            in3 => \N__9417\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10720\,
            ce => \N__8292\,
            sr => \N__11185\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6719\,
            in1 => \N__7044\,
            in2 => \_gnd_net_\,
            in3 => \N__9419\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9035\,
            in1 => \N__9442\,
            in2 => \N__6684\,
            in3 => \N__9981\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__6879\,
            in1 => \N__8377\,
            in2 => \N__6681\,
            in3 => \N__11298\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10723\,
            ce => \N__8300\,
            sr => \N__11176\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9034\,
            in2 => \_gnd_net_\,
            in3 => \N__9418\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__10314\,
            in1 => \N__8378\,
            in2 => \N__6894\,
            in3 => \N__7110\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10723\,
            ce => \N__8300\,
            sr => \N__11176\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7005\,
            in1 => \N__7092\,
            in2 => \_gnd_net_\,
            in3 => \N__7073\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10728\,
            ce => 'H',
            sr => \N__11169\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7059\,
            in1 => \N__7043\,
            in2 => \_gnd_net_\,
            in3 => \N__7004\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10728\,
            ce => 'H',
            sr => \N__11169\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7029\,
            in1 => \N__8226\,
            in2 => \_gnd_net_\,
            in3 => \N__7006\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10728\,
            ce => 'H',
            sr => \N__11169\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__8375\,
            in1 => \N__6892\,
            in2 => \N__10254\,
            in3 => \N__8106\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10733\,
            ce => \N__8301\,
            sr => \N__11161\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8373\,
            in1 => \N__9255\,
            in2 => \N__6898\,
            in3 => \N__8631\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10733\,
            ce => \N__8301\,
            sr => \N__11161\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__8376\,
            in1 => \N__6893\,
            in2 => \N__9948\,
            in3 => \N__8211\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10733\,
            ce => \N__8301\,
            sr => \N__11161\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8374\,
            in1 => \N__9246\,
            in2 => \N__6899\,
            in3 => \N__6846\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10733\,
            ce => \N__8301\,
            sr => \N__11161\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7755\,
            in1 => \N__7597\,
            in2 => \N__7452\,
            in3 => \N__7380\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10736\,
            ce => \N__7341\,
            sr => \N__11157\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8429\,
            in2 => \_gnd_net_\,
            in3 => \N__7276\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_401_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__7335\,
            in1 => \N__7314\,
            in2 => \N__7281\,
            in3 => \N__10941\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10741\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7270\,
            in1 => \N__9192\,
            in2 => \N__9619\,
            in3 => \N__7253\,
            lcout => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__9194\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7237\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000100010"
        )
    port map (
            in0 => \N__10947\,
            in1 => \N__7164\,
            in2 => \N__7194\,
            in3 => \N__9613\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111101"
        )
    port map (
            in0 => \N__9143\,
            in1 => \N__9193\,
            in2 => \N__9620\,
            in3 => \N__7187\,
            lcout => \U712_REG_SM.STATE_COUNTc_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_170_i_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__7157\,
            in1 => \N__9801\,
            in2 => \N__8673\,
            in3 => \N__7145\,
            lcout => \N_170_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9197\,
            in2 => \_gnd_net_\,
            in3 => \N__9593\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__10959\,
            in1 => \N__8448\,
            in2 => \N__7968\,
            in3 => \N__9145\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10750\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__9234\,
            in1 => \N__9196\,
            in2 => \_gnd_net_\,
            in3 => \N__9592\,
            lcout => \U712_REG_SM.N_302\,
            ltout => \U712_REG_SM.N_302_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__10960\,
            in1 => \N__7910\,
            in2 => \N__7959\,
            in3 => \N__9235\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10750\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.N_160_i_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001010000"
        )
    port map (
            in0 => \N__7949\,
            in1 => \N__11952\,
            in2 => \N__9055\,
            in3 => \N__11874\,
            lcout => \N_160_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__7909\,
            in1 => \N__9195\,
            in2 => \_gnd_net_\,
            in3 => \N__9591\,
            lcout => \U712_REG_SM.N_404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111100011111100"
        )
    port map (
            in0 => \N__9101\,
            in1 => \N__7815\,
            in2 => \N__8664\,
            in3 => \N__9724\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10757\,
            ce => 'H',
            sr => \N__11154\
        );

    \U712_REG_SM.C1_SYNC_0_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7797\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10757\,
            ce => 'H',
            sr => \N__11154\
        );

    \U712_REG_SM.C1_SYNC_1_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7761\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10757\,
            ce => 'H',
            sr => \N__11154\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__9529\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11216\,
            lcout => \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10998\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8100\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8659\,
            in2 => \_gnd_net_\,
            in3 => \N__8099\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__9729\,
            in1 => \_gnd_net_\,
            in2 => \N__9105\,
            in3 => \N__10997\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9617\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10764\,
            ce => \N__8067\,
            sr => \N__11150\
        );

    \U712_CHIP_RAM.RASn_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8019\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10718\,
            ce => 'H',
            sr => \N__11197\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11733\,
            in1 => \N__11548\,
            in2 => \_gnd_net_\,
            in3 => \N__10147\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11286\,
            ce => \N__11255\,
            sr => \N__11167\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10148\,
            in1 => \_gnd_net_\,
            in2 => \N__11553\,
            in3 => \N__11042\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11286\,
            ce => \N__11255\,
            sr => \N__11167\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNIE8IL_0_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8010\,
            in2 => \_gnd_net_\,
            in3 => \N__10027\,
            lcout => \U712_CHIP_RAM.N_309\,
            ltout => \U712_CHIP_RAM.N_309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__9043\,
            in1 => \N__11792\,
            in2 => \N__7971\,
            in3 => \N__9448\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001111"
        )
    port map (
            in0 => \N__9044\,
            in1 => \N__11793\,
            in2 => \N__8388\,
            in3 => \N__9449\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8322\,
            in2 => \N__8316\,
            in3 => \N__8145\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10721\,
            ce => \N__8291\,
            sr => \N__11159\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8241\,
            in1 => \N__8225\,
            in2 => \_gnd_net_\,
            in3 => \N__9452\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9455\,
            in1 => \N__9047\,
            in2 => \N__8214\,
            in3 => \N__11685\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8195\,
            in1 => \N__8163\,
            in2 => \_gnd_net_\,
            in3 => \N__9450\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9453\,
            in1 => \N__9045\,
            in2 => \N__8148\,
            in3 => \N__11565\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8139\,
            in1 => \N__8124\,
            in2 => \_gnd_net_\,
            in3 => \N__9451\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9454\,
            in1 => \N__9046\,
            in2 => \N__8109\,
            in3 => \N__10164\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9039\,
            in1 => \N__8643\,
            in2 => \N__9446\,
            in3 => \N__9936\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_3_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10840\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10779\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10730\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_RNI8MQ3_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9097\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__9684\,
            in1 => \N__8514\,
            in2 => \_gnd_net_\,
            in3 => \N__8859\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10737\,
            ce => 'H',
            sr => \N__11155\
        );

    \U712_REG_SM.C3_SYNC_0_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8477\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10737\,
            ce => 'H',
            sr => \N__11155\
        );

    \U712_REG_SM.C3_SYNC_1_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8454\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10737\,
            ce => 'H',
            sr => \N__11155\
        );

    \U712_REG_SM.START_RST_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__8430\,
            in1 => \N__8447\,
            in2 => \_gnd_net_\,
            in3 => \N__9144\,
            lcout => \U712_REG_SM.START_RSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10737\,
            ce => 'H',
            sr => \N__11155\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000000"
        )
    port map (
            in0 => \N__9789\,
            in1 => \N__9869\,
            in2 => \N__9921\,
            in3 => \N__9051\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_443_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_54_i_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__8779\,
            in1 => \N__11951\,
            in2 => \N__8418\,
            in3 => \N__8722\,
            lcout => \N_54_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001111"
        )
    port map (
            in0 => \N__9228\,
            in1 => \N__9181\,
            in2 => \N__9146\,
            in3 => \N__9577\,
            lcout => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110111"
        )
    port map (
            in0 => \N__8814\,
            in1 => \N__9668\,
            in2 => \N__8853\,
            in3 => \N__9720\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_452_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__9669\,
            in1 => \N__10961\,
            in2 => \N__9108\,
            in3 => \N__9096\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10742\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__9870\,
            in1 => \N__9790\,
            in2 => \N__9057\,
            in3 => \N__9920\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_421_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_168_i_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__8721\,
            in1 => \N__11950\,
            in2 => \N__8883\,
            in3 => \N__8778\,
            lcout => \N_168_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__8813\,
            in1 => \N__8849\,
            in2 => \_gnd_net_\,
            in3 => \N__9667\,
            lcout => \U712_CYCLE_TERM.N_326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8848\,
            in2 => \_gnd_net_\,
            in3 => \N__8812\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__11850\,
            in1 => \N__8780\,
            in2 => \_gnd_net_\,
            in3 => \N__8723\,
            lcout => \U712_BYTE_ENABLE.N_425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10962\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8663\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__9728\,
            in1 => \N__9699\,
            in2 => \N__9693\,
            in3 => \N__9680\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10752\,
            ce => 'H',
            sr => \N__11149\
        );

    \U712_REG_SM.LDSn_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__9600\,
            in1 => \N__9654\,
            in2 => \N__9638\,
            in3 => \N__9533\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10752\,
            ce => 'H',
            sr => \N__11149\
        );

    \U712_REG_SM.UDSn_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111110101100"
        )
    port map (
            in0 => \N__9494\,
            in1 => \N__9601\,
            in2 => \N__9534\,
            in3 => \N__9909\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10752\,
            ce => 'H',
            sr => \N__11149\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10999\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_i_i_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010110000"
        )
    port map (
            in0 => \N__9775\,
            in1 => \N__9867\,
            in2 => \N__10397\,
            in3 => \N__10478\,
            lcout => \N_166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9456\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10719\,
            ce => 'H',
            sr => \N__11191\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10305\,
            in1 => \N__11530\,
            in2 => \_gnd_net_\,
            in3 => \N__11673\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__11256\,
            sr => \N__11170\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11669\,
            in1 => \N__11495\,
            in2 => \_gnd_net_\,
            in3 => \N__10304\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11284\,
            ce => \N__11253\,
            sr => \N__11162\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11500\,
            in1 => \N__11732\,
            in2 => \_gnd_net_\,
            in3 => \N__11767\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11284\,
            ce => \N__11253\,
            sr => \N__11162\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10206\,
            in1 => \N__11496\,
            in2 => \_gnd_net_\,
            in3 => \N__10241\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11284\,
            ce => \N__11253\,
            sr => \N__11162\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10242\,
            in1 => \_gnd_net_\,
            in2 => \N__11529\,
            in3 => \N__11766\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11284\,
            ce => \N__11253\,
            sr => \N__11162\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10202\,
            in1 => \N__11490\,
            in2 => \_gnd_net_\,
            in3 => \N__10296\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__11251\,
            sr => \N__11158\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__11778\,
            in1 => \_gnd_net_\,
            in2 => \N__11528\,
            in3 => \N__10240\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__11251\,
            sr => \N__11158\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__10509\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10420\,
            lcout => \U712_BYTE_ENABLE.N_298_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_RNO_0_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__10584\,
            in1 => \N__9854\,
            in2 => \N__10422\,
            in3 => \N__10508\,
            lcout => \U712_REG_SM.N_459\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_390_i_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000101000"
        )
    port map (
            in0 => \N__9793\,
            in1 => \N__10499\,
            in2 => \N__10416\,
            in3 => \N__9873\,
            lcout => \N_390_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_389_i_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000010100"
        )
    port map (
            in0 => \N__9792\,
            in1 => \N__10498\,
            in2 => \N__10415\,
            in3 => \N__9872\,
            lcout => \N_389_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100110000"
        )
    port map (
            in0 => \N__9871\,
            in1 => \N__9791\,
            in2 => \N__10507\,
            in3 => \N__10398\,
            lcout => \N_189\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11535\,
            in1 => \N__11610\,
            in2 => \_gnd_net_\,
            in3 => \N__11667\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11285\,
            ce => \N__11259\,
            sr => \N__11186\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10303\,
            in1 => \N__11494\,
            in2 => \_gnd_net_\,
            in3 => \N__10195\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11282\,
            ce => \N__11257\,
            sr => \N__11171\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10231\,
            in1 => \N__11470\,
            in2 => \_gnd_net_\,
            in3 => \N__10194\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__11252\,
            sr => \N__11163\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10133\,
            in1 => \N__11471\,
            in2 => \_gnd_net_\,
            in3 => \N__11731\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__11252\,
            sr => \N__11163\
        );

    \U712_CHIP_RAM.CRCSn_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10091\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10724\,
            ce => 'H',
            sr => \N__11196\
        );

    \U712_CHIP_RAM.WEn_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10032\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10729\,
            ce => 'H',
            sr => \N__11193\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11534\,
            in1 => \N__11622\,
            in2 => \_gnd_net_\,
            in3 => \N__11372\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__11261\,
            sr => \N__11192\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11321\,
            in1 => \N__11533\,
            in2 => \_gnd_net_\,
            in3 => \N__11364\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__11260\,
            sr => \N__11187\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11532\,
            in1 => \N__11618\,
            in2 => \_gnd_net_\,
            in3 => \N__11371\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11281\,
            ce => \N__11258\,
            sr => \N__11177\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11777\,
            in1 => \N__11446\,
            in2 => \_gnd_net_\,
            in3 => \N__11730\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__11254\,
            sr => \N__11172\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11668\,
            in1 => \N__11445\,
            in2 => \_gnd_net_\,
            in3 => \N__11611\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__11254\,
            sr => \N__11172\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11539\,
            in1 => \N__11373\,
            in2 => \_gnd_net_\,
            in3 => \N__11325\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11283\,
            ce => \N__11262\,
            sr => \N__11194\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10876\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11016\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11058\,
            in1 => \N__10875\,
            in2 => \_gnd_net_\,
            in3 => \N__11043\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_2_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10785\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_0_m2_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010101010101"
        )
    port map (
            in0 => \N__10620\,
            in1 => \N__10583\,
            in2 => \N__11923\,
            in3 => \N__11835\,
            lcout => \DRDDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

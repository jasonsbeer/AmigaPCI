-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 7 2025 10:58:53

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    TT : in std_logic_vector(1 downto 0);
    TM : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(31 downto 1);
    D : inout std_logic_vector(7 downto 4);
    RESETn : in std_logic;
    OVL : in std_logic;
    CONFIGENn : out std_logic;
    PIO_S0 : out std_logic;
    PORTSIZE : out std_logic;
    TICK60 : out std_logic;
    CIACS0n : out std_logic;
    CPUCONFn : in std_logic;
    CLK6 : in std_logic;
    CLK_CIA : out std_logic;
    BUFENn : out std_logic;
    AUTOBOOT : in std_logic;
    RnW : in std_logic;
    PIO_P2 : out std_logic;
    CIACS1n : out std_logic;
    BRIDGE_ENn : out std_logic;
    PIO_S1 : out std_logic;
    ATA_MODE_S : in std_logic;
    PIO_P0 : out std_logic;
    TICK50 : out std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : out std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    REGSPACEn : out std_logic;
    TSn : in std_logic;
    RTC_ENn : out std_logic;
    PIO_S2 : out std_logic;
    ATA_ENn : out std_logic;
    TACKn : inout std_logic;
    ATA_MODE_P : in std_logic;
    ROMENn : out std_logic;
    PIO_P1 : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__11402\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4077\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \PIO_S0_c\ : std_logic;
signal \GNDG0\ : std_logic;
signal \PIO_P0_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_25\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_26\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_8_cascade_\ : std_logic;
signal \A_c_24\ : std_logic;
signal \U409_AUTOCONFIG.N_270\ : std_logic;
signal \U409_AUTOCONFIG.N_271\ : std_logic;
signal \U409_AUTOCONFIG.N_433_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_433\ : std_logic;
signal \U409_AUTOCONFIG.N_373\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_2_3_0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0_0\ : std_logic;
signal \U409_AUTOCONFIG.N_269\ : std_logic;
signal \U409_AUTOCONFIG.N_370\ : std_logic;
signal \U409_AUTOCONFIG.N_195_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_383\ : std_logic;
signal \U409_AUTOCONFIG.N_274\ : std_logic;
signal \U409_AUTOCONFIG.N_383_cascade_\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \U409_ADDRESS_DECODE.N_345\ : std_logic;
signal \U409_ADDRESS_DECODE.N_344\ : std_logic;
signal \U409_AUTOCONFIG.N_288_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_a2Z0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.N_405_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_414\ : std_logic;
signal \U409_AUTOCONFIG.N_285\ : std_logic;
signal \U409_AUTOCONFIG.N_9\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0_1\ : std_logic;
signal \U409_AUTOCONFIG.N_405\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTc_0_1\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTc_0_0\ : std_logic;
signal \U409_AUTOCONFIG.N_286\ : std_logic;
signal \U409_AUTOCONFIG.AC_START_RNI3D7VZ0Z2\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\ : std_logic;
signal \U409_AUTOCONFIG.N_287\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U409_AUTOCONFIG.N_273\ : std_logic;
signal \U409_AUTOCONFIG.N_400\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_10\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_11\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_9_cascade_\ : std_logic;
signal \N_374\ : std_logic;
signal \N_401_cascade_\ : std_logic;
signal \N_436\ : std_logic;
signal \N_265_i\ : std_logic;
signal \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_o2_4\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ1Z_0\ : std_logic;
signal \N_124\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_1_0_a2_0Z0Z_2\ : std_logic;
signal \CPUCONFn_c\ : std_logic;
signal \U409_AUTOCONFIG.AC_STARTZ0\ : std_logic;
signal \INVU409_AUTOCONFIG.STATE_0C_net\ : std_logic;
signal \N_354_cascade_\ : std_logic;
signal \D_1_i\ : std_logic;
signal \AUTOBOOT_c\ : std_logic;
signal \U409_AUTOCONFIG.N_360\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U409_AUTOCONFIG.N_276\ : std_logic;
signal \U409_ADDRESS_DECODE.PORTSIZE_iZ0Z_1_cascade_\ : std_logic;
signal \N_139\ : std_logic;
signal \U409_ADDRESS_DECODE.N_343\ : std_logic;
signal \TM_c_1\ : std_logic;
signal \TM_c_0\ : std_logic;
signal \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_o2_5\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\ : std_logic;
signal \N_126\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net\ : std_logic;
signal \N_96\ : std_logic;
signal \A_c_29\ : std_logic;
signal \BRIDGE_BASE_1\ : std_logic;
signal \A_c_28\ : std_logic;
signal \BRIDGE_BASE_0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0Z0Z_0\ : std_logic;
signal \A_c_31\ : std_logic;
signal \BRIDGE_BASE_3\ : std_logic;
signal \BRIDGE_BASE_2\ : std_logic;
signal \A_c_30\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0Z0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\ : std_logic;
signal \U409_AUTOCONFIG.STATEZ0Z_0\ : std_logic;
signal \INVU409_AUTOCONFIG.AC_TACKC_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_a2_3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_268_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\ : std_logic;
signal \N_130\ : std_logic;
signal \ATA_BASE_4\ : std_logic;
signal \ATA_BASE_5\ : std_logic;
signal \D_in_4\ : std_logic;
signal \D_in_5\ : std_logic;
signal \D_in_6\ : std_logic;
signal \INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net\ : std_logic;
signal \ATA_BASE_6\ : std_logic;
signal \ATA_BASE_1\ : std_logic;
signal \ATA_BASE_0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7Z0Z_0_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_7_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_EN_2_0_o2_3_cascade_\ : std_logic;
signal \A_c_18\ : std_logic;
signal \ATA_BASE_2\ : std_logic;
signal \U409_ADDRESS_DECODE.N_183_i\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_EN_2_0_o2_2\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_2\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_7\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_o2dupZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_ATA_ENn_i_0Z0Z_3_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_ENZ0\ : std_logic;
signal \N_107\ : std_logic;
signal \A_c_16\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_CONFZ0\ : std_logic;
signal \N_128\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_268\ : std_logic;
signal \U409_TRANSFER_ACK.N_237\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\ : std_logic;
signal \RnW_c\ : std_logic;
signal \N_356\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_TRANSFER_ACK.N_346_cascade_\ : std_logic;
signal \N_434\ : std_logic;
signal \N_190_cascade_\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \A_c_21\ : std_logic;
signal \N_351\ : std_logic;
signal \N_436_i\ : std_logic;
signal \A_c_17\ : std_logic;
signal \N_431\ : std_logic;
signal \A_c_22\ : std_logic;
signal \N_401\ : std_logic;
signal \N_431_cascade_\ : std_logic;
signal \N_422\ : std_logic;
signal \A_c_19\ : std_logic;
signal \ATA_BASE_7\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_5\ : std_logic;
signal \N_361\ : std_logic;
signal \D_in_7\ : std_logic;
signal \ATA_BASE_3\ : std_logic;
signal \INVU409_AUTOCONFIG.ATA_BASE_ness_3C_net\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_1_0_0\ : std_logic;
signal \U409_AUTOCONFIG.N_172\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONFZ0\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_1_0_a2_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \CONFIGENn_c\ : std_logic;
signal \INVU409_AUTOCONFIG.CONFIGENnC_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \AC_TACK\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_159\ : std_logic;
signal \U409_TRANSFER_ACK.N_380\ : std_logic;
signal \U409_TRANSFER_ACK.N_380_cascade_\ : std_logic;
signal \N_190\ : std_logic;
signal \N_297\ : std_logic;
signal \N_94_i\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS1n_i\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_289\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_OUTnC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_379\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_307\ : std_logic;
signal \U409_TRANSFER_ACK.N_381\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROMENn_e_1\ : std_logic;
signal \ROMENn_c\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \N_357\ : std_logic;
signal \N_339\ : std_logic;
signal \TCIn_1_i\ : std_logic;
signal \CLK40_IN_c_g\ : std_logic;
signal \GB_BUFFER_CLK40_IN_c_g_THRU_CO\ : std_logic;
signal \CIA_ENABLE\ : std_logic;
signal \CIA_ENABLE_cascade_\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS0n_i\ : std_logic;
signal \U409_TICK.TICK603_10_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.m12_i_a2_1_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.m12_i_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_293\ : std_logic;
signal \U409_TRANSFER_ACK.N_191\ : std_logic;
signal \U409_TRANSFER_ACK.N_191_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_223\ : std_logic;
signal \U409_TRANSFER_ACK.i5_mux_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_290\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \OVL_c\ : std_logic;
signal \N_429\ : std_logic;
signal \N_348\ : std_logic;
signal \N_156_i\ : std_logic;
signal \N_264_i\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \bfn_13_6_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.TICK603_11\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_CIA.CLK_CIA6_0_a2_0_cascade_\ : std_logic;
signal \U409_CIA.CLK_CIA6_cascade_\ : std_logic;
signal \CLK_CIA_c\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_3_0_a2_0_cascade_\ : std_logic;
signal \U409_CIA.VMA_3_0_a2_2\ : std_logic;
signal \U409_CIA.VMA_RNOZ0Z_1_cascade_\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \bfn_14_5_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.TICK603_8\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_5\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_6\ : std_logic;
signal \U409_CIA.N_427\ : std_logic;
signal \U409_CIA.N_427_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_6\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_7\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_2_0_a2_2_cascade_\ : std_logic;
signal \U409_CIA.N_420\ : std_logic;
signal \U409_CIA.CLK_CIA_RNOZ0Z_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a2_2\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \PIO_P1_wire\ : std_logic;
signal \CPUCONFn_wire\ : std_logic;
signal \RTC_ENn_wire\ : std_logic;
signal \ATA_MODE_P_wire\ : std_logic;
signal \TM_wire\ : std_logic_vector(1 downto 0);
signal \RAMSPACEn_wire\ : std_logic;
signal \ROMENn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \AUTOBOOT_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \PIO_P2_wire\ : std_logic;
signal \BRIDGE_ENn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CIACS0n_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CONFIGENn_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \PIO_P0_wire\ : std_logic;
signal \ATA_MODE_S_wire\ : std_logic;
signal \ATA_ENn_wire\ : std_logic;
signal \CIACS1n_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \CLK_CIA_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \PIO_S0_wire\ : std_logic;
signal \PIO_S2_wire\ : std_logic;
signal \PIO_S1_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    \CLK40_IN_wire\ <= CLK40_IN;
    \A_wire\ <= A;
    \TT_wire\ <= TT;
    PIO_P1 <= \PIO_P1_wire\;
    \CPUCONFn_wire\ <= CPUCONFn;
    RTC_ENn <= \RTC_ENn_wire\;
    \ATA_MODE_P_wire\ <= ATA_MODE_P;
    \TM_wire\ <= TM;
    RAMSPACEn <= \RAMSPACEn_wire\;
    ROMENn <= \ROMENn_wire\;
    TBIn <= \TBIn_wire\;
    \AUTOBOOT_wire\ <= AUTOBOOT;
    \TSn_wire\ <= TSn;
    PORTSIZE <= \PORTSIZE_wire\;
    PIO_P2 <= \PIO_P2_wire\;
    BRIDGE_ENn <= \BRIDGE_ENn_wire\;
    \RESETn_wire\ <= RESETn;
    CIACS0n <= \CIACS0n_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TCIn <= \TCIn_wire\;
    \RnW_wire\ <= RnW;
    CONFIGENn <= \CONFIGENn_wire\;
    TICK60 <= \TICK60_wire\;
    PIO_P0 <= \PIO_P0_wire\;
    \ATA_MODE_S_wire\ <= ATA_MODE_S;
    ATA_ENn <= \ATA_ENn_wire\;
    CIACS1n <= \CIACS1n_wire\;
    REGSPACEn <= \REGSPACEn_wire\;
    CLK_CIA <= \CLK_CIA_wire\;
    BUFENn <= \BUFENn_wire\;
    PIO_S0 <= \PIO_S0_wire\;
    PIO_S2 <= \PIO_S2_wire\;
    PIO_S1 <= \PIO_S1_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__8292\,
            RESETB => \N__10619\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11400\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11402\,
            DIN => \N__11401\,
            DOUT => \N__11400\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11402\,
            PADOUT => \N__11401\,
            PADIN => \N__11400\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11390\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11392\,
            DIN => \N__11391\,
            DOUT => \N__11390\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11392\,
            PADOUT => \N__11391\,
            PADIN => \N__11390\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11380\,
            GLOBALBUFFEROUTPUT => \CLK40_IN_c_g\
        );

    \CLK40_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11382\,
            DIN => \N__11381\,
            DOUT => \N__11380\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11382\,
            PADOUT => \N__11381\,
            PADIN => \N__11380\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11371\,
            DIN => \N__11370\,
            DOUT => \N__11369\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11371\,
            PADOUT => \N__11370\,
            PADIN => \N__11369\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11362\,
            DIN => \N__11361\,
            DOUT => \N__11360\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11362\,
            PADOUT => \N__11361\,
            PADIN => \N__11360\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_P1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11353\,
            DIN => \N__11352\,
            DOUT => \N__11351\,
            PACKAGEPIN => \PIO_P1_wire\
        );

    \PIO_P1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11353\,
            PADOUT => \N__11352\,
            PADIN => \N__11351\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10623\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11344\,
            DIN => \N__11343\,
            DOUT => \N__11342\,
            PACKAGEPIN => D(7)
        );

    \D_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11344\,
            PADOUT => \N__11343\,
            PADIN => \N__11342\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5328\,
            DIN0 => \D_in_7\,
            DOUT0 => \N__5907\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11335\,
            DIN => \N__11334\,
            DOUT => \N__11333\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11335\,
            PADOUT => \N__11334\,
            PADIN => \N__11333\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUCONFn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11326\,
            DIN => \N__11325\,
            DOUT => \N__11324\,
            PACKAGEPIN => \CPUCONFn_wire\
        );

    \CPUCONFn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11326\,
            PADOUT => \N__11325\,
            PADIN => \N__11324\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CPUCONFn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RTC_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11317\,
            DIN => \N__11316\,
            DOUT => \N__11315\,
            PACKAGEPIN => \RTC_ENn_wire\
        );

    \RTC_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11317\,
            PADOUT => \N__11316\,
            PADIN => \N__11315\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6639\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11308\,
            DIN => \N__11307\,
            DOUT => \N__11306\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11308\,
            PADOUT => \N__11307\,
            PADIN => \N__11306\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ATA_MODE_P_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11299\,
            DIN => \N__11298\,
            DOUT => \N__11297\,
            PACKAGEPIN => \ATA_MODE_P_wire\
        );

    \ATA_MODE_P_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11299\,
            PADOUT => \N__11298\,
            PADIN => \N__11297\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PIO_P0_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11290\,
            DIN => \N__11289\,
            DOUT => \N__11288\,
            PACKAGEPIN => D(4)
        );

    \D_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11290\,
            PADOUT => \N__11289\,
            PADIN => \N__11288\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5306\,
            DIN0 => \D_in_4\,
            DOUT0 => \N__4923\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11281\,
            DIN => \N__11280\,
            DOUT => \N__11279\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11281\,
            PADOUT => \N__11280\,
            PADIN => \N__11279\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11272\,
            DIN => \N__11271\,
            DOUT => \N__11270\,
            PACKAGEPIN => \TM_wire\(1)
        );

    \TM_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11272\,
            PADOUT => \N__11271\,
            PADIN => \N__11270\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11263\,
            DIN => \N__11262\,
            DOUT => \N__11261\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11263\,
            PADOUT => \N__11262\,
            PADIN => \N__11261\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11254\,
            DIN => \N__11253\,
            DOUT => \N__11252\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11254\,
            PADOUT => \N__11253\,
            PADIN => \N__11252\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9192\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11245\,
            DIN => \N__11244\,
            DOUT => \N__11243\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11245\,
            PADOUT => \N__11244\,
            PADIN => \N__11243\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11236\,
            DIN => \N__11235\,
            DOUT => \N__11234\,
            PACKAGEPIN => \ROMENn_wire\
        );

    \ROMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11236\,
            PADOUT => \N__11235\,
            PADIN => \N__11234\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8664\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11227\,
            DIN => \N__11226\,
            DOUT => \N__11225\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11227\,
            PADOUT => \N__11226\,
            PADIN => \N__11225\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8490\,
            DIN0 => OPEN,
            DOUT0 => \N__8258\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AUTOBOOT_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11218\,
            DIN => \N__11217\,
            DOUT => \N__11216\,
            PACKAGEPIN => \AUTOBOOT_wire\
        );

    \AUTOBOOT_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11218\,
            PADOUT => \N__11217\,
            PADIN => \N__11216\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AUTOBOOT_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11209\,
            DIN => \N__11208\,
            DOUT => \N__11207\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11209\,
            PADOUT => \N__11208\,
            PADIN => \N__11207\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11200\,
            DIN => \N__11199\,
            DOUT => \N__11198\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11200\,
            PADOUT => \N__11199\,
            PADIN => \N__11198\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5085\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_P2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11191\,
            DIN => \N__11190\,
            DOUT => \N__11189\,
            PACKAGEPIN => \PIO_P2_wire\
        );

    \PIO_P2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11191\,
            PADOUT => \N__11190\,
            PADIN => \N__11189\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10605\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11182\,
            DIN => \N__11181\,
            DOUT => \N__11180\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11182\,
            PADOUT => \N__11181\,
            PADIN => \N__11180\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BRIDGE_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11173\,
            DIN => \N__11172\,
            DOUT => \N__11171\,
            PACKAGEPIN => \BRIDGE_ENn_wire\
        );

    \BRIDGE_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11173\,
            PADOUT => \N__11172\,
            PADIN => \N__11171\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5472\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11164\,
            DIN => \N__11163\,
            DOUT => \N__11162\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11164\,
            PADOUT => \N__11163\,
            PADIN => \N__11162\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11155\,
            DIN => \N__11154\,
            DOUT => \N__11153\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11155\,
            PADOUT => \N__11154\,
            PADIN => \N__11153\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11146\,
            DIN => \N__11145\,
            DOUT => \N__11144\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11146\,
            PADOUT => \N__11145\,
            PADIN => \N__11144\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11137\,
            DIN => \N__11136\,
            DOUT => \N__11135\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11137\,
            PADOUT => \N__11136\,
            PADIN => \N__11135\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11128\,
            DIN => \N__11127\,
            DOUT => \N__11126\,
            PACKAGEPIN => \CIACS0n_wire\
        );

    \CIACS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11128\,
            PADOUT => \N__11127\,
            PADIN => \N__11126\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8757\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11119\,
            DIN => \N__11118\,
            DOUT => \N__11117\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11119\,
            PADOUT => \N__11118\,
            PADIN => \N__11117\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10185\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11110\,
            DIN => \N__11109\,
            DOUT => \N__11108\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11110\,
            PADOUT => \N__11109\,
            PADIN => \N__11108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11101\,
            DIN => \N__11100\,
            DOUT => \N__11099\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11101\,
            PADOUT => \N__11100\,
            PADIN => \N__11099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11092\,
            DIN => \N__11091\,
            DOUT => \N__11090\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11092\,
            PADOUT => \N__11091\,
            PADIN => \N__11090\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11083\,
            DIN => \N__11082\,
            DOUT => \N__11081\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11083\,
            PADOUT => \N__11082\,
            PADIN => \N__11081\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11074\,
            DIN => \N__11073\,
            DOUT => \N__11072\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11074\,
            PADOUT => \N__11073\,
            PADIN => \N__11072\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8406\,
            DIN0 => OPEN,
            DOUT0 => \N__8259\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11065\,
            DIN => \N__11064\,
            DOUT => \N__11063\,
            PACKAGEPIN => D(5)
        );

    \D_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11065\,
            PADOUT => \N__11064\,
            PADIN => \N__11063\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5323\,
            DIN0 => \D_in_5\,
            DOUT0 => \N__5487\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11056\,
            DIN => \N__11055\,
            DOUT => \N__11054\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11056\,
            PADOUT => \N__11055\,
            PADIN => \N__11054\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11047\,
            DIN => \N__11046\,
            DOUT => \N__11045\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11047\,
            PADOUT => \N__11046\,
            PADIN => \N__11045\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11038\,
            DIN => \N__11037\,
            DOUT => \N__11036\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11038\,
            PADOUT => \N__11037\,
            PADIN => \N__11036\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CONFIGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11029\,
            DIN => \N__11028\,
            DOUT => \N__11027\,
            PACKAGEPIN => \CONFIGENn_wire\
        );

    \CONFIGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11029\,
            PADOUT => \N__11028\,
            PADIN => \N__11027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7212\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11020\,
            DIN => \N__11019\,
            DOUT => \N__11018\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11020\,
            PADOUT => \N__11019\,
            PADIN => \N__11018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9597\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11011\,
            DIN => \N__11010\,
            DOUT => \N__11009\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11011\,
            PADOUT => \N__11010\,
            PADIN => \N__11009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_P0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11002\,
            DIN => \N__11001\,
            DOUT => \N__11000\,
            PACKAGEPIN => \PIO_P0_wire\
        );

    \PIO_P0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11002\,
            PADOUT => \N__11001\,
            PADIN => \N__11000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4155\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ATA_MODE_S_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__10993\,
            DIN => \N__10992\,
            DOUT => \N__10991\,
            PACKAGEPIN => \ATA_MODE_S_wire\
        );

    \ATA_MODE_S_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10993\,
            PADOUT => \N__10992\,
            PADIN => \N__10991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PIO_S0_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10984\,
            DIN => \N__10983\,
            DOUT => \N__10982\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10984\,
            PADOUT => \N__10983\,
            PADIN => \N__10982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ATA_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10975\,
            DIN => \N__10974\,
            DOUT => \N__10973\,
            PACKAGEPIN => \ATA_ENn_wire\
        );

    \ATA_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10975\,
            PADOUT => \N__10974\,
            PADIN => \N__10973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6468\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10966\,
            DIN => \N__10965\,
            DOUT => \N__10964\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10966\,
            PADOUT => \N__10965\,
            PADIN => \N__10964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10957\,
            DIN => \N__10956\,
            DOUT => \N__10955\,
            PACKAGEPIN => \CIACS1n_wire\
        );

    \CIACS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10957\,
            PADOUT => \N__10956\,
            PADIN => \N__10955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7989\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10948\,
            DIN => \N__10947\,
            DOUT => \N__10946\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10948\,
            PADOUT => \N__10947\,
            PADIN => \N__10946\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4989\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10939\,
            DIN => \N__10938\,
            DOUT => \N__10937\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10939\,
            PADOUT => \N__10938\,
            PADIN => \N__10937\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_CIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10930\,
            DIN => \N__10929\,
            DOUT => \N__10928\,
            PACKAGEPIN => \CLK_CIA_wire\
        );

    \CLK_CIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10930\,
            PADOUT => \N__10929\,
            PADIN => \N__10928\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9564\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10921\,
            DIN => \N__10920\,
            DOUT => \N__10919\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10921\,
            PADOUT => \N__10920\,
            PADIN => \N__10919\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10912\,
            DIN => \N__10911\,
            DOUT => \N__10910\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__10912\,
            PADOUT => \N__10911\,
            PADIN => \N__10910\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8486\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__8246\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10903\,
            DIN => \N__10902\,
            DOUT => \N__10901\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10903\,
            PADOUT => \N__10902\,
            PADIN => \N__10901\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10894\,
            DIN => \N__10893\,
            DOUT => \N__10892\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10894\,
            PADOUT => \N__10893\,
            PADIN => \N__10892\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8022\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_S0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10885\,
            DIN => \N__10884\,
            DOUT => \N__10883\,
            PACKAGEPIN => \PIO_S0_wire\
        );

    \PIO_S0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10885\,
            PADOUT => \N__10884\,
            PADIN => \N__10883\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4134\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10876\,
            DIN => \N__10875\,
            DOUT => \N__10874\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10876\,
            PADOUT => \N__10875\,
            PADIN => \N__10874\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_S2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10867\,
            DIN => \N__10866\,
            DOUT => \N__10865\,
            PACKAGEPIN => \PIO_S2_wire\
        );

    \PIO_S2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10867\,
            PADOUT => \N__10866\,
            PADIN => \N__10865\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10618\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10858\,
            DIN => \N__10857\,
            DOUT => \N__10856\,
            PACKAGEPIN => D(6)
        );

    \D_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__10858\,
            PADOUT => \N__10857\,
            PADIN => \N__10856\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5324\,
            DIN0 => \D_in_6\,
            DOUT0 => \N__6339\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10849\,
            DIN => \N__10848\,
            DOUT => \N__10847\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10849\,
            PADOUT => \N__10848\,
            PADIN => \N__10847\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10840\,
            DIN => \N__10839\,
            DOUT => \N__10838\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10840\,
            PADOUT => \N__10839\,
            PADIN => \N__10838\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_S1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10831\,
            DIN => \N__10830\,
            DOUT => \N__10829\,
            PACKAGEPIN => \PIO_S1_wire\
        );

    \PIO_S1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10831\,
            PADOUT => \N__10830\,
            PADIN => \N__10829\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10598\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10822\,
            DIN => \N__10821\,
            DOUT => \N__10820\,
            PACKAGEPIN => \TM_wire\(0)
        );

    \TM_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10822\,
            PADOUT => \N__10821\,
            PADIN => \N__10820\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10813\,
            DIN => \N__10812\,
            DOUT => \N__10811\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10813\,
            PADOUT => \N__10812\,
            PADIN => \N__10811\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10804\,
            DIN => \N__10803\,
            DOUT => \N__10802\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10804\,
            PADOUT => \N__10803\,
            PADIN => \N__10802\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2593\ : InMux
    port map (
            O => \N__10785\,
            I => \N__10782\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__10782\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__2591\ : InMux
    port map (
            O => \N__10779\,
            I => \N__10761\
        );

    \I__2590\ : InMux
    port map (
            O => \N__10778\,
            I => \N__10761\
        );

    \I__2589\ : InMux
    port map (
            O => \N__10777\,
            I => \N__10761\
        );

    \I__2588\ : InMux
    port map (
            O => \N__10776\,
            I => \N__10761\
        );

    \I__2587\ : InMux
    port map (
            O => \N__10775\,
            I => \N__10761\
        );

    \I__2586\ : InMux
    port map (
            O => \N__10774\,
            I => \N__10754\
        );

    \I__2585\ : InMux
    port map (
            O => \N__10773\,
            I => \N__10754\
        );

    \I__2584\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10754\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__10761\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__10754\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2581\ : CascadeMux
    port map (
            O => \N__10749\,
            I => \N__10742\
        );

    \I__2580\ : InMux
    port map (
            O => \N__10748\,
            I => \N__10730\
        );

    \I__2579\ : InMux
    port map (
            O => \N__10747\,
            I => \N__10730\
        );

    \I__2578\ : InMux
    port map (
            O => \N__10746\,
            I => \N__10730\
        );

    \I__2577\ : InMux
    port map (
            O => \N__10745\,
            I => \N__10730\
        );

    \I__2576\ : InMux
    port map (
            O => \N__10742\,
            I => \N__10721\
        );

    \I__2575\ : InMux
    port map (
            O => \N__10741\,
            I => \N__10721\
        );

    \I__2574\ : InMux
    port map (
            O => \N__10740\,
            I => \N__10721\
        );

    \I__2573\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10721\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__10730\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__10721\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2570\ : CascadeMux
    port map (
            O => \N__10716\,
            I => \N__10709\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__10715\,
            I => \N__10706\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__10714\,
            I => \N__10702\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__10713\,
            I => \N__10697\
        );

    \I__2566\ : InMux
    port map (
            O => \N__10712\,
            I => \N__10688\
        );

    \I__2565\ : InMux
    port map (
            O => \N__10709\,
            I => \N__10688\
        );

    \I__2564\ : InMux
    port map (
            O => \N__10706\,
            I => \N__10688\
        );

    \I__2563\ : InMux
    port map (
            O => \N__10705\,
            I => \N__10688\
        );

    \I__2562\ : InMux
    port map (
            O => \N__10702\,
            I => \N__10683\
        );

    \I__2561\ : InMux
    port map (
            O => \N__10701\,
            I => \N__10683\
        );

    \I__2560\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10678\
        );

    \I__2559\ : InMux
    port map (
            O => \N__10697\,
            I => \N__10678\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__10688\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__10683\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__10678\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__10671\,
            I => \N__10668\
        );

    \I__2554\ : InMux
    port map (
            O => \N__10668\,
            I => \N__10664\
        );

    \I__2553\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10661\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10664\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__10661\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2550\ : ClkMux
    port map (
            O => \N__10656\,
            I => \N__10629\
        );

    \I__2549\ : ClkMux
    port map (
            O => \N__10655\,
            I => \N__10629\
        );

    \I__2548\ : ClkMux
    port map (
            O => \N__10654\,
            I => \N__10629\
        );

    \I__2547\ : ClkMux
    port map (
            O => \N__10653\,
            I => \N__10629\
        );

    \I__2546\ : ClkMux
    port map (
            O => \N__10652\,
            I => \N__10629\
        );

    \I__2545\ : ClkMux
    port map (
            O => \N__10651\,
            I => \N__10629\
        );

    \I__2544\ : ClkMux
    port map (
            O => \N__10650\,
            I => \N__10629\
        );

    \I__2543\ : ClkMux
    port map (
            O => \N__10649\,
            I => \N__10629\
        );

    \I__2542\ : ClkMux
    port map (
            O => \N__10648\,
            I => \N__10629\
        );

    \I__2541\ : GlobalMux
    port map (
            O => \N__10629\,
            I => \N__10626\
        );

    \I__2540\ : gio2CtrlBuf
    port map (
            O => \N__10626\,
            I => \CLK6_c_g\
        );

    \I__2539\ : IoInMux
    port map (
            O => \N__10623\,
            I => \N__10620\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__10620\,
            I => \N__10615\
        );

    \I__2537\ : IoInMux
    port map (
            O => \N__10619\,
            I => \N__10612\
        );

    \I__2536\ : IoInMux
    port map (
            O => \N__10618\,
            I => \N__10609\
        );

    \I__2535\ : IoSpan4Mux
    port map (
            O => \N__10615\,
            I => \N__10606\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__10612\,
            I => \N__10602\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__10609\,
            I => \N__10599\
        );

    \I__2532\ : Span4Mux_s2_h
    port map (
            O => \N__10606\,
            I => \N__10595\
        );

    \I__2531\ : IoInMux
    port map (
            O => \N__10605\,
            I => \N__10592\
        );

    \I__2530\ : IoSpan4Mux
    port map (
            O => \N__10602\,
            I => \N__10589\
        );

    \I__2529\ : IoSpan4Mux
    port map (
            O => \N__10599\,
            I => \N__10586\
        );

    \I__2528\ : IoInMux
    port map (
            O => \N__10598\,
            I => \N__10583\
        );

    \I__2527\ : Sp12to4
    port map (
            O => \N__10595\,
            I => \N__10578\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__10592\,
            I => \N__10578\
        );

    \I__2525\ : Sp12to4
    port map (
            O => \N__10589\,
            I => \N__10575\
        );

    \I__2524\ : Sp12to4
    port map (
            O => \N__10586\,
            I => \N__10570\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__10583\,
            I => \N__10570\
        );

    \I__2522\ : Span12Mux_s9_h
    port map (
            O => \N__10578\,
            I => \N__10567\
        );

    \I__2521\ : Span12Mux_s9_v
    port map (
            O => \N__10575\,
            I => \N__10564\
        );

    \I__2520\ : Span12Mux_s1_h
    port map (
            O => \N__10570\,
            I => \N__10561\
        );

    \I__2519\ : Odrv12
    port map (
            O => \N__10567\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2518\ : Odrv12
    port map (
            O => \N__10564\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2517\ : Odrv12
    port map (
            O => \N__10561\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__10554\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__2515\ : InMux
    port map (
            O => \N__10551\,
            I => \N__10547\
        );

    \I__2514\ : InMux
    port map (
            O => \N__10550\,
            I => \N__10544\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__10547\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__10544\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2511\ : InMux
    port map (
            O => \N__10539\,
            I => \N__10535\
        );

    \I__2510\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10532\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__10535\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10532\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__10527\,
            I => \N__10521\
        );

    \I__2506\ : InMux
    port map (
            O => \N__10526\,
            I => \N__10518\
        );

    \I__2505\ : InMux
    port map (
            O => \N__10525\,
            I => \N__10515\
        );

    \I__2504\ : InMux
    port map (
            O => \N__10524\,
            I => \N__10512\
        );

    \I__2503\ : InMux
    port map (
            O => \N__10521\,
            I => \N__10509\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__10518\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__10515\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__10512\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__10509\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2498\ : InMux
    port map (
            O => \N__10500\,
            I => \N__10496\
        );

    \I__2497\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10493\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__10496\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__10493\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10488\,
            I => \N__10485\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__10485\,
            I => \N__10482\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__10482\,
            I => \U409_TICK.TICK503_11\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__10479\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__2490\ : InMux
    port map (
            O => \N__10476\,
            I => \N__10472\
        );

    \I__2489\ : InMux
    port map (
            O => \N__10475\,
            I => \N__10469\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__10472\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__10469\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__10464\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__2485\ : InMux
    port map (
            O => \N__10461\,
            I => \N__10458\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__10458\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__2483\ : InMux
    port map (
            O => \N__10455\,
            I => \N__10451\
        );

    \I__2482\ : InMux
    port map (
            O => \N__10454\,
            I => \N__10448\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__10451\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__10448\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__2479\ : InMux
    port map (
            O => \N__10443\,
            I => \N__10440\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__10440\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__2477\ : InMux
    port map (
            O => \N__10437\,
            I => \N__10434\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__10434\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__2475\ : InMux
    port map (
            O => \N__10431\,
            I => \N__10427\
        );

    \I__2474\ : InMux
    port map (
            O => \N__10430\,
            I => \N__10424\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__10427\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__10424\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__2471\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10415\
        );

    \I__2470\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10412\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__10415\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__10412\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2467\ : InMux
    port map (
            O => \N__10407\,
            I => \N__10403\
        );

    \I__2466\ : InMux
    port map (
            O => \N__10406\,
            I => \N__10400\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__10403\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__10400\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__10395\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__2462\ : InMux
    port map (
            O => \N__10392\,
            I => \N__10389\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__10389\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__2460\ : InMux
    port map (
            O => \N__10386\,
            I => \N__10382\
        );

    \I__2459\ : InMux
    port map (
            O => \N__10385\,
            I => \N__10379\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__10382\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__10379\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__10374\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_2_0_a2_2_cascade_\
        );

    \I__2455\ : InMux
    port map (
            O => \N__10371\,
            I => \N__10367\
        );

    \I__2454\ : InMux
    port map (
            O => \N__10370\,
            I => \N__10364\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__10367\,
            I => \U409_CIA.N_420\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__10364\,
            I => \U409_CIA.N_420\
        );

    \I__2451\ : InMux
    port map (
            O => \N__10359\,
            I => \N__10356\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10356\,
            I => \U409_CIA.CLK_CIA_RNOZ0Z_1\
        );

    \I__2449\ : CascadeMux
    port map (
            O => \N__10353\,
            I => \N__10345\
        );

    \I__2448\ : InMux
    port map (
            O => \N__10352\,
            I => \N__10337\
        );

    \I__2447\ : InMux
    port map (
            O => \N__10351\,
            I => \N__10337\
        );

    \I__2446\ : InMux
    port map (
            O => \N__10350\,
            I => \N__10337\
        );

    \I__2445\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10334\
        );

    \I__2444\ : InMux
    port map (
            O => \N__10348\,
            I => \N__10327\
        );

    \I__2443\ : InMux
    port map (
            O => \N__10345\,
            I => \N__10327\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10344\,
            I => \N__10327\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__10337\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__10334\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__10327\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__2438\ : CascadeMux
    port map (
            O => \N__10320\,
            I => \N__10313\
        );

    \I__2437\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10308\
        );

    \I__2436\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10301\
        );

    \I__2435\ : InMux
    port map (
            O => \N__10317\,
            I => \N__10301\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10316\,
            I => \N__10301\
        );

    \I__2433\ : InMux
    port map (
            O => \N__10313\,
            I => \N__10298\
        );

    \I__2432\ : InMux
    port map (
            O => \N__10312\,
            I => \N__10293\
        );

    \I__2431\ : InMux
    port map (
            O => \N__10311\,
            I => \N__10293\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__10308\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__10301\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__10298\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__10293\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2426\ : ClkMux
    port map (
            O => \N__10284\,
            I => \N__10275\
        );

    \I__2425\ : ClkMux
    port map (
            O => \N__10283\,
            I => \N__10275\
        );

    \I__2424\ : ClkMux
    port map (
            O => \N__10282\,
            I => \N__10275\
        );

    \I__2423\ : GlobalMux
    port map (
            O => \N__10275\,
            I => \N__10272\
        );

    \I__2422\ : gio2CtrlBuf
    port map (
            O => \N__10272\,
            I => \CLK28_IN_c_g\
        );

    \I__2421\ : InMux
    port map (
            O => \N__10269\,
            I => \N__10263\
        );

    \I__2420\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10260\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10267\,
            I => \N__10255\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10266\,
            I => \N__10255\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__10263\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__10260\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__10255\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10248\,
            I => \N__10241\
        );

    \I__2413\ : InMux
    port map (
            O => \N__10247\,
            I => \N__10236\
        );

    \I__2412\ : InMux
    port map (
            O => \N__10246\,
            I => \N__10236\
        );

    \I__2411\ : InMux
    port map (
            O => \N__10245\,
            I => \N__10231\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10231\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__10241\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__10236\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__10231\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2406\ : InMux
    port map (
            O => \N__10224\,
            I => \N__10218\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10223\,
            I => \N__10215\
        );

    \I__2404\ : InMux
    port map (
            O => \N__10222\,
            I => \N__10210\
        );

    \I__2403\ : InMux
    port map (
            O => \N__10221\,
            I => \N__10210\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__10218\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__10215\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__10210\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10203\,
            I => \N__10200\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__10200\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\
        );

    \I__2397\ : CascadeMux
    port map (
            O => \N__10197\,
            I => \N__10194\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10191\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__10191\,
            I => \N__10188\
        );

    \I__2394\ : Odrv4
    port map (
            O => \N__10188\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__2393\ : IoInMux
    port map (
            O => \N__10185\,
            I => \N__10182\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__10182\,
            I => \N__10179\
        );

    \I__2391\ : Span4Mux_s3_v
    port map (
            O => \N__10179\,
            I => \N__10176\
        );

    \I__2390\ : Span4Mux_v
    port map (
            O => \N__10176\,
            I => \N__10173\
        );

    \I__2389\ : Span4Mux_h
    port map (
            O => \N__10173\,
            I => \N__10169\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10172\,
            I => \N__10166\
        );

    \I__2387\ : Odrv4
    port map (
            O => \N__10169\,
            I => \TICK50_c\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__10166\,
            I => \TICK50_c\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10158\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10158\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10155\,
            I => \N__10151\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10148\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__10151\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__10148\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2379\ : InMux
    port map (
            O => \N__10143\,
            I => \N__10139\
        );

    \I__2378\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10136\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__10139\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__10136\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__10131\,
            I => \N__10127\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__10130\,
            I => \N__10124\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10127\,
            I => \N__10118\
        );

    \I__2372\ : InMux
    port map (
            O => \N__10124\,
            I => \N__10118\
        );

    \I__2371\ : InMux
    port map (
            O => \N__10123\,
            I => \N__10115\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__10118\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__10115\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10110\,
            I => \N__10106\
        );

    \I__2367\ : InMux
    port map (
            O => \N__10109\,
            I => \N__10103\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__10106\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__10103\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10098\,
            I => \N__10094\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10097\,
            I => \N__10091\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10094\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__10091\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__10086\,
            I => \N__10083\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10083\,
            I => \N__10079\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10076\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__10079\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10076\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10071\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__2354\ : InMux
    port map (
            O => \N__10068\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__2353\ : InMux
    port map (
            O => \N__10065\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__2352\ : InMux
    port map (
            O => \N__10062\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\
        );

    \I__2351\ : InMux
    port map (
            O => \N__10059\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\
        );

    \I__2350\ : InMux
    port map (
            O => \N__10056\,
            I => \N__10050\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10055\,
            I => \N__10050\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__10050\,
            I => \U409_CIA.N_427\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__10047\,
            I => \U409_CIA.N_427_cascade_\
        );

    \I__2346\ : InMux
    port map (
            O => \N__10044\,
            I => \N__10038\
        );

    \I__2345\ : InMux
    port map (
            O => \N__10043\,
            I => \N__10038\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__10038\,
            I => \N__10035\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__10035\,
            I => \U409_CIA.CIA_CLK_COUNT11\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10032\,
            I => \N__10027\
        );

    \I__2341\ : InMux
    port map (
            O => \N__10031\,
            I => \N__10022\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10030\,
            I => \N__10022\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__10027\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__10022\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__10017\,
            I => \N__10013\
        );

    \I__2336\ : InMux
    port map (
            O => \N__10016\,
            I => \N__10009\
        );

    \I__2335\ : InMux
    port map (
            O => \N__10013\,
            I => \N__10004\
        );

    \I__2334\ : InMux
    port map (
            O => \N__10012\,
            I => \N__10004\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__10009\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__10004\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__2331\ : InMux
    port map (
            O => \N__9999\,
            I => \N__9994\
        );

    \I__2330\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9989\
        );

    \I__2329\ : InMux
    port map (
            O => \N__9997\,
            I => \N__9989\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__9994\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__9989\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__2326\ : InMux
    port map (
            O => \N__9984\,
            I => \N__9981\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__9981\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__2324\ : InMux
    port map (
            O => \N__9978\,
            I => \N__9974\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__9977\,
            I => \N__9969\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__9974\,
            I => \N__9966\
        );

    \I__2321\ : InMux
    port map (
            O => \N__9973\,
            I => \N__9961\
        );

    \I__2320\ : InMux
    port map (
            O => \N__9972\,
            I => \N__9961\
        );

    \I__2319\ : InMux
    port map (
            O => \N__9969\,
            I => \N__9958\
        );

    \I__2318\ : Odrv4
    port map (
            O => \N__9966\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__9961\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__9958\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2315\ : InMux
    port map (
            O => \N__9951\,
            I => \N__9948\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__9948\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__2313\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9941\
        );

    \I__2312\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9938\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__9941\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__9938\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__2309\ : InMux
    port map (
            O => \N__9933\,
            I => \N__9929\
        );

    \I__2308\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9926\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__9929\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__9926\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__9921\,
            I => \N__9918\
        );

    \I__2304\ : InMux
    port map (
            O => \N__9918\,
            I => \N__9915\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__9915\,
            I => \N__9911\
        );

    \I__2302\ : InMux
    port map (
            O => \N__9914\,
            I => \N__9908\
        );

    \I__2301\ : Odrv4
    port map (
            O => \N__9911\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__9908\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__9903\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__2298\ : InMux
    port map (
            O => \N__9900\,
            I => \N__9897\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__9897\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__2296\ : InMux
    port map (
            O => \N__9894\,
            I => \N__9890\
        );

    \I__2295\ : InMux
    port map (
            O => \N__9893\,
            I => \N__9887\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__9890\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__9887\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__9882\,
            I => \N__9874\
        );

    \I__2291\ : InMux
    port map (
            O => \N__9881\,
            I => \N__9866\
        );

    \I__2290\ : InMux
    port map (
            O => \N__9880\,
            I => \N__9866\
        );

    \I__2289\ : InMux
    port map (
            O => \N__9879\,
            I => \N__9866\
        );

    \I__2288\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9861\
        );

    \I__2287\ : InMux
    port map (
            O => \N__9877\,
            I => \N__9861\
        );

    \I__2286\ : InMux
    port map (
            O => \N__9874\,
            I => \N__9856\
        );

    \I__2285\ : InMux
    port map (
            O => \N__9873\,
            I => \N__9856\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__9866\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__9861\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__9856\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2281\ : InMux
    port map (
            O => \N__9849\,
            I => \N__9838\
        );

    \I__2280\ : InMux
    port map (
            O => \N__9848\,
            I => \N__9838\
        );

    \I__2279\ : InMux
    port map (
            O => \N__9847\,
            I => \N__9835\
        );

    \I__2278\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9826\
        );

    \I__2277\ : InMux
    port map (
            O => \N__9845\,
            I => \N__9826\
        );

    \I__2276\ : InMux
    port map (
            O => \N__9844\,
            I => \N__9826\
        );

    \I__2275\ : InMux
    port map (
            O => \N__9843\,
            I => \N__9826\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__9838\,
            I => \N__9823\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__9835\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__9826\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__9823\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2270\ : CascadeMux
    port map (
            O => \N__9816\,
            I => \N__9810\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__9815\,
            I => \N__9807\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__9814\,
            I => \N__9804\
        );

    \I__2267\ : InMux
    port map (
            O => \N__9813\,
            I => \N__9790\
        );

    \I__2266\ : InMux
    port map (
            O => \N__9810\,
            I => \N__9790\
        );

    \I__2265\ : InMux
    port map (
            O => \N__9807\,
            I => \N__9790\
        );

    \I__2264\ : InMux
    port map (
            O => \N__9804\,
            I => \N__9790\
        );

    \I__2263\ : InMux
    port map (
            O => \N__9803\,
            I => \N__9790\
        );

    \I__2262\ : InMux
    port map (
            O => \N__9802\,
            I => \N__9787\
        );

    \I__2261\ : InMux
    port map (
            O => \N__9801\,
            I => \N__9784\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__9790\,
            I => \N__9781\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__9787\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__9784\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2257\ : Odrv12
    port map (
            O => \N__9781\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2256\ : InMux
    port map (
            O => \N__9774\,
            I => \N__9771\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__9771\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__2254\ : InMux
    port map (
            O => \N__9768\,
            I => \N__9764\
        );

    \I__2253\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9761\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__9764\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__9761\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2250\ : InMux
    port map (
            O => \N__9756\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__2249\ : InMux
    port map (
            O => \N__9753\,
            I => \bfn_14_6_0_\
        );

    \I__2248\ : InMux
    port map (
            O => \N__9750\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__2247\ : InMux
    port map (
            O => \N__9747\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__2246\ : InMux
    port map (
            O => \N__9744\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__2245\ : InMux
    port map (
            O => \N__9741\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__2244\ : InMux
    port map (
            O => \N__9738\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9735\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9732\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9729\,
            I => \N__9725\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9722\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__9725\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__9722\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9714\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__9714\,
            I => \U409_TICK.TICK603_8\
        );

    \I__2235\ : InMux
    port map (
            O => \N__9711\,
            I => \N__9708\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__9708\,
            I => \N__9705\
        );

    \I__2233\ : Span4Mux_h
    port map (
            O => \N__9705\,
            I => \N__9702\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__9702\,
            I => \U409_CIA.VMA_3_0_a2_2\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__9699\,
            I => \U409_CIA.VMA_RNOZ0Z_1_cascade_\
        );

    \I__2230\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9693\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__9693\,
            I => \N__9690\
        );

    \I__2228\ : Span4Mux_v
    port map (
            O => \N__9690\,
            I => \N__9685\
        );

    \I__2227\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9682\
        );

    \I__2226\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9679\
        );

    \I__2225\ : Odrv4
    port map (
            O => \N__9685\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__9682\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__9679\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2222\ : InMux
    port map (
            O => \N__9672\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__2221\ : InMux
    port map (
            O => \N__9669\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9666\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__2219\ : InMux
    port map (
            O => \N__9663\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__2218\ : InMux
    port map (
            O => \N__9660\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__2217\ : InMux
    port map (
            O => \N__9657\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__2216\ : InMux
    port map (
            O => \N__9654\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__2215\ : InMux
    port map (
            O => \N__9651\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__2214\ : InMux
    port map (
            O => \N__9648\,
            I => \N__9644\
        );

    \I__2213\ : InMux
    port map (
            O => \N__9647\,
            I => \N__9641\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__9644\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__9641\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__2210\ : InMux
    port map (
            O => \N__9636\,
            I => \N__9632\
        );

    \I__2209\ : InMux
    port map (
            O => \N__9635\,
            I => \N__9629\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__9632\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__9629\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__9624\,
            I => \N__9621\
        );

    \I__2205\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9618\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__9618\,
            I => \N__9614\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9611\
        );

    \I__2202\ : Odrv12
    port map (
            O => \N__9614\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__9611\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__2200\ : InMux
    port map (
            O => \N__9606\,
            I => \N__9603\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__9603\,
            I => \U409_TICK.TICK603_11\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__9600\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__2197\ : IoInMux
    port map (
            O => \N__9597\,
            I => \N__9594\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__9594\,
            I => \N__9591\
        );

    \I__2195\ : Span4Mux_s3_v
    port map (
            O => \N__9591\,
            I => \N__9588\
        );

    \I__2194\ : Span4Mux_v
    port map (
            O => \N__9588\,
            I => \N__9585\
        );

    \I__2193\ : Span4Mux_v
    port map (
            O => \N__9585\,
            I => \N__9582\
        );

    \I__2192\ : Span4Mux_h
    port map (
            O => \N__9582\,
            I => \N__9578\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9575\
        );

    \I__2190\ : Odrv4
    port map (
            O => \N__9578\,
            I => \TICK60_c\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__9575\,
            I => \TICK60_c\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__9570\,
            I => \U409_CIA.CLK_CIA6_0_a2_0_cascade_\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__9567\,
            I => \U409_CIA.CLK_CIA6_cascade_\
        );

    \I__2186\ : IoInMux
    port map (
            O => \N__9564\,
            I => \N__9561\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__9561\,
            I => \N__9558\
        );

    \I__2184\ : IoSpan4Mux
    port map (
            O => \N__9558\,
            I => \N__9555\
        );

    \I__2183\ : Span4Mux_s2_v
    port map (
            O => \N__9555\,
            I => \N__9552\
        );

    \I__2182\ : Span4Mux_v
    port map (
            O => \N__9552\,
            I => \N__9549\
        );

    \I__2181\ : Sp12to4
    port map (
            O => \N__9549\,
            I => \N__9544\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9548\,
            I => \N__9541\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9547\,
            I => \N__9538\
        );

    \I__2178\ : Odrv12
    port map (
            O => \N__9544\,
            I => \CLK_CIA_c\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__9541\,
            I => \CLK_CIA_c\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9538\,
            I => \CLK_CIA_c\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__9531\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_3_0_a2_0_cascade_\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9525\,
            I => \N__9521\
        );

    \I__2172\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9518\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9521\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9518\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__2169\ : InMux
    port map (
            O => \N__9513\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9510\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9507\,
            I => \bfn_13_7_0_\
        );

    \I__2166\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9500\
        );

    \I__2165\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9497\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9500\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__9497\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9492\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9489\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__2160\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9482\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9485\,
            I => \N__9479\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__9482\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9479\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9474\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9471\,
            I => \N__9467\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9470\,
            I => \N__9464\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__9467\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__9464\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9459\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9456\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__9453\,
            I => \N__9449\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9452\,
            I => \N__9446\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9443\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__9446\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__9443\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9438\,
            I => \N__9435\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9435\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9432\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__2141\ : InMux
    port map (
            O => \N__9429\,
            I => \N__9426\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__9426\,
            I => \N__9421\
        );

    \I__2139\ : SRMux
    port map (
            O => \N__9425\,
            I => \N__9387\
        );

    \I__2138\ : SRMux
    port map (
            O => \N__9424\,
            I => \N__9387\
        );

    \I__2137\ : Glb2LocalMux
    port map (
            O => \N__9421\,
            I => \N__9387\
        );

    \I__2136\ : SRMux
    port map (
            O => \N__9420\,
            I => \N__9387\
        );

    \I__2135\ : SRMux
    port map (
            O => \N__9419\,
            I => \N__9387\
        );

    \I__2134\ : SRMux
    port map (
            O => \N__9418\,
            I => \N__9387\
        );

    \I__2133\ : SRMux
    port map (
            O => \N__9417\,
            I => \N__9387\
        );

    \I__2132\ : SRMux
    port map (
            O => \N__9416\,
            I => \N__9387\
        );

    \I__2131\ : SRMux
    port map (
            O => \N__9415\,
            I => \N__9387\
        );

    \I__2130\ : SRMux
    port map (
            O => \N__9414\,
            I => \N__9387\
        );

    \I__2129\ : SRMux
    port map (
            O => \N__9413\,
            I => \N__9387\
        );

    \I__2128\ : SRMux
    port map (
            O => \N__9412\,
            I => \N__9387\
        );

    \I__2127\ : GlobalMux
    port map (
            O => \N__9387\,
            I => \N__9384\
        );

    \I__2126\ : gio2CtrlBuf
    port map (
            O => \N__9384\,
            I => \RESETn_c_i_g\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9381\,
            I => \N__9377\
        );

    \I__2124\ : InMux
    port map (
            O => \N__9380\,
            I => \N__9374\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__9377\,
            I => \N__9369\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9374\,
            I => \N__9369\
        );

    \I__2121\ : Span4Mux_v
    port map (
            O => \N__9369\,
            I => \N__9366\
        );

    \I__2120\ : Span4Mux_h
    port map (
            O => \N__9366\,
            I => \N__9362\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9365\,
            I => \N__9359\
        );

    \I__2118\ : Sp12to4
    port map (
            O => \N__9362\,
            I => \N__9356\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9359\,
            I => \N__9353\
        );

    \I__2116\ : Span12Mux_h
    port map (
            O => \N__9356\,
            I => \N__9350\
        );

    \I__2115\ : Span12Mux_v
    port map (
            O => \N__9353\,
            I => \N__9347\
        );

    \I__2114\ : Span12Mux_v
    port map (
            O => \N__9350\,
            I => \N__9342\
        );

    \I__2113\ : Span12Mux_h
    port map (
            O => \N__9347\,
            I => \N__9342\
        );

    \I__2112\ : Odrv12
    port map (
            O => \N__9342\,
            I => \OVL_c\
        );

    \I__2111\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9336\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9336\,
            I => \N__9332\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__9335\,
            I => \N__9329\
        );

    \I__2108\ : Span4Mux_v
    port map (
            O => \N__9332\,
            I => \N__9325\
        );

    \I__2107\ : InMux
    port map (
            O => \N__9329\,
            I => \N__9322\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9319\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__9325\,
            I => \N_429\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9322\,
            I => \N_429\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__9319\,
            I => \N_429\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__9312\,
            I => \N__9309\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9309\,
            I => \N__9305\
        );

    \I__2100\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9298\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9305\,
            I => \N__9295\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9304\,
            I => \N__9290\
        );

    \I__2097\ : InMux
    port map (
            O => \N__9303\,
            I => \N__9290\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9302\,
            I => \N__9287\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9301\,
            I => \N__9284\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__9298\,
            I => \N__9281\
        );

    \I__2093\ : Span4Mux_h
    port map (
            O => \N__9295\,
            I => \N__9272\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__9290\,
            I => \N__9272\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__9287\,
            I => \N__9272\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9284\,
            I => \N__9272\
        );

    \I__2089\ : Span4Mux_v
    port map (
            O => \N__9281\,
            I => \N__9267\
        );

    \I__2088\ : Span4Mux_v
    port map (
            O => \N__9272\,
            I => \N__9264\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9271\,
            I => \N__9261\
        );

    \I__2086\ : InMux
    port map (
            O => \N__9270\,
            I => \N__9258\
        );

    \I__2085\ : Odrv4
    port map (
            O => \N__9267\,
            I => \N_348\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__9264\,
            I => \N_348\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__9261\,
            I => \N_348\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__9258\,
            I => \N_348\
        );

    \I__2081\ : CascadeMux
    port map (
            O => \N__9249\,
            I => \N__9243\
        );

    \I__2080\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9240\
        );

    \I__2079\ : InMux
    port map (
            O => \N__9247\,
            I => \N__9237\
        );

    \I__2078\ : InMux
    port map (
            O => \N__9246\,
            I => \N__9231\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9243\,
            I => \N__9231\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9240\,
            I => \N__9227\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__9237\,
            I => \N__9224\
        );

    \I__2074\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9221\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__9231\,
            I => \N__9218\
        );

    \I__2072\ : InMux
    port map (
            O => \N__9230\,
            I => \N__9215\
        );

    \I__2071\ : Span4Mux_h
    port map (
            O => \N__9227\,
            I => \N__9208\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__9224\,
            I => \N__9208\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__9221\,
            I => \N__9208\
        );

    \I__2068\ : Span12Mux_v
    port map (
            O => \N__9218\,
            I => \N__9205\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__9215\,
            I => \N__9202\
        );

    \I__2066\ : Span4Mux_v
    port map (
            O => \N__9208\,
            I => \N__9199\
        );

    \I__2065\ : Odrv12
    port map (
            O => \N__9205\,
            I => \N_156_i\
        );

    \I__2064\ : Odrv12
    port map (
            O => \N__9202\,
            I => \N_156_i\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__9199\,
            I => \N_156_i\
        );

    \I__2062\ : IoInMux
    port map (
            O => \N__9192\,
            I => \N__9189\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__9189\,
            I => \N__9186\
        );

    \I__2060\ : Span12Mux_s11_v
    port map (
            O => \N__9186\,
            I => \N__9183\
        );

    \I__2059\ : Odrv12
    port map (
            O => \N__9183\,
            I => \N_264_i\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9174\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__9179\,
            I => \N__9171\
        );

    \I__2056\ : CascadeMux
    port map (
            O => \N__9178\,
            I => \N__9164\
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__9177\,
            I => \N__9160\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__9174\,
            I => \N__9155\
        );

    \I__2053\ : InMux
    port map (
            O => \N__9171\,
            I => \N__9152\
        );

    \I__2052\ : InMux
    port map (
            O => \N__9170\,
            I => \N__9149\
        );

    \I__2051\ : InMux
    port map (
            O => \N__9169\,
            I => \N__9146\
        );

    \I__2050\ : InMux
    port map (
            O => \N__9168\,
            I => \N__9137\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9167\,
            I => \N__9137\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9137\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9137\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9160\,
            I => \N__9132\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9159\,
            I => \N__9127\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9127\
        );

    \I__2043\ : Span4Mux_h
    port map (
            O => \N__9155\,
            I => \N__9122\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9152\,
            I => \N__9122\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__9149\,
            I => \N__9119\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__9146\,
            I => \N__9114\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__9137\,
            I => \N__9114\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9111\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9108\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9132\,
            I => \N__9100\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__9127\,
            I => \N__9100\
        );

    \I__2034\ : Span4Mux_v
    port map (
            O => \N__9122\,
            I => \N__9090\
        );

    \I__2033\ : Span4Mux_h
    port map (
            O => \N__9119\,
            I => \N__9090\
        );

    \I__2032\ : Span4Mux_h
    port map (
            O => \N__9114\,
            I => \N__9090\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9111\,
            I => \N__9090\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9108\,
            I => \N__9087\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9107\,
            I => \N__9084\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9106\,
            I => \N__9079\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9105\,
            I => \N__9079\
        );

    \I__2026\ : Span4Mux_h
    port map (
            O => \N__9100\,
            I => \N__9076\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9073\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__9090\,
            I => \N__9067\
        );

    \I__2023\ : Span4Mux_h
    port map (
            O => \N__9087\,
            I => \N__9062\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__9084\,
            I => \N__9062\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9079\,
            I => \N__9059\
        );

    \I__2020\ : Span4Mux_h
    port map (
            O => \N__9076\,
            I => \N__9056\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__9073\,
            I => \N__9053\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9072\,
            I => \N__9050\
        );

    \I__2017\ : InMux
    port map (
            O => \N__9071\,
            I => \N__9045\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9070\,
            I => \N__9045\
        );

    \I__2015\ : Span4Mux_h
    port map (
            O => \N__9067\,
            I => \N__9037\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__9062\,
            I => \N__9037\
        );

    \I__2013\ : Span4Mux_v
    port map (
            O => \N__9059\,
            I => \N__9037\
        );

    \I__2012\ : Sp12to4
    port map (
            O => \N__9056\,
            I => \N__9028\
        );

    \I__2011\ : Span12Mux_s7_v
    port map (
            O => \N__9053\,
            I => \N__9028\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__9050\,
            I => \N__9028\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__9045\,
            I => \N__9028\
        );

    \I__2008\ : InMux
    port map (
            O => \N__9044\,
            I => \N__9025\
        );

    \I__2007\ : Sp12to4
    port map (
            O => \N__9037\,
            I => \N__9018\
        );

    \I__2006\ : Span12Mux_v
    port map (
            O => \N__9028\,
            I => \N__9018\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__9025\,
            I => \N__9018\
        );

    \I__2004\ : Span12Mux_v
    port map (
            O => \N__9018\,
            I => \N__9015\
        );

    \I__2003\ : Span12Mux_h
    port map (
            O => \N__9015\,
            I => \N__9012\
        );

    \I__2002\ : Odrv12
    port map (
            O => \N__9012\,
            I => \RESETn_c\
        );

    \I__2001\ : IoInMux
    port map (
            O => \N__9009\,
            I => \N__9006\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9006\,
            I => \N__9003\
        );

    \I__1999\ : Odrv12
    port map (
            O => \N__9003\,
            I => \RESETn_c_i\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__9000\,
            I => \N__8996\
        );

    \I__1997\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8991\
        );

    \I__1996\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8991\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__8991\,
            I => \N__8987\
        );

    \I__1994\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8984\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__8987\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__8984\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1991\ : InMux
    port map (
            O => \N__8979\,
            I => \N__8975\
        );

    \I__1990\ : InMux
    port map (
            O => \N__8978\,
            I => \N__8972\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__8975\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__8972\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1987\ : InMux
    port map (
            O => \N__8967\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__1986\ : InMux
    port map (
            O => \N__8964\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__1985\ : InMux
    port map (
            O => \N__8961\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__1984\ : InMux
    port map (
            O => \N__8958\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__8955\,
            I => \N__8952\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8952\,
            I => \N__8949\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__8949\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__1980\ : InMux
    port map (
            O => \N__8946\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__8943\,
            I => \U409_TRANSFER_ACK.m12_i_0_cascade_\
        );

    \I__1978\ : InMux
    port map (
            O => \N__8940\,
            I => \N__8937\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__8937\,
            I => \U409_TRANSFER_ACK.N_293\
        );

    \I__1976\ : InMux
    port map (
            O => \N__8934\,
            I => \N__8931\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__8931\,
            I => \U409_TRANSFER_ACK.N_191\
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__8928\,
            I => \U409_TRANSFER_ACK.N_191_cascade_\
        );

    \I__1973\ : InMux
    port map (
            O => \N__8925\,
            I => \N__8922\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__8922\,
            I => \U409_TRANSFER_ACK.N_223\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__8919\,
            I => \U409_TRANSFER_ACK.i5_mux_cascade_\
        );

    \I__1970\ : InMux
    port map (
            O => \N__8916\,
            I => \N__8913\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__8913\,
            I => \N__8905\
        );

    \I__1968\ : InMux
    port map (
            O => \N__8912\,
            I => \N__8900\
        );

    \I__1967\ : InMux
    port map (
            O => \N__8911\,
            I => \N__8900\
        );

    \I__1966\ : InMux
    port map (
            O => \N__8910\,
            I => \N__8897\
        );

    \I__1965\ : InMux
    port map (
            O => \N__8909\,
            I => \N__8892\
        );

    \I__1964\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8892\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__8905\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__8900\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__8897\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__8892\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__8883\,
            I => \N__8880\
        );

    \I__1958\ : InMux
    port map (
            O => \N__8880\,
            I => \N__8877\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__8877\,
            I => \N__8870\
        );

    \I__1956\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8863\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8875\,
            I => \N__8863\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8863\
        );

    \I__1953\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8860\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__8870\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__8863\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__8860\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1949\ : InMux
    port map (
            O => \N__8853\,
            I => \N__8850\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__8850\,
            I => \U409_TRANSFER_ACK.N_290\
        );

    \I__1947\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8841\
        );

    \I__1946\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8834\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8834\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8844\,
            I => \N__8834\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__8841\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__8834\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__8829\,
            I => \N__8825\
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__8828\,
            I => \N__8822\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8814\
        );

    \I__1938\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8814\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8821\,
            I => \N__8814\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8814\,
            I => \N__8811\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__8811\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__1934\ : InMux
    port map (
            O => \N__8808\,
            I => \N__8802\
        );

    \I__1933\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8797\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8806\,
            I => \N__8797\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8805\,
            I => \N__8794\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__8802\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__8797\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__8794\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1927\ : InMux
    port map (
            O => \N__8787\,
            I => \N__8780\
        );

    \I__1926\ : InMux
    port map (
            O => \N__8786\,
            I => \N__8780\
        );

    \I__1925\ : InMux
    port map (
            O => \N__8785\,
            I => \N__8777\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8780\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__8777\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__8772\,
            I => \CIA_ENABLE_cascade_\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8766\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__8766\,
            I => \N__8763\
        );

    \I__1919\ : Span12Mux_h
    port map (
            O => \N__8763\,
            I => \N__8760\
        );

    \I__1918\ : Odrv12
    port map (
            O => \N__8760\,
            I => \A_c_12\
        );

    \I__1917\ : IoInMux
    port map (
            O => \N__8757\,
            I => \N__8754\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__8754\,
            I => \N__8751\
        );

    \I__1915\ : Span4Mux_s0_h
    port map (
            O => \N__8751\,
            I => \N__8748\
        );

    \I__1914\ : Span4Mux_h
    port map (
            O => \N__8748\,
            I => \N__8745\
        );

    \I__1913\ : Sp12to4
    port map (
            O => \N__8745\,
            I => \N__8742\
        );

    \I__1912\ : Span12Mux_s8_v
    port map (
            O => \N__8742\,
            I => \N__8739\
        );

    \I__1911\ : Span12Mux_h
    port map (
            O => \N__8739\,
            I => \N__8736\
        );

    \I__1910\ : Odrv12
    port map (
            O => \N__8736\,
            I => \U409_ADDRESS_DECODE_un1_CIACS0n_i\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__8733\,
            I => \U409_TICK.TICK603_10_cascade_\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__8730\,
            I => \U409_TRANSFER_ACK.m12_i_a2_1_0_cascade_\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__8727\,
            I => \N__8724\
        );

    \I__1906\ : InMux
    port map (
            O => \N__8724\,
            I => \N__8721\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__8721\,
            I => \U409_TRANSFER_ACK.N_379\
        );

    \I__1904\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8715\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__8715\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8712\,
            I => \N__8709\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__8709\,
            I => \U409_TRANSFER_ACK.N_307\
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__8706\,
            I => \N__8703\
        );

    \I__1899\ : InMux
    port map (
            O => \N__8703\,
            I => \N__8699\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8695\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__8699\,
            I => \N__8692\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8698\,
            I => \N__8689\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__8695\,
            I => \N__8686\
        );

    \I__1894\ : Span4Mux_v
    port map (
            O => \N__8692\,
            I => \N__8681\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__8689\,
            I => \N__8681\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__8686\,
            I => \U409_TRANSFER_ACK.N_381\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__8681\,
            I => \U409_TRANSFER_ACK.N_381\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8673\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__8673\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0\
        );

    \I__1888\ : InMux
    port map (
            O => \N__8670\,
            I => \N__8667\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8667\,
            I => \U409_TRANSFER_ACK.ROMENn_e_1\
        );

    \I__1886\ : IoInMux
    port map (
            O => \N__8664\,
            I => \N__8661\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8661\,
            I => \N__8658\
        );

    \I__1884\ : Span4Mux_s2_v
    port map (
            O => \N__8658\,
            I => \N__8655\
        );

    \I__1883\ : Sp12to4
    port map (
            O => \N__8655\,
            I => \N__8652\
        );

    \I__1882\ : Span12Mux_h
    port map (
            O => \N__8652\,
            I => \N__8648\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__8651\,
            I => \N__8645\
        );

    \I__1880\ : Span12Mux_v
    port map (
            O => \N__8648\,
            I => \N__8642\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8639\
        );

    \I__1878\ : Odrv12
    port map (
            O => \N__8642\,
            I => \ROMENn_c\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8639\,
            I => \ROMENn_c\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__8634\,
            I => \N__8627\
        );

    \I__1875\ : InMux
    port map (
            O => \N__8633\,
            I => \N__8620\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8632\,
            I => \N__8620\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8631\,
            I => \N__8617\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8630\,
            I => \N__8614\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8627\,
            I => \N__8611\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8626\,
            I => \N__8608\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8605\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8620\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8617\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__8614\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8611\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8608\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__8605\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__8592\,
            I => \N__8587\
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__8591\,
            I => \N__8582\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8578\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8587\,
            I => \N__8575\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8586\,
            I => \N__8572\
        );

    \I__1857\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8569\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8564\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8564\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8578\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8575\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__8572\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__8569\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8564\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__8553\,
            I => \N__8548\
        );

    \I__1848\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8540\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8540\
        );

    \I__1846\ : InMux
    port map (
            O => \N__8548\,
            I => \N__8535\
        );

    \I__1845\ : InMux
    port map (
            O => \N__8547\,
            I => \N__8535\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8546\,
            I => \N__8532\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8545\,
            I => \N__8529\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__8540\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8535\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8532\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8529\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8520\,
            I => \N__8512\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8507\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8518\,
            I => \N__8507\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8504\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8499\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8515\,
            I => \N__8499\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8512\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__8507\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8504\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__8499\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1828\ : IoInMux
    port map (
            O => \N__8490\,
            I => \N__8487\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8487\,
            I => \N__8483\
        );

    \I__1826\ : IoInMux
    port map (
            O => \N__8486\,
            I => \N__8480\
        );

    \I__1825\ : IoSpan4Mux
    port map (
            O => \N__8483\,
            I => \N__8477\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__8480\,
            I => \N__8474\
        );

    \I__1823\ : Span4Mux_s2_v
    port map (
            O => \N__8477\,
            I => \N__8469\
        );

    \I__1822\ : Span4Mux_s2_v
    port map (
            O => \N__8474\,
            I => \N__8469\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__8469\,
            I => \N__8466\
        );

    \I__1820\ : Sp12to4
    port map (
            O => \N__8466\,
            I => \N__8461\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8458\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__8464\,
            I => \N__8455\
        );

    \I__1817\ : Span12Mux_h
    port map (
            O => \N__8461\,
            I => \N__8450\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8458\,
            I => \N__8450\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8447\
        );

    \I__1814\ : Odrv12
    port map (
            O => \N__8450\,
            I => \TACK_EN\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8447\,
            I => \TACK_EN\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8442\,
            I => \N__8439\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8439\,
            I => \N__8435\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8432\
        );

    \I__1809\ : Span4Mux_v
    port map (
            O => \N__8435\,
            I => \N__8429\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8432\,
            I => \N__8426\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__8429\,
            I => \N_357\
        );

    \I__1806\ : Odrv4
    port map (
            O => \N__8426\,
            I => \N_357\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8418\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__8418\,
            I => \N__8414\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8411\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__8414\,
            I => \N_339\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8411\,
            I => \N_339\
        );

    \I__1800\ : IoInMux
    port map (
            O => \N__8406\,
            I => \N__8403\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8403\,
            I => \N__8400\
        );

    \I__1798\ : IoSpan4Mux
    port map (
            O => \N__8400\,
            I => \N__8397\
        );

    \I__1797\ : IoSpan4Mux
    port map (
            O => \N__8397\,
            I => \N__8394\
        );

    \I__1796\ : Sp12to4
    port map (
            O => \N__8394\,
            I => \N__8391\
        );

    \I__1795\ : Span12Mux_v
    port map (
            O => \N__8391\,
            I => \N__8388\
        );

    \I__1794\ : Odrv12
    port map (
            O => \N__8388\,
            I => \TCIn_1_i\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__8385\,
            I => \N__8377\
        );

    \I__1792\ : CascadeMux
    port map (
            O => \N__8384\,
            I => \N__8374\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8383\,
            I => \N__8370\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8382\,
            I => \N__8365\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8381\,
            I => \N__8365\
        );

    \I__1788\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8362\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8359\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8354\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8373\,
            I => \N__8354\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8370\,
            I => \N__8351\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8365\,
            I => \N__8339\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8362\,
            I => \N__8336\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__8359\,
            I => \N__8333\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8354\,
            I => \N__8330\
        );

    \I__1779\ : Glb2LocalMux
    port map (
            O => \N__8351\,
            I => \N__8298\
        );

    \I__1778\ : ClkMux
    port map (
            O => \N__8350\,
            I => \N__8298\
        );

    \I__1777\ : ClkMux
    port map (
            O => \N__8349\,
            I => \N__8298\
        );

    \I__1776\ : ClkMux
    port map (
            O => \N__8348\,
            I => \N__8298\
        );

    \I__1775\ : ClkMux
    port map (
            O => \N__8347\,
            I => \N__8298\
        );

    \I__1774\ : ClkMux
    port map (
            O => \N__8346\,
            I => \N__8298\
        );

    \I__1773\ : ClkMux
    port map (
            O => \N__8345\,
            I => \N__8298\
        );

    \I__1772\ : ClkMux
    port map (
            O => \N__8344\,
            I => \N__8298\
        );

    \I__1771\ : ClkMux
    port map (
            O => \N__8343\,
            I => \N__8298\
        );

    \I__1770\ : ClkMux
    port map (
            O => \N__8342\,
            I => \N__8298\
        );

    \I__1769\ : Glb2LocalMux
    port map (
            O => \N__8339\,
            I => \N__8298\
        );

    \I__1768\ : Glb2LocalMux
    port map (
            O => \N__8336\,
            I => \N__8298\
        );

    \I__1767\ : Glb2LocalMux
    port map (
            O => \N__8333\,
            I => \N__8298\
        );

    \I__1766\ : Glb2LocalMux
    port map (
            O => \N__8330\,
            I => \N__8298\
        );

    \I__1765\ : ClkMux
    port map (
            O => \N__8329\,
            I => \N__8298\
        );

    \I__1764\ : GlobalMux
    port map (
            O => \N__8298\,
            I => \N__8295\
        );

    \I__1763\ : gio2CtrlBuf
    port map (
            O => \N__8295\,
            I => \CLK40_IN_c_g\
        );

    \I__1762\ : IoInMux
    port map (
            O => \N__8292\,
            I => \N__8289\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8289\,
            I => \N__8286\
        );

    \I__1760\ : Span4Mux_s2_v
    port map (
            O => \N__8286\,
            I => \N__8283\
        );

    \I__1759\ : Span4Mux_v
    port map (
            O => \N__8283\,
            I => \N__8280\
        );

    \I__1758\ : Odrv4
    port map (
            O => \N__8280\,
            I => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\
        );

    \I__1757\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8274\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8274\,
            I => \CIA_ENABLE\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__8271\,
            I => \U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8268\,
            I => \N__8265\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__8265\,
            I => \U409_TRANSFER_ACK.N_289\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__8262\,
            I => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\
        );

    \I__1751\ : IoInMux
    port map (
            O => \N__8259\,
            I => \N__8255\
        );

    \I__1750\ : IoInMux
    port map (
            O => \N__8258\,
            I => \N__8252\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__8255\,
            I => \N__8247\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8252\,
            I => \N__8247\
        );

    \I__1747\ : IoSpan4Mux
    port map (
            O => \N__8247\,
            I => \N__8243\
        );

    \I__1746\ : IoInMux
    port map (
            O => \N__8246\,
            I => \N__8240\
        );

    \I__1745\ : Span4Mux_s1_v
    port map (
            O => \N__8243\,
            I => \N__8237\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__8240\,
            I => \N__8234\
        );

    \I__1743\ : Span4Mux_v
    port map (
            O => \N__8237\,
            I => \N__8229\
        );

    \I__1742\ : Span4Mux_s1_v
    port map (
            O => \N__8234\,
            I => \N__8229\
        );

    \I__1741\ : Sp12to4
    port map (
            O => \N__8229\,
            I => \N__8226\
        );

    \I__1740\ : Span12Mux_h
    port map (
            O => \N__8226\,
            I => \N__8223\
        );

    \I__1739\ : Span12Mux_v
    port map (
            O => \N__8223\,
            I => \N__8218\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8222\,
            I => \N__8213\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8221\,
            I => \N__8213\
        );

    \I__1736\ : Odrv12
    port map (
            O => \N__8218\,
            I => \TACK_OUTn\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8213\,
            I => \TACK_OUTn\
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__8208\,
            I => \N__8202\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__8207\,
            I => \N__8199\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__8206\,
            I => \N__8196\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8193\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8202\,
            I => \N__8186\
        );

    \I__1729\ : InMux
    port map (
            O => \N__8199\,
            I => \N__8186\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8196\,
            I => \N__8186\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__8193\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__8186\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8181\,
            I => \N__8175\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8180\,
            I => \N__8168\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8179\,
            I => \N__8168\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8178\,
            I => \N__8168\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__8175\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8168\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8158\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8162\,
            I => \N__8153\
        );

    \I__1717\ : InMux
    port map (
            O => \N__8161\,
            I => \N__8153\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__8158\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8153\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1714\ : InMux
    port map (
            O => \N__8148\,
            I => \N__8145\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__8145\,
            I => \N__8141\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8144\,
            I => \N__8138\
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__8141\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__8138\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__1709\ : CascadeMux
    port map (
            O => \N__8133\,
            I => \N__8130\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8130\,
            I => \N__8126\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__8129\,
            I => \N__8123\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8126\,
            I => \N__8120\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8123\,
            I => \N__8117\
        );

    \I__1704\ : Span4Mux_h
    port map (
            O => \N__8120\,
            I => \N__8112\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__8117\,
            I => \N__8112\
        );

    \I__1702\ : Span4Mux_h
    port map (
            O => \N__8112\,
            I => \N__8109\
        );

    \I__1701\ : Odrv4
    port map (
            O => \N__8109\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz\
        );

    \I__1700\ : InMux
    port map (
            O => \N__8106\,
            I => \N__8102\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8105\,
            I => \N__8099\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__8102\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__8099\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__8094\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\
        );

    \I__1695\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8087\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8090\,
            I => \N__8084\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8087\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__8084\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8079\,
            I => \N__8075\
        );

    \I__1690\ : InMux
    port map (
            O => \N__8078\,
            I => \N__8072\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__8075\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8072\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8067\,
            I => \N__8061\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8066\,
            I => \N__8061\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8061\,
            I => \U409_TRANSFER_ACK.N_159\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8058\,
            I => \N__8055\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8055\,
            I => \U409_TRANSFER_ACK.N_380\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__8052\,
            I => \U409_TRANSFER_ACK.N_380_cascade_\
        );

    \I__1681\ : InMux
    port map (
            O => \N__8049\,
            I => \N__8046\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__8046\,
            I => \N_190\
        );

    \I__1679\ : InMux
    port map (
            O => \N__8043\,
            I => \N__8040\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__8040\,
            I => \N__8036\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8039\,
            I => \N__8033\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__8036\,
            I => \N__8030\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__8033\,
            I => \N__8027\
        );

    \I__1674\ : Odrv4
    port map (
            O => \N__8030\,
            I => \N_297\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__8027\,
            I => \N_297\
        );

    \I__1672\ : IoInMux
    port map (
            O => \N__8022\,
            I => \N__8019\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__8019\,
            I => \N__8016\
        );

    \I__1670\ : Span12Mux_s7_v
    port map (
            O => \N__8016\,
            I => \N__8013\
        );

    \I__1669\ : Span12Mux_h
    port map (
            O => \N__8013\,
            I => \N__8010\
        );

    \I__1668\ : Odrv12
    port map (
            O => \N__8010\,
            I => \N_94_i\
        );

    \I__1667\ : InMux
    port map (
            O => \N__8007\,
            I => \N__8004\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__8004\,
            I => \N__8001\
        );

    \I__1665\ : Span4Mux_v
    port map (
            O => \N__8001\,
            I => \N__7998\
        );

    \I__1664\ : Sp12to4
    port map (
            O => \N__7998\,
            I => \N__7995\
        );

    \I__1663\ : Span12Mux_h
    port map (
            O => \N__7995\,
            I => \N__7992\
        );

    \I__1662\ : Odrv12
    port map (
            O => \N__7992\,
            I => \A_c_13\
        );

    \I__1661\ : IoInMux
    port map (
            O => \N__7989\,
            I => \N__7986\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7986\,
            I => \N__7983\
        );

    \I__1659\ : Span4Mux_s1_h
    port map (
            O => \N__7983\,
            I => \N__7980\
        );

    \I__1658\ : Sp12to4
    port map (
            O => \N__7980\,
            I => \N__7977\
        );

    \I__1657\ : Span12Mux_s9_v
    port map (
            O => \N__7977\,
            I => \N__7974\
        );

    \I__1656\ : Span12Mux_h
    port map (
            O => \N__7974\,
            I => \N__7971\
        );

    \I__1655\ : Odrv12
    port map (
            O => \N__7971\,
            I => \U409_ADDRESS_DECODE_un1_CIACS1n_i\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7968\,
            I => \N__7965\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__7965\,
            I => \N__7959\
        );

    \I__1652\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7956\
        );

    \I__1651\ : InMux
    port map (
            O => \N__7963\,
            I => \N__7953\
        );

    \I__1650\ : InMux
    port map (
            O => \N__7962\,
            I => \N__7949\
        );

    \I__1649\ : Span4Mux_v
    port map (
            O => \N__7959\,
            I => \N__7944\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__7956\,
            I => \N__7944\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__7953\,
            I => \N__7941\
        );

    \I__1646\ : InMux
    port map (
            O => \N__7952\,
            I => \N__7938\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__7949\,
            I => \N__7933\
        );

    \I__1644\ : Span4Mux_v
    port map (
            O => \N__7944\,
            I => \N__7926\
        );

    \I__1643\ : Span4Mux_h
    port map (
            O => \N__7941\,
            I => \N__7926\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__7938\,
            I => \N__7926\
        );

    \I__1641\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7923\
        );

    \I__1640\ : InMux
    port map (
            O => \N__7936\,
            I => \N__7920\
        );

    \I__1639\ : Span4Mux_v
    port map (
            O => \N__7933\,
            I => \N__7917\
        );

    \I__1638\ : Span4Mux_h
    port map (
            O => \N__7926\,
            I => \N__7912\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__7923\,
            I => \N__7912\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__7920\,
            I => \N__7909\
        );

    \I__1635\ : Span4Mux_v
    port map (
            O => \N__7917\,
            I => \N__7906\
        );

    \I__1634\ : Span4Mux_v
    port map (
            O => \N__7912\,
            I => \N__7903\
        );

    \I__1633\ : Span12Mux_h
    port map (
            O => \N__7909\,
            I => \N__7900\
        );

    \I__1632\ : Span4Mux_v
    port map (
            O => \N__7906\,
            I => \N__7897\
        );

    \I__1631\ : Span4Mux_v
    port map (
            O => \N__7903\,
            I => \N__7894\
        );

    \I__1630\ : Span12Mux_v
    port map (
            O => \N__7900\,
            I => \N__7891\
        );

    \I__1629\ : Sp12to4
    port map (
            O => \N__7897\,
            I => \N__7886\
        );

    \I__1628\ : Sp12to4
    port map (
            O => \N__7894\,
            I => \N__7886\
        );

    \I__1627\ : Odrv12
    port map (
            O => \N__7891\,
            I => \A_c_22\
        );

    \I__1626\ : Odrv12
    port map (
            O => \N__7886\,
            I => \A_c_22\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__7881\,
            I => \N__7878\
        );

    \I__1624\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7875\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7875\,
            I => \N__7871\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__7874\,
            I => \N__7867\
        );

    \I__1621\ : Span4Mux_v
    port map (
            O => \N__7871\,
            I => \N__7864\
        );

    \I__1620\ : InMux
    port map (
            O => \N__7870\,
            I => \N__7861\
        );

    \I__1619\ : InMux
    port map (
            O => \N__7867\,
            I => \N__7858\
        );

    \I__1618\ : Sp12to4
    port map (
            O => \N__7864\,
            I => \N__7850\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__7861\,
            I => \N__7850\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__7858\,
            I => \N__7850\
        );

    \I__1615\ : InMux
    port map (
            O => \N__7857\,
            I => \N__7847\
        );

    \I__1614\ : Odrv12
    port map (
            O => \N__7850\,
            I => \N_401\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__7847\,
            I => \N_401\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__7842\,
            I => \N_431_cascade_\
        );

    \I__1611\ : InMux
    port map (
            O => \N__7839\,
            I => \N__7836\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__7836\,
            I => \N__7832\
        );

    \I__1609\ : InMux
    port map (
            O => \N__7835\,
            I => \N__7829\
        );

    \I__1608\ : Span4Mux_h
    port map (
            O => \N__7832\,
            I => \N__7823\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__7829\,
            I => \N__7823\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7828\,
            I => \N__7820\
        );

    \I__1605\ : Sp12to4
    port map (
            O => \N__7823\,
            I => \N__7815\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__7820\,
            I => \N__7815\
        );

    \I__1603\ : Odrv12
    port map (
            O => \N__7815\,
            I => \N_422\
        );

    \I__1602\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7808\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7805\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7808\,
            I => \N__7797\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__7805\,
            I => \N__7797\
        );

    \I__1598\ : InMux
    port map (
            O => \N__7804\,
            I => \N__7794\
        );

    \I__1597\ : InMux
    port map (
            O => \N__7803\,
            I => \N__7791\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7802\,
            I => \N__7788\
        );

    \I__1595\ : Span4Mux_v
    port map (
            O => \N__7797\,
            I => \N__7784\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__7794\,
            I => \N__7781\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__7791\,
            I => \N__7778\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__7788\,
            I => \N__7775\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7787\,
            I => \N__7772\
        );

    \I__1590\ : Span4Mux_h
    port map (
            O => \N__7784\,
            I => \N__7767\
        );

    \I__1589\ : Span4Mux_v
    port map (
            O => \N__7781\,
            I => \N__7767\
        );

    \I__1588\ : Span4Mux_v
    port map (
            O => \N__7778\,
            I => \N__7764\
        );

    \I__1587\ : Span4Mux_v
    port map (
            O => \N__7775\,
            I => \N__7759\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__7772\,
            I => \N__7759\
        );

    \I__1585\ : Span4Mux_v
    port map (
            O => \N__7767\,
            I => \N__7756\
        );

    \I__1584\ : Span4Mux_h
    port map (
            O => \N__7764\,
            I => \N__7751\
        );

    \I__1583\ : Span4Mux_v
    port map (
            O => \N__7759\,
            I => \N__7751\
        );

    \I__1582\ : Sp12to4
    port map (
            O => \N__7756\,
            I => \N__7746\
        );

    \I__1581\ : Sp12to4
    port map (
            O => \N__7751\,
            I => \N__7746\
        );

    \I__1580\ : Span12Mux_h
    port map (
            O => \N__7746\,
            I => \N__7743\
        );

    \I__1579\ : Span12Mux_v
    port map (
            O => \N__7743\,
            I => \N__7740\
        );

    \I__1578\ : Odrv12
    port map (
            O => \N__7740\,
            I => \A_c_19\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7737\,
            I => \N__7733\
        );

    \I__1576\ : InMux
    port map (
            O => \N__7736\,
            I => \N__7730\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7733\,
            I => \ATA_BASE_7\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__7730\,
            I => \ATA_BASE_7\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__7725\,
            I => \N__7722\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7722\,
            I => \N__7719\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__7719\,
            I => \N__7715\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7718\,
            I => \N__7712\
        );

    \I__1569\ : Span4Mux_v
    port map (
            O => \N__7715\,
            I => \N__7708\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7712\,
            I => \N__7705\
        );

    \I__1567\ : InMux
    port map (
            O => \N__7711\,
            I => \N__7702\
        );

    \I__1566\ : Span4Mux_v
    port map (
            O => \N__7708\,
            I => \N__7696\
        );

    \I__1565\ : Span4Mux_h
    port map (
            O => \N__7705\,
            I => \N__7691\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__7702\,
            I => \N__7691\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7701\,
            I => \N__7688\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__7700\,
            I => \N__7685\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__7699\,
            I => \N__7682\
        );

    \I__1560\ : Span4Mux_h
    port map (
            O => \N__7696\,
            I => \N__7679\
        );

    \I__1559\ : Span4Mux_v
    port map (
            O => \N__7691\,
            I => \N__7676\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7688\,
            I => \N__7673\
        );

    \I__1557\ : InMux
    port map (
            O => \N__7685\,
            I => \N__7668\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7668\
        );

    \I__1555\ : Sp12to4
    port map (
            O => \N__7679\,
            I => \N__7659\
        );

    \I__1554\ : Sp12to4
    port map (
            O => \N__7676\,
            I => \N__7659\
        );

    \I__1553\ : Span12Mux_h
    port map (
            O => \N__7673\,
            I => \N__7659\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7668\,
            I => \N__7659\
        );

    \I__1551\ : Odrv12
    port map (
            O => \N__7659\,
            I => \A_c_23\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7656\,
            I => \N__7650\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7655\,
            I => \N__7650\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7650\,
            I => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_5\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__7647\,
            I => \N__7640\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7646\,
            I => \N__7629\
        );

    \I__1545\ : InMux
    port map (
            O => \N__7645\,
            I => \N__7629\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7644\,
            I => \N__7629\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7643\,
            I => \N__7629\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7626\
        );

    \I__1541\ : CascadeMux
    port map (
            O => \N__7639\,
            I => \N__7620\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__7638\,
            I => \N__7615\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__7629\,
            I => \N__7612\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7626\,
            I => \N__7609\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7625\,
            I => \N__7594\
        );

    \I__1536\ : InMux
    port map (
            O => \N__7624\,
            I => \N__7594\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7623\,
            I => \N__7594\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7620\,
            I => \N__7594\
        );

    \I__1533\ : InMux
    port map (
            O => \N__7619\,
            I => \N__7594\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7618\,
            I => \N__7594\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7615\,
            I => \N__7594\
        );

    \I__1530\ : Span4Mux_v
    port map (
            O => \N__7612\,
            I => \N__7591\
        );

    \I__1529\ : Span4Mux_v
    port map (
            O => \N__7609\,
            I => \N__7588\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7594\,
            I => \N__7585\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__7591\,
            I => \N_361\
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__7588\,
            I => \N_361\
        );

    \I__1525\ : Odrv12
    port map (
            O => \N__7585\,
            I => \N_361\
        );

    \I__1524\ : CascadeMux
    port map (
            O => \N__7578\,
            I => \N__7574\
        );

    \I__1523\ : CascadeMux
    port map (
            O => \N__7577\,
            I => \N__7571\
        );

    \I__1522\ : InMux
    port map (
            O => \N__7574\,
            I => \N__7568\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7565\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7568\,
            I => \N__7562\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7565\,
            I => \N__7559\
        );

    \I__1518\ : Span4Mux_v
    port map (
            O => \N__7562\,
            I => \N__7555\
        );

    \I__1517\ : Span4Mux_v
    port map (
            O => \N__7559\,
            I => \N__7552\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7558\,
            I => \N__7549\
        );

    \I__1515\ : Span4Mux_h
    port map (
            O => \N__7555\,
            I => \N__7546\
        );

    \I__1514\ : Span4Mux_v
    port map (
            O => \N__7552\,
            I => \N__7543\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7549\,
            I => \N__7540\
        );

    \I__1512\ : Sp12to4
    port map (
            O => \N__7546\,
            I => \N__7535\
        );

    \I__1511\ : Sp12to4
    port map (
            O => \N__7543\,
            I => \N__7535\
        );

    \I__1510\ : Span4Mux_v
    port map (
            O => \N__7540\,
            I => \N__7532\
        );

    \I__1509\ : Span12Mux_h
    port map (
            O => \N__7535\,
            I => \N__7527\
        );

    \I__1508\ : Sp12to4
    port map (
            O => \N__7532\,
            I => \N__7527\
        );

    \I__1507\ : Odrv12
    port map (
            O => \N__7527\,
            I => \D_in_7\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7518\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7518\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7518\,
            I => \ATA_BASE_3\
        );

    \I__1503\ : CEMux
    port map (
            O => \N__7515\,
            I => \N__7512\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7512\,
            I => \N__7509\
        );

    \I__1501\ : Span4Mux_h
    port map (
            O => \N__7509\,
            I => \N__7506\
        );

    \I__1500\ : Span4Mux_h
    port map (
            O => \N__7506\,
            I => \N__7502\
        );

    \I__1499\ : CEMux
    port map (
            O => \N__7505\,
            I => \N__7499\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__7502\,
            I => \U409_AUTOCONFIG.un1_STATE_1_0_0\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7499\,
            I => \U409_AUTOCONFIG.un1_STATE_1_0_0\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7494\,
            I => \N__7482\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7493\,
            I => \N__7482\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7492\,
            I => \N__7482\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7491\,
            I => \N__7482\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7482\,
            I => \U409_AUTOCONFIG.N_172\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__7479\,
            I => \N__7476\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7476\,
            I => \N__7472\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7475\,
            I => \N__7465\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7472\,
            I => \N__7461\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7471\,
            I => \N__7458\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7470\,
            I => \N__7455\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__7469\,
            I => \N__7452\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7468\,
            I => \N__7447\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7465\,
            I => \N__7444\
        );

    \I__1482\ : CascadeMux
    port map (
            O => \N__7464\,
            I => \N__7440\
        );

    \I__1481\ : Span4Mux_h
    port map (
            O => \N__7461\,
            I => \N__7435\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__7458\,
            I => \N__7435\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7455\,
            I => \N__7432\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7452\,
            I => \N__7429\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7451\,
            I => \N__7424\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7450\,
            I => \N__7424\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__7447\,
            I => \N__7421\
        );

    \I__1474\ : Span4Mux_h
    port map (
            O => \N__7444\,
            I => \N__7418\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7443\,
            I => \N__7413\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7440\,
            I => \N__7413\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__7435\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1470\ : Odrv12
    port map (
            O => \N__7432\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7429\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7424\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1467\ : Odrv12
    port map (
            O => \N__7421\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1466\ : Odrv4
    port map (
            O => \N__7418\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7413\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7398\,
            I => \N__7395\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7395\,
            I => \N__7388\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7394\,
            I => \N__7383\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7393\,
            I => \N__7383\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7392\,
            I => \N__7378\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7391\,
            I => \N__7378\
        );

    \I__1458\ : Odrv4
    port map (
            O => \N__7388\,
            I => \U409_AUTOCONFIG.un1_STATE_1_0_a2_0\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7383\,
            I => \U409_AUTOCONFIG.un1_STATE_1_0_a2_0\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7378\,
            I => \U409_AUTOCONFIG.un1_STATE_1_0_a2_0\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7371\,
            I => \N__7357\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7370\,
            I => \N__7357\
        );

    \I__1453\ : InMux
    port map (
            O => \N__7369\,
            I => \N__7350\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7368\,
            I => \N__7350\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7367\,
            I => \N__7350\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__7366\,
            I => \N__7347\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__7365\,
            I => \N__7343\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__7364\,
            I => \N__7340\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__7363\,
            I => \N__7337\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__7362\,
            I => \N__7334\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7357\,
            I => \N__7320\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__7350\,
            I => \N__7320\
        );

    \I__1443\ : InMux
    port map (
            O => \N__7347\,
            I => \N__7317\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7346\,
            I => \N__7312\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7343\,
            I => \N__7312\
        );

    \I__1440\ : InMux
    port map (
            O => \N__7340\,
            I => \N__7305\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7337\,
            I => \N__7305\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7334\,
            I => \N__7305\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7294\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7294\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7331\,
            I => \N__7294\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7330\,
            I => \N__7294\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7329\,
            I => \N__7294\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7328\,
            I => \N__7291\
        );

    \I__1431\ : InMux
    port map (
            O => \N__7327\,
            I => \N__7286\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7326\,
            I => \N__7286\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__7325\,
            I => \N__7281\
        );

    \I__1428\ : Span4Mux_v
    port map (
            O => \N__7320\,
            I => \N__7275\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__7317\,
            I => \N__7275\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__7312\,
            I => \N__7272\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7305\,
            I => \N__7263\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__7294\,
            I => \N__7263\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__7291\,
            I => \N__7263\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7286\,
            I => \N__7263\
        );

    \I__1421\ : InMux
    port map (
            O => \N__7285\,
            I => \N__7258\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7284\,
            I => \N__7258\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7281\,
            I => \N__7255\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7280\,
            I => \N__7252\
        );

    \I__1417\ : Span4Mux_v
    port map (
            O => \N__7275\,
            I => \N__7249\
        );

    \I__1416\ : Span4Mux_v
    port map (
            O => \N__7272\,
            I => \N__7246\
        );

    \I__1415\ : Span4Mux_v
    port map (
            O => \N__7263\,
            I => \N__7243\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__7258\,
            I => \N__7236\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__7255\,
            I => \N__7236\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__7252\,
            I => \N__7236\
        );

    \I__1411\ : Sp12to4
    port map (
            O => \N__7249\,
            I => \N__7229\
        );

    \I__1410\ : Sp12to4
    port map (
            O => \N__7246\,
            I => \N__7229\
        );

    \I__1409\ : Sp12to4
    port map (
            O => \N__7243\,
            I => \N__7229\
        );

    \I__1408\ : Span12Mux_h
    port map (
            O => \N__7236\,
            I => \N__7226\
        );

    \I__1407\ : Span12Mux_h
    port map (
            O => \N__7229\,
            I => \N__7223\
        );

    \I__1406\ : Span12Mux_v
    port map (
            O => \N__7226\,
            I => \N__7220\
        );

    \I__1405\ : Span12Mux_v
    port map (
            O => \N__7223\,
            I => \N__7217\
        );

    \I__1404\ : Odrv12
    port map (
            O => \N__7220\,
            I => \A_c_1\
        );

    \I__1403\ : Odrv12
    port map (
            O => \N__7217\,
            I => \A_c_1\
        );

    \I__1402\ : IoInMux
    port map (
            O => \N__7212\,
            I => \N__7209\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7209\,
            I => \N__7206\
        );

    \I__1400\ : Span4Mux_s3_v
    port map (
            O => \N__7206\,
            I => \N__7203\
        );

    \I__1399\ : Sp12to4
    port map (
            O => \N__7203\,
            I => \N__7198\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7202\,
            I => \N__7195\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7201\,
            I => \N__7192\
        );

    \I__1396\ : Span12Mux_h
    port map (
            O => \N__7198\,
            I => \N__7189\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7195\,
            I => \N__7183\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__7192\,
            I => \N__7183\
        );

    \I__1393\ : Span12Mux_v
    port map (
            O => \N__7189\,
            I => \N__7179\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7188\,
            I => \N__7176\
        );

    \I__1391\ : Span4Mux_h
    port map (
            O => \N__7183\,
            I => \N__7173\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7182\,
            I => \N__7170\
        );

    \I__1389\ : Odrv12
    port map (
            O => \N__7179\,
            I => \CONFIGENn_c\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__7176\,
            I => \CONFIGENn_c\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__7173\,
            I => \CONFIGENn_c\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7170\,
            I => \CONFIGENn_c\
        );

    \I__1385\ : InMux
    port map (
            O => \N__7161\,
            I => \N__7157\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7160\,
            I => \N__7154\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__7157\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__7154\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7149\,
            I => \N__7146\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7146\,
            I => \N__7143\
        );

    \I__1379\ : Odrv4
    port map (
            O => \N__7143\,
            I => \AC_TACK\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7136\
        );

    \I__1377\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7131\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__7136\,
            I => \N__7128\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7125\
        );

    \I__1374\ : CascadeMux
    port map (
            O => \N__7134\,
            I => \N__7122\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__7131\,
            I => \N__7118\
        );

    \I__1372\ : Span4Mux_v
    port map (
            O => \N__7128\,
            I => \N__7113\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7125\,
            I => \N__7113\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7122\,
            I => \N__7110\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7121\,
            I => \N__7107\
        );

    \I__1368\ : Span4Mux_v
    port map (
            O => \N__7118\,
            I => \N__7104\
        );

    \I__1367\ : Span4Mux_h
    port map (
            O => \N__7113\,
            I => \N__7101\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__7110\,
            I => \N__7094\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__7107\,
            I => \N__7094\
        );

    \I__1364\ : Sp12to4
    port map (
            O => \N__7104\,
            I => \N__7094\
        );

    \I__1363\ : Span4Mux_h
    port map (
            O => \N__7101\,
            I => \N__7091\
        );

    \I__1362\ : Span12Mux_h
    port map (
            O => \N__7094\,
            I => \N__7088\
        );

    \I__1361\ : Sp12to4
    port map (
            O => \N__7091\,
            I => \N__7085\
        );

    \I__1360\ : Span12Mux_v
    port map (
            O => \N__7088\,
            I => \N__7082\
        );

    \I__1359\ : Span12Mux_v
    port map (
            O => \N__7085\,
            I => \N__7079\
        );

    \I__1358\ : Odrv12
    port map (
            O => \N__7082\,
            I => \RnW_c\
        );

    \I__1357\ : Odrv12
    port map (
            O => \N__7079\,
            I => \RnW_c\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__7074\,
            I => \N__7071\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7071\,
            I => \N__7068\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7068\,
            I => \N__7064\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7067\,
            I => \N__7061\
        );

    \I__1352\ : Span4Mux_v
    port map (
            O => \N__7064\,
            I => \N__7056\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7061\,
            I => \N__7053\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7060\,
            I => \N__7048\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7059\,
            I => \N__7048\
        );

    \I__1348\ : Odrv4
    port map (
            O => \N__7056\,
            I => \N_356\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__7053\,
            I => \N_356\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7048\,
            I => \N_356\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7032\
        );

    \I__1344\ : InMux
    port map (
            O => \N__7040\,
            I => \N__7027\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7039\,
            I => \N__7027\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7038\,
            I => \N__7024\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7037\,
            I => \N__7017\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7036\,
            I => \N__7017\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7035\,
            I => \N__7017\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__7032\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__7027\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7024\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7017\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1334\ : InMux
    port map (
            O => \N__7008\,
            I => \N__7002\
        );

    \I__1333\ : InMux
    port map (
            O => \N__7007\,
            I => \N__6999\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7006\,
            I => \N__6994\
        );

    \I__1331\ : InMux
    port map (
            O => \N__7005\,
            I => \N__6994\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__7002\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6999\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__6994\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1327\ : InMux
    port map (
            O => \N__6987\,
            I => \N__6980\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6986\,
            I => \N__6977\
        );

    \I__1325\ : InMux
    port map (
            O => \N__6985\,
            I => \N__6974\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6984\,
            I => \N__6971\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6983\,
            I => \N__6968\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6980\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6977\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6974\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6971\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__6968\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__6957\,
            I => \N__6953\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6956\,
            I => \N__6949\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6953\,
            I => \N__6944\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6952\,
            I => \N__6944\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6949\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6944\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__1311\ : CascadeMux
    port map (
            O => \N__6939\,
            I => \N__6936\
        );

    \I__1310\ : InMux
    port map (
            O => \N__6936\,
            I => \N__6933\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6933\,
            I => \N__6928\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6925\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__6931\,
            I => \N__6922\
        );

    \I__1306\ : Span4Mux_h
    port map (
            O => \N__6928\,
            I => \N__6915\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6925\,
            I => \N__6915\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6922\,
            I => \N__6912\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6921\,
            I => \N__6906\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6920\,
            I => \N__6906\
        );

    \I__1301\ : Span4Mux_v
    port map (
            O => \N__6915\,
            I => \N__6901\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6912\,
            I => \N__6901\
        );

    \I__1299\ : CascadeMux
    port map (
            O => \N__6911\,
            I => \N__6897\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6906\,
            I => \N__6894\
        );

    \I__1297\ : Span4Mux_v
    port map (
            O => \N__6901\,
            I => \N__6890\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6887\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6897\,
            I => \N__6884\
        );

    \I__1294\ : Span4Mux_v
    port map (
            O => \N__6894\,
            I => \N__6881\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6878\
        );

    \I__1292\ : Sp12to4
    port map (
            O => \N__6890\,
            I => \N__6867\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__6887\,
            I => \N__6867\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__6884\,
            I => \N__6867\
        );

    \I__1289\ : Sp12to4
    port map (
            O => \N__6881\,
            I => \N__6867\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6878\,
            I => \N__6867\
        );

    \I__1287\ : Span12Mux_h
    port map (
            O => \N__6867\,
            I => \N__6864\
        );

    \I__1286\ : Odrv12
    port map (
            O => \N__6864\,
            I => \A_c_20\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__6861\,
            I => \U409_TRANSFER_ACK.N_346_cascade_\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6858\,
            I => \N__6855\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6855\,
            I => \N__6851\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6854\,
            I => \N__6848\
        );

    \I__1281\ : Span4Mux_v
    port map (
            O => \N__6851\,
            I => \N__6843\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__6848\,
            I => \N__6843\
        );

    \I__1279\ : Span4Mux_h
    port map (
            O => \N__6843\,
            I => \N__6839\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6836\
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__6839\,
            I => \N_434\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__6836\,
            I => \N_434\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__6831\,
            I => \N_190_cascade_\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6828\,
            I => \N__6825\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__6825\,
            I => \N__6822\
        );

    \I__1272\ : Span12Mux_h
    port map (
            O => \N__6822\,
            I => \N__6819\
        );

    \I__1271\ : Span12Mux_h
    port map (
            O => \N__6819\,
            I => \N__6816\
        );

    \I__1270\ : Span12Mux_v
    port map (
            O => \N__6816\,
            I => \N__6813\
        );

    \I__1269\ : Odrv12
    port map (
            O => \N__6813\,
            I => \TACKn_in\
        );

    \I__1268\ : SRMux
    port map (
            O => \N__6810\,
            I => \N__6805\
        );

    \I__1267\ : SRMux
    port map (
            O => \N__6809\,
            I => \N__6802\
        );

    \I__1266\ : SRMux
    port map (
            O => \N__6808\,
            I => \N__6799\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6805\,
            I => \N__6792\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6802\,
            I => \N__6792\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__6799\,
            I => \N__6792\
        );

    \I__1262\ : Span4Mux_v
    port map (
            O => \N__6792\,
            I => \N__6789\
        );

    \I__1261\ : Span4Mux_v
    port map (
            O => \N__6789\,
            I => \N__6786\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__6786\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1259\ : InMux
    port map (
            O => \N__6783\,
            I => \N__6779\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6776\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6779\,
            I => \N__6771\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__6776\,
            I => \N__6768\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6765\
        );

    \I__1254\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6760\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__6771\,
            I => \N__6753\
        );

    \I__1252\ : Span4Mux_h
    port map (
            O => \N__6768\,
            I => \N__6753\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__6765\,
            I => \N__6753\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6764\,
            I => \N__6750\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6763\,
            I => \N__6747\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6760\,
            I => \N__6738\
        );

    \I__1247\ : Span4Mux_h
    port map (
            O => \N__6753\,
            I => \N__6738\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6750\,
            I => \N__6738\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6747\,
            I => \N__6738\
        );

    \I__1244\ : Span4Mux_v
    port map (
            O => \N__6738\,
            I => \N__6732\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6727\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6727\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6735\,
            I => \N__6724\
        );

    \I__1240\ : Sp12to4
    port map (
            O => \N__6732\,
            I => \N__6717\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__6727\,
            I => \N__6717\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6724\,
            I => \N__6714\
        );

    \I__1237\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6709\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6722\,
            I => \N__6709\
        );

    \I__1235\ : Span12Mux_h
    port map (
            O => \N__6717\,
            I => \N__6702\
        );

    \I__1234\ : Sp12to4
    port map (
            O => \N__6714\,
            I => \N__6702\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6709\,
            I => \N__6702\
        );

    \I__1232\ : Odrv12
    port map (
            O => \N__6702\,
            I => \A_c_21\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6699\,
            I => \N__6689\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6698\,
            I => \N__6689\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6697\,
            I => \N__6686\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6696\,
            I => \N__6683\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6695\,
            I => \N__6680\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__6694\,
            I => \N__6677\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6689\,
            I => \N__6674\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6686\,
            I => \N__6671\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6683\,
            I => \N__6666\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__6680\,
            I => \N__6666\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6677\,
            I => \N__6663\
        );

    \I__1220\ : Span4Mux_v
    port map (
            O => \N__6674\,
            I => \N__6654\
        );

    \I__1219\ : Span4Mux_v
    port map (
            O => \N__6671\,
            I => \N__6654\
        );

    \I__1218\ : Span4Mux_v
    port map (
            O => \N__6666\,
            I => \N__6654\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__6663\,
            I => \N__6651\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6662\,
            I => \N__6646\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6646\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__6654\,
            I => \N_351\
        );

    \I__1213\ : Odrv12
    port map (
            O => \N__6651\,
            I => \N_351\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6646\,
            I => \N_351\
        );

    \I__1211\ : IoInMux
    port map (
            O => \N__6639\,
            I => \N__6636\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6636\,
            I => \N__6633\
        );

    \I__1209\ : IoSpan4Mux
    port map (
            O => \N__6633\,
            I => \N__6630\
        );

    \I__1208\ : Sp12to4
    port map (
            O => \N__6630\,
            I => \N__6627\
        );

    \I__1207\ : Span12Mux_s7_h
    port map (
            O => \N__6627\,
            I => \N__6624\
        );

    \I__1206\ : Span12Mux_h
    port map (
            O => \N__6624\,
            I => \N__6621\
        );

    \I__1205\ : Span12Mux_v
    port map (
            O => \N__6621\,
            I => \N__6618\
        );

    \I__1204\ : Odrv12
    port map (
            O => \N__6618\,
            I => \N_436_i\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6615\,
            I => \N__6609\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6603\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6600\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6612\,
            I => \N__6597\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6609\,
            I => \N__6594\
        );

    \I__1198\ : CascadeMux
    port map (
            O => \N__6608\,
            I => \N__6591\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__6607\,
            I => \N__6587\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__6606\,
            I => \N__6583\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__6603\,
            I => \N__6578\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__6600\,
            I => \N__6578\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6597\,
            I => \N__6573\
        );

    \I__1192\ : Span4Mux_v
    port map (
            O => \N__6594\,
            I => \N__6573\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6591\,
            I => \N__6570\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6590\,
            I => \N__6567\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6587\,
            I => \N__6564\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6561\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6558\
        );

    \I__1186\ : Span4Mux_v
    port map (
            O => \N__6578\,
            I => \N__6551\
        );

    \I__1185\ : Span4Mux_h
    port map (
            O => \N__6573\,
            I => \N__6551\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6570\,
            I => \N__6551\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6567\,
            I => \N__6548\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6564\,
            I => \N__6541\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6561\,
            I => \N__6541\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6558\,
            I => \N__6541\
        );

    \I__1179\ : Sp12to4
    port map (
            O => \N__6551\,
            I => \N__6538\
        );

    \I__1178\ : Span4Mux_v
    port map (
            O => \N__6548\,
            I => \N__6533\
        );

    \I__1177\ : Span4Mux_v
    port map (
            O => \N__6541\,
            I => \N__6533\
        );

    \I__1176\ : Span12Mux_v
    port map (
            O => \N__6538\,
            I => \N__6528\
        );

    \I__1175\ : Sp12to4
    port map (
            O => \N__6533\,
            I => \N__6528\
        );

    \I__1174\ : Span12Mux_h
    port map (
            O => \N__6528\,
            I => \N__6525\
        );

    \I__1173\ : Span12Mux_v
    port map (
            O => \N__6525\,
            I => \N__6522\
        );

    \I__1172\ : Odrv12
    port map (
            O => \N__6522\,
            I => \A_c_17\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6516\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6516\,
            I => \N__6512\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6515\,
            I => \N__6509\
        );

    \I__1168\ : Odrv4
    port map (
            O => \N__6512\,
            I => \N_431\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__6509\,
            I => \N_431\
        );

    \I__1166\ : CascadeMux
    port map (
            O => \N__6504\,
            I => \N__6501\
        );

    \I__1165\ : InMux
    port map (
            O => \N__6501\,
            I => \N__6498\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__6498\,
            I => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_7\
        );

    \I__1163\ : CascadeMux
    port map (
            O => \N__6495\,
            I => \N__6491\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6494\,
            I => \N__6488\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6485\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__6488\,
            I => \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_o2dupZ0\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6485\,
            I => \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_o2dupZ0\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__6480\,
            I => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_0Z0Z_3_cascade_\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6477\,
            I => \N__6471\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6476\,
            I => \N__6471\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6471\,
            I => \U409_ADDRESS_DECODE.ATA_ENZ0\
        );

    \I__1154\ : IoInMux
    port map (
            O => \N__6468\,
            I => \N__6465\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6465\,
            I => \N__6462\
        );

    \I__1152\ : Span12Mux_s10_h
    port map (
            O => \N__6462\,
            I => \N__6459\
        );

    \I__1151\ : Odrv12
    port map (
            O => \N__6459\,
            I => \N_107\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6456\,
            I => \N__6452\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6455\,
            I => \N__6449\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6452\,
            I => \N__6443\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6449\,
            I => \N__6443\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6448\,
            I => \N__6440\
        );

    \I__1145\ : Span4Mux_v
    port map (
            O => \N__6443\,
            I => \N__6437\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6440\,
            I => \N__6434\
        );

    \I__1143\ : Span4Mux_v
    port map (
            O => \N__6437\,
            I => \N__6431\
        );

    \I__1142\ : Span4Mux_v
    port map (
            O => \N__6434\,
            I => \N__6428\
        );

    \I__1141\ : Span4Mux_v
    port map (
            O => \N__6431\,
            I => \N__6425\
        );

    \I__1140\ : Sp12to4
    port map (
            O => \N__6428\,
            I => \N__6422\
        );

    \I__1139\ : Sp12to4
    port map (
            O => \N__6425\,
            I => \N__6417\
        );

    \I__1138\ : Span12Mux_v
    port map (
            O => \N__6422\,
            I => \N__6417\
        );

    \I__1137\ : Odrv12
    port map (
            O => \N__6417\,
            I => \A_c_16\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6414\,
            I => \N__6411\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6411\,
            I => \N__6407\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__6410\,
            I => \N__6404\
        );

    \I__1133\ : Span4Mux_v
    port map (
            O => \N__6407\,
            I => \N__6401\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6404\,
            I => \N__6398\
        );

    \I__1131\ : Odrv4
    port map (
            O => \N__6401\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__6398\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6393\,
            I => \N__6390\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6390\,
            I => \N__6386\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6389\,
            I => \N__6383\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__6386\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6383\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__6378\,
            I => \N__6373\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6377\,
            I => \N__6370\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6376\,
            I => \N__6367\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6373\,
            I => \N__6364\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__6370\,
            I => \N__6359\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6367\,
            I => \N__6354\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6364\,
            I => \N__6354\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6363\,
            I => \N__6351\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6362\,
            I => \N__6348\
        );

    \I__1115\ : Odrv4
    port map (
            O => \N__6359\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1114\ : Odrv4
    port map (
            O => \N__6354\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__6351\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6348\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1111\ : IoInMux
    port map (
            O => \N__6339\,
            I => \N__6336\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6336\,
            I => \N__6333\
        );

    \I__1109\ : IoSpan4Mux
    port map (
            O => \N__6333\,
            I => \N__6330\
        );

    \I__1108\ : Sp12to4
    port map (
            O => \N__6330\,
            I => \N__6327\
        );

    \I__1107\ : Span12Mux_s9_v
    port map (
            O => \N__6327\,
            I => \N__6324\
        );

    \I__1106\ : Odrv12
    port map (
            O => \N__6324\,
            I => \N_128\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6321\,
            I => \N__6313\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6320\,
            I => \N__6313\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6319\,
            I => \N__6310\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6318\,
            I => \N__6307\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__6313\,
            I => \N__6303\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6310\,
            I => \N__6300\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6307\,
            I => \N__6297\
        );

    \I__1098\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6294\
        );

    \I__1097\ : Span4Mux_v
    port map (
            O => \N__6303\,
            I => \N__6291\
        );

    \I__1096\ : Span4Mux_h
    port map (
            O => \N__6300\,
            I => \N__6284\
        );

    \I__1095\ : Span4Mux_v
    port map (
            O => \N__6297\,
            I => \N__6284\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6294\,
            I => \N__6284\
        );

    \I__1093\ : Span4Mux_v
    port map (
            O => \N__6291\,
            I => \N__6281\
        );

    \I__1092\ : Span4Mux_v
    port map (
            O => \N__6284\,
            I => \N__6278\
        );

    \I__1091\ : Sp12to4
    port map (
            O => \N__6281\,
            I => \N__6275\
        );

    \I__1090\ : Span4Mux_h
    port map (
            O => \N__6278\,
            I => \N__6272\
        );

    \I__1089\ : Span12Mux_h
    port map (
            O => \N__6275\,
            I => \N__6267\
        );

    \I__1088\ : Sp12to4
    port map (
            O => \N__6272\,
            I => \N__6267\
        );

    \I__1087\ : Odrv12
    port map (
            O => \N__6267\,
            I => \TSn_c\
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__6264\,
            I => \N__6257\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6263\,
            I => \N__6253\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6262\,
            I => \N__6248\
        );

    \I__1083\ : InMux
    port map (
            O => \N__6261\,
            I => \N__6248\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6241\
        );

    \I__1081\ : InMux
    port map (
            O => \N__6257\,
            I => \N__6241\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6256\,
            I => \N__6241\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6253\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6248\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__6241\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6234\,
            I => \N__6230\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6233\,
            I => \N__6227\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__6230\,
            I => \U409_TRANSFER_ACK.N_268\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__6227\,
            I => \U409_TRANSFER_ACK.N_268\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6222\,
            I => \N__6218\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6221\,
            I => \N__6215\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__6218\,
            I => \U409_TRANSFER_ACK.N_237\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6215\,
            I => \U409_TRANSFER_ACK.N_237\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__6210\,
            I => \N__6206\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__6209\,
            I => \N__6203\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6206\,
            I => \N__6200\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6197\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__6200\,
            I => \N__6192\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__6197\,
            I => \N__6192\
        );

    \I__1062\ : Span4Mux_v
    port map (
            O => \N__6192\,
            I => \N__6188\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__6191\,
            I => \N__6185\
        );

    \I__1060\ : Span4Mux_v
    port map (
            O => \N__6188\,
            I => \N__6182\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6179\
        );

    \I__1058\ : Sp12to4
    port map (
            O => \N__6182\,
            I => \N__6176\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6179\,
            I => \N__6173\
        );

    \I__1056\ : Span12Mux_h
    port map (
            O => \N__6176\,
            I => \N__6168\
        );

    \I__1055\ : Span12Mux_v
    port map (
            O => \N__6173\,
            I => \N__6168\
        );

    \I__1054\ : Odrv12
    port map (
            O => \N__6168\,
            I => \D_in_6\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6165\,
            I => \N__6161\
        );

    \I__1052\ : InMux
    port map (
            O => \N__6164\,
            I => \N__6158\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6161\,
            I => \ATA_BASE_6\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6158\,
            I => \ATA_BASE_6\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__6153\,
            I => \N__6150\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6150\,
            I => \N__6146\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6149\,
            I => \N__6143\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6146\,
            I => \ATA_BASE_1\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__6143\,
            I => \ATA_BASE_1\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6138\,
            I => \N__6134\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6137\,
            I => \N__6131\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6134\,
            I => \ATA_BASE_0\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__6131\,
            I => \ATA_BASE_0\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__6126\,
            I => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7Z0Z_0_cascade_\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__6123\,
            I => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_7_cascade_\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__6120\,
            I => \U409_ADDRESS_DECODE.ATA_EN_2_0_o2_3_cascade_\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6117\,
            I => \N__6113\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6116\,
            I => \N__6108\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6113\,
            I => \N__6105\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6112\,
            I => \N__6102\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6111\,
            I => \N__6099\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6108\,
            I => \N__6092\
        );

    \I__1031\ : Span4Mux_h
    port map (
            O => \N__6105\,
            I => \N__6092\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6102\,
            I => \N__6092\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6099\,
            I => \N__6089\
        );

    \I__1028\ : Span4Mux_v
    port map (
            O => \N__6092\,
            I => \N__6085\
        );

    \I__1027\ : Span4Mux_v
    port map (
            O => \N__6089\,
            I => \N__6082\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6079\
        );

    \I__1025\ : Sp12to4
    port map (
            O => \N__6085\,
            I => \N__6072\
        );

    \I__1024\ : Sp12to4
    port map (
            O => \N__6082\,
            I => \N__6072\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__6079\,
            I => \N__6072\
        );

    \I__1022\ : Span12Mux_h
    port map (
            O => \N__6072\,
            I => \N__6069\
        );

    \I__1021\ : Span12Mux_v
    port map (
            O => \N__6069\,
            I => \N__6066\
        );

    \I__1020\ : Odrv12
    port map (
            O => \N__6066\,
            I => \A_c_18\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6063\,
            I => \N__6059\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6062\,
            I => \N__6056\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__6059\,
            I => \ATA_BASE_2\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__6056\,
            I => \ATA_BASE_2\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6048\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__6048\,
            I => \U409_ADDRESS_DECODE.N_183_i\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6045\,
            I => \N__6042\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6042\,
            I => \U409_ADDRESS_DECODE.ATA_EN_2_0_o2_2\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6039\,
            I => \N__6033\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6033\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6033\,
            I => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_2\
        );

    \I__1008\ : InMux
    port map (
            O => \N__6030\,
            I => \N__6024\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6029\,
            I => \N__6024\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6024\,
            I => \N__6021\
        );

    \I__1005\ : Span4Mux_v
    port map (
            O => \N__6021\,
            I => \N__6018\
        );

    \I__1004\ : Span4Mux_v
    port map (
            O => \N__6018\,
            I => \N__6015\
        );

    \I__1003\ : Odrv4
    port map (
            O => \N__6015\,
            I => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_0\
        );

    \I__1002\ : CascadeMux
    port map (
            O => \N__6012\,
            I => \N__6008\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6011\,
            I => \N__6003\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6008\,
            I => \N__5996\
        );

    \I__999\ : InMux
    port map (
            O => \N__6007\,
            I => \N__5996\
        );

    \I__998\ : InMux
    port map (
            O => \N__6006\,
            I => \N__5993\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__6003\,
            I => \N__5990\
        );

    \I__996\ : InMux
    port map (
            O => \N__6002\,
            I => \N__5985\
        );

    \I__995\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5985\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5996\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5993\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__992\ : Odrv12
    port map (
            O => \N__5990\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5985\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__990\ : InMux
    port map (
            O => \N__5976\,
            I => \N__5971\
        );

    \I__989\ : InMux
    port map (
            O => \N__5975\,
            I => \N__5966\
        );

    \I__988\ : InMux
    port map (
            O => \N__5974\,
            I => \N__5963\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__5971\,
            I => \N__5960\
        );

    \I__986\ : InMux
    port map (
            O => \N__5970\,
            I => \N__5955\
        );

    \I__985\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5955\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5966\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5963\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__982\ : Odrv4
    port map (
            O => \N__5960\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5955\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__980\ : InMux
    port map (
            O => \N__5946\,
            I => \N__5943\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__5943\,
            I => \N__5939\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__5942\,
            I => \N__5936\
        );

    \I__977\ : Span4Mux_v
    port map (
            O => \N__5939\,
            I => \N__5933\
        );

    \I__976\ : InMux
    port map (
            O => \N__5936\,
            I => \N__5930\
        );

    \I__975\ : Odrv4
    port map (
            O => \N__5933\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__5930\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\
        );

    \I__973\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5922\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5922\,
            I => \N__5919\
        );

    \I__971\ : Span4Mux_v
    port map (
            O => \N__5919\,
            I => \N__5915\
        );

    \I__970\ : InMux
    port map (
            O => \N__5918\,
            I => \N__5912\
        );

    \I__969\ : Odrv4
    port map (
            O => \N__5915\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5912\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\
        );

    \I__967\ : IoInMux
    port map (
            O => \N__5907\,
            I => \N__5904\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5904\,
            I => \N__5901\
        );

    \I__965\ : IoSpan4Mux
    port map (
            O => \N__5901\,
            I => \N__5898\
        );

    \I__964\ : Span4Mux_s2_v
    port map (
            O => \N__5898\,
            I => \N__5895\
        );

    \I__963\ : Sp12to4
    port map (
            O => \N__5895\,
            I => \N__5892\
        );

    \I__962\ : Odrv12
    port map (
            O => \N__5892\,
            I => \N_130\
        );

    \I__961\ : InMux
    port map (
            O => \N__5889\,
            I => \N__5883\
        );

    \I__960\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5883\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__5883\,
            I => \ATA_BASE_4\
        );

    \I__958\ : InMux
    port map (
            O => \N__5880\,
            I => \N__5874\
        );

    \I__957\ : InMux
    port map (
            O => \N__5879\,
            I => \N__5874\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__5874\,
            I => \ATA_BASE_5\
        );

    \I__955\ : CascadeMux
    port map (
            O => \N__5871\,
            I => \N__5866\
        );

    \I__954\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5861\
        );

    \I__953\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5861\
        );

    \I__952\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5858\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__5861\,
            I => \N__5855\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5858\,
            I => \N__5852\
        );

    \I__949\ : Span4Mux_v
    port map (
            O => \N__5855\,
            I => \N__5849\
        );

    \I__948\ : Span4Mux_v
    port map (
            O => \N__5852\,
            I => \N__5846\
        );

    \I__947\ : Sp12to4
    port map (
            O => \N__5849\,
            I => \N__5841\
        );

    \I__946\ : Sp12to4
    port map (
            O => \N__5846\,
            I => \N__5841\
        );

    \I__945\ : Span12Mux_h
    port map (
            O => \N__5841\,
            I => \N__5838\
        );

    \I__944\ : Odrv12
    port map (
            O => \N__5838\,
            I => \D_in_4\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__5835\,
            I => \N__5832\
        );

    \I__942\ : InMux
    port map (
            O => \N__5832\,
            I => \N__5826\
        );

    \I__941\ : InMux
    port map (
            O => \N__5831\,
            I => \N__5826\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5826\,
            I => \N__5823\
        );

    \I__939\ : Span4Mux_v
    port map (
            O => \N__5823\,
            I => \N__5819\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__5822\,
            I => \N__5816\
        );

    \I__937\ : Span4Mux_v
    port map (
            O => \N__5819\,
            I => \N__5813\
        );

    \I__936\ : InMux
    port map (
            O => \N__5816\,
            I => \N__5810\
        );

    \I__935\ : Sp12to4
    port map (
            O => \N__5813\,
            I => \N__5807\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5810\,
            I => \N__5804\
        );

    \I__933\ : Span12Mux_h
    port map (
            O => \N__5807\,
            I => \N__5799\
        );

    \I__932\ : Span12Mux_v
    port map (
            O => \N__5804\,
            I => \N__5799\
        );

    \I__931\ : Odrv12
    port map (
            O => \N__5799\,
            I => \D_in_5\
        );

    \I__930\ : InMux
    port map (
            O => \N__5796\,
            I => \N__5793\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5793\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3\
        );

    \I__928\ : InMux
    port map (
            O => \N__5790\,
            I => \N__5782\
        );

    \I__927\ : InMux
    port map (
            O => \N__5789\,
            I => \N__5782\
        );

    \I__926\ : InMux
    port map (
            O => \N__5788\,
            I => \N__5777\
        );

    \I__925\ : InMux
    port map (
            O => \N__5787\,
            I => \N__5777\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5782\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5777\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__5772\,
            I => \N__5768\
        );

    \I__921\ : InMux
    port map (
            O => \N__5771\,
            I => \N__5764\
        );

    \I__920\ : InMux
    port map (
            O => \N__5768\,
            I => \N__5759\
        );

    \I__919\ : InMux
    port map (
            O => \N__5767\,
            I => \N__5759\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5764\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__5759\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__5754\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_a2_3_cascade_\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__5751\,
            I => \U409_TRANSFER_ACK.N_268_cascade_\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__5748\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__5745\,
            I => \N__5742\
        );

    \I__912\ : InMux
    port map (
            O => \N__5742\,
            I => \N__5736\
        );

    \I__911\ : InMux
    port map (
            O => \N__5741\,
            I => \N__5736\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__5736\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__909\ : CascadeMux
    port map (
            O => \N__5733\,
            I => \N__5729\
        );

    \I__908\ : InMux
    port map (
            O => \N__5732\,
            I => \N__5724\
        );

    \I__907\ : InMux
    port map (
            O => \N__5729\,
            I => \N__5724\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5724\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__905\ : InMux
    port map (
            O => \N__5721\,
            I => \N__5718\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5718\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__5715\,
            I => \N__5710\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__5714\,
            I => \N__5707\
        );

    \I__901\ : InMux
    port map (
            O => \N__5713\,
            I => \N__5703\
        );

    \I__900\ : InMux
    port map (
            O => \N__5710\,
            I => \N__5696\
        );

    \I__899\ : InMux
    port map (
            O => \N__5707\,
            I => \N__5696\
        );

    \I__898\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5696\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5703\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5696\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__895\ : InMux
    port map (
            O => \N__5691\,
            I => \N__5688\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__5688\,
            I => \N__5685\
        );

    \I__893\ : Span4Mux_h
    port map (
            O => \N__5685\,
            I => \N__5680\
        );

    \I__892\ : InMux
    port map (
            O => \N__5684\,
            I => \N__5677\
        );

    \I__891\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5674\
        );

    \I__890\ : Span4Mux_h
    port map (
            O => \N__5680\,
            I => \N__5669\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__5677\,
            I => \N__5669\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5674\,
            I => \N__5666\
        );

    \I__887\ : Span4Mux_h
    port map (
            O => \N__5669\,
            I => \N__5663\
        );

    \I__886\ : Span12Mux_v
    port map (
            O => \N__5666\,
            I => \N__5660\
        );

    \I__885\ : Span4Mux_v
    port map (
            O => \N__5663\,
            I => \N__5657\
        );

    \I__884\ : Odrv12
    port map (
            O => \N__5660\,
            I => \A_c_31\
        );

    \I__883\ : Odrv4
    port map (
            O => \N__5657\,
            I => \A_c_31\
        );

    \I__882\ : InMux
    port map (
            O => \N__5652\,
            I => \N__5648\
        );

    \I__881\ : InMux
    port map (
            O => \N__5651\,
            I => \N__5645\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5648\,
            I => \BRIDGE_BASE_3\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5645\,
            I => \BRIDGE_BASE_3\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__5640\,
            I => \N__5637\
        );

    \I__877\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5633\
        );

    \I__876\ : InMux
    port map (
            O => \N__5636\,
            I => \N__5630\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5633\,
            I => \BRIDGE_BASE_2\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5630\,
            I => \BRIDGE_BASE_2\
        );

    \I__873\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5621\
        );

    \I__872\ : InMux
    port map (
            O => \N__5624\,
            I => \N__5618\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5621\,
            I => \N__5615\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5618\,
            I => \N__5611\
        );

    \I__869\ : Span4Mux_h
    port map (
            O => \N__5615\,
            I => \N__5608\
        );

    \I__868\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5605\
        );

    \I__867\ : Span4Mux_h
    port map (
            O => \N__5611\,
            I => \N__5602\
        );

    \I__866\ : Span4Mux_h
    port map (
            O => \N__5608\,
            I => \N__5597\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5605\,
            I => \N__5597\
        );

    \I__864\ : Sp12to4
    port map (
            O => \N__5602\,
            I => \N__5594\
        );

    \I__863\ : Span4Mux_h
    port map (
            O => \N__5597\,
            I => \N__5591\
        );

    \I__862\ : Span12Mux_v
    port map (
            O => \N__5594\,
            I => \N__5588\
        );

    \I__861\ : Span4Mux_v
    port map (
            O => \N__5591\,
            I => \N__5585\
        );

    \I__860\ : Odrv12
    port map (
            O => \N__5588\,
            I => \A_c_30\
        );

    \I__859\ : Odrv4
    port map (
            O => \N__5585\,
            I => \A_c_30\
        );

    \I__858\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5577\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__5577\,
            I => \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0Z0Z_1\
        );

    \I__856\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5562\
        );

    \I__855\ : InMux
    port map (
            O => \N__5573\,
            I => \N__5562\
        );

    \I__854\ : InMux
    port map (
            O => \N__5572\,
            I => \N__5562\
        );

    \I__853\ : InMux
    port map (
            O => \N__5571\,
            I => \N__5562\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5562\,
            I => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\
        );

    \I__851\ : InMux
    port map (
            O => \N__5559\,
            I => \N__5553\
        );

    \I__850\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5548\
        );

    \I__849\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5548\
        );

    \I__848\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5545\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__5553\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5548\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5545\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__844\ : InMux
    port map (
            O => \N__5538\,
            I => \N__5529\
        );

    \I__843\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5529\
        );

    \I__842\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5529\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5529\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_o2_5\
        );

    \I__840\ : InMux
    port map (
            O => \N__5526\,
            I => \N__5522\
        );

    \I__839\ : CascadeMux
    port map (
            O => \N__5525\,
            I => \N__5519\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5522\,
            I => \N__5516\
        );

    \I__837\ : InMux
    port map (
            O => \N__5519\,
            I => \N__5513\
        );

    \I__836\ : Span4Mux_v
    port map (
            O => \N__5516\,
            I => \N__5508\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__5513\,
            I => \N__5508\
        );

    \I__834\ : Odrv4
    port map (
            O => \N__5508\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\
        );

    \I__833\ : InMux
    port map (
            O => \N__5505\,
            I => \N__5502\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5502\,
            I => \N__5499\
        );

    \I__831\ : Span4Mux_v
    port map (
            O => \N__5499\,
            I => \N__5495\
        );

    \I__830\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5492\
        );

    \I__829\ : Odrv4
    port map (
            O => \N__5495\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5492\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\
        );

    \I__827\ : IoInMux
    port map (
            O => \N__5487\,
            I => \N__5484\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5484\,
            I => \N__5481\
        );

    \I__825\ : Sp12to4
    port map (
            O => \N__5481\,
            I => \N__5478\
        );

    \I__824\ : Span12Mux_s10_v
    port map (
            O => \N__5478\,
            I => \N__5475\
        );

    \I__823\ : Odrv12
    port map (
            O => \N__5475\,
            I => \N_126\
        );

    \I__822\ : IoInMux
    port map (
            O => \N__5472\,
            I => \N__5469\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5469\,
            I => \N__5466\
        );

    \I__820\ : IoSpan4Mux
    port map (
            O => \N__5466\,
            I => \N__5463\
        );

    \I__819\ : Span4Mux_s1_h
    port map (
            O => \N__5463\,
            I => \N__5460\
        );

    \I__818\ : Sp12to4
    port map (
            O => \N__5460\,
            I => \N__5457\
        );

    \I__817\ : Span12Mux_h
    port map (
            O => \N__5457\,
            I => \N__5454\
        );

    \I__816\ : Odrv12
    port map (
            O => \N__5454\,
            I => \N_96\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__5451\,
            I => \N__5448\
        );

    \I__814\ : InMux
    port map (
            O => \N__5448\,
            I => \N__5443\
        );

    \I__813\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5440\
        );

    \I__812\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5437\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5443\,
            I => \N__5432\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__5440\,
            I => \N__5432\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__5437\,
            I => \N__5429\
        );

    \I__808\ : Span4Mux_v
    port map (
            O => \N__5432\,
            I => \N__5426\
        );

    \I__807\ : Span12Mux_h
    port map (
            O => \N__5429\,
            I => \N__5423\
        );

    \I__806\ : Span4Mux_v
    port map (
            O => \N__5426\,
            I => \N__5420\
        );

    \I__805\ : Span12Mux_v
    port map (
            O => \N__5423\,
            I => \N__5417\
        );

    \I__804\ : Sp12to4
    port map (
            O => \N__5420\,
            I => \N__5414\
        );

    \I__803\ : Odrv12
    port map (
            O => \N__5417\,
            I => \A_c_29\
        );

    \I__802\ : Odrv12
    port map (
            O => \N__5414\,
            I => \A_c_29\
        );

    \I__801\ : InMux
    port map (
            O => \N__5409\,
            I => \N__5405\
        );

    \I__800\ : InMux
    port map (
            O => \N__5408\,
            I => \N__5402\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__5405\,
            I => \BRIDGE_BASE_1\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5402\,
            I => \BRIDGE_BASE_1\
        );

    \I__797\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5392\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__5396\,
            I => \N__5389\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__5395\,
            I => \N__5386\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__5392\,
            I => \N__5383\
        );

    \I__793\ : InMux
    port map (
            O => \N__5389\,
            I => \N__5380\
        );

    \I__792\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5377\
        );

    \I__791\ : Span4Mux_v
    port map (
            O => \N__5383\,
            I => \N__5374\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5380\,
            I => \N__5371\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5377\,
            I => \N__5368\
        );

    \I__788\ : Span4Mux_v
    port map (
            O => \N__5374\,
            I => \N__5365\
        );

    \I__787\ : Span12Mux_v
    port map (
            O => \N__5371\,
            I => \N__5360\
        );

    \I__786\ : Sp12to4
    port map (
            O => \N__5368\,
            I => \N__5360\
        );

    \I__785\ : Span4Mux_v
    port map (
            O => \N__5365\,
            I => \N__5357\
        );

    \I__784\ : Span12Mux_v
    port map (
            O => \N__5360\,
            I => \N__5354\
        );

    \I__783\ : Span4Mux_h
    port map (
            O => \N__5357\,
            I => \N__5351\
        );

    \I__782\ : Odrv12
    port map (
            O => \N__5354\,
            I => \A_c_28\
        );

    \I__781\ : Odrv4
    port map (
            O => \N__5351\,
            I => \A_c_28\
        );

    \I__780\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5342\
        );

    \I__779\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5339\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5342\,
            I => \BRIDGE_BASE_0\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5339\,
            I => \BRIDGE_BASE_0\
        );

    \I__776\ : InMux
    port map (
            O => \N__5334\,
            I => \N__5331\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5331\,
            I => \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0Z0Z_0\
        );

    \I__774\ : IoInMux
    port map (
            O => \N__5328\,
            I => \N__5325\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__5325\,
            I => \N__5320\
        );

    \I__772\ : IoInMux
    port map (
            O => \N__5324\,
            I => \N__5317\
        );

    \I__771\ : IoInMux
    port map (
            O => \N__5323\,
            I => \N__5314\
        );

    \I__770\ : IoSpan4Mux
    port map (
            O => \N__5320\,
            I => \N__5307\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5317\,
            I => \N__5307\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5314\,
            I => \N__5307\
        );

    \I__767\ : IoSpan4Mux
    port map (
            O => \N__5307\,
            I => \N__5303\
        );

    \I__766\ : IoInMux
    port map (
            O => \N__5306\,
            I => \N__5300\
        );

    \I__765\ : Span4Mux_s2_v
    port map (
            O => \N__5303\,
            I => \N__5297\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5300\,
            I => \N__5294\
        );

    \I__763\ : Sp12to4
    port map (
            O => \N__5297\,
            I => \N__5289\
        );

    \I__762\ : Span12Mux_s4_v
    port map (
            O => \N__5294\,
            I => \N__5289\
        );

    \I__761\ : Odrv12
    port map (
            O => \N__5289\,
            I => \D_1_i\
        );

    \I__760\ : InMux
    port map (
            O => \N__5286\,
            I => \N__5283\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5283\,
            I => \N__5280\
        );

    \I__758\ : Span4Mux_v
    port map (
            O => \N__5280\,
            I => \N__5277\
        );

    \I__757\ : Sp12to4
    port map (
            O => \N__5277\,
            I => \N__5274\
        );

    \I__756\ : Span12Mux_h
    port map (
            O => \N__5274\,
            I => \N__5271\
        );

    \I__755\ : Span12Mux_h
    port map (
            O => \N__5271\,
            I => \N__5268\
        );

    \I__754\ : Span12Mux_v
    port map (
            O => \N__5268\,
            I => \N__5265\
        );

    \I__753\ : Odrv12
    port map (
            O => \N__5265\,
            I => \AUTOBOOT_c\
        );

    \I__752\ : InMux
    port map (
            O => \N__5262\,
            I => \N__5258\
        );

    \I__751\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5255\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__5258\,
            I => \U409_AUTOCONFIG.N_360\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__5255\,
            I => \U409_AUTOCONFIG.N_360\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__5250\,
            I => \N__5244\
        );

    \I__747\ : InMux
    port map (
            O => \N__5249\,
            I => \N__5241\
        );

    \I__746\ : InMux
    port map (
            O => \N__5248\,
            I => \N__5236\
        );

    \I__745\ : InMux
    port map (
            O => \N__5247\,
            I => \N__5236\
        );

    \I__744\ : InMux
    port map (
            O => \N__5244\,
            I => \N__5233\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__5241\,
            I => \N__5224\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__5236\,
            I => \N__5221\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__5233\,
            I => \N__5218\
        );

    \I__740\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5211\
        );

    \I__739\ : InMux
    port map (
            O => \N__5231\,
            I => \N__5211\
        );

    \I__738\ : InMux
    port map (
            O => \N__5230\,
            I => \N__5211\
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__5229\,
            I => \N__5208\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__5228\,
            I => \N__5205\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__5227\,
            I => \N__5201\
        );

    \I__734\ : Span4Mux_v
    port map (
            O => \N__5224\,
            I => \N__5196\
        );

    \I__733\ : Span4Mux_v
    port map (
            O => \N__5221\,
            I => \N__5196\
        );

    \I__732\ : Span4Mux_v
    port map (
            O => \N__5218\,
            I => \N__5191\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__5211\,
            I => \N__5191\
        );

    \I__730\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5182\
        );

    \I__729\ : InMux
    port map (
            O => \N__5205\,
            I => \N__5182\
        );

    \I__728\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5182\
        );

    \I__727\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5182\
        );

    \I__726\ : Sp12to4
    port map (
            O => \N__5196\,
            I => \N__5175\
        );

    \I__725\ : Sp12to4
    port map (
            O => \N__5191\,
            I => \N__5175\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5182\,
            I => \N__5175\
        );

    \I__723\ : Odrv12
    port map (
            O => \N__5175\,
            I => \A_c_5\
        );

    \I__722\ : InMux
    port map (
            O => \N__5172\,
            I => \N__5169\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__5169\,
            I => \N__5162\
        );

    \I__720\ : InMux
    port map (
            O => \N__5168\,
            I => \N__5155\
        );

    \I__719\ : InMux
    port map (
            O => \N__5167\,
            I => \N__5155\
        );

    \I__718\ : InMux
    port map (
            O => \N__5166\,
            I => \N__5155\
        );

    \I__717\ : InMux
    port map (
            O => \N__5165\,
            I => \N__5148\
        );

    \I__716\ : Span4Mux_h
    port map (
            O => \N__5162\,
            I => \N__5143\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5155\,
            I => \N__5143\
        );

    \I__714\ : InMux
    port map (
            O => \N__5154\,
            I => \N__5140\
        );

    \I__713\ : InMux
    port map (
            O => \N__5153\,
            I => \N__5137\
        );

    \I__712\ : InMux
    port map (
            O => \N__5152\,
            I => \N__5132\
        );

    \I__711\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5132\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5148\,
            I => \N__5125\
        );

    \I__709\ : Span4Mux_h
    port map (
            O => \N__5143\,
            I => \N__5125\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__5140\,
            I => \N__5125\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__5137\,
            I => \N__5120\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5132\,
            I => \N__5120\
        );

    \I__705\ : Sp12to4
    port map (
            O => \N__5125\,
            I => \N__5117\
        );

    \I__704\ : Span12Mux_h
    port map (
            O => \N__5120\,
            I => \N__5114\
        );

    \I__703\ : Span12Mux_v
    port map (
            O => \N__5117\,
            I => \N__5111\
        );

    \I__702\ : Span12Mux_v
    port map (
            O => \N__5114\,
            I => \N__5108\
        );

    \I__701\ : Odrv12
    port map (
            O => \N__5111\,
            I => \A_c_3\
        );

    \I__700\ : Odrv12
    port map (
            O => \N__5108\,
            I => \A_c_3\
        );

    \I__699\ : CascadeMux
    port map (
            O => \N__5103\,
            I => \N__5100\
        );

    \I__698\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5097\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5097\,
            I => \N__5094\
        );

    \I__696\ : Span4Mux_v
    port map (
            O => \N__5094\,
            I => \N__5091\
        );

    \I__695\ : Odrv4
    port map (
            O => \N__5091\,
            I => \U409_AUTOCONFIG.N_276\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__5088\,
            I => \U409_ADDRESS_DECODE.PORTSIZE_iZ0Z_1_cascade_\
        );

    \I__693\ : IoInMux
    port map (
            O => \N__5085\,
            I => \N__5082\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5082\,
            I => \N__5079\
        );

    \I__691\ : IoSpan4Mux
    port map (
            O => \N__5079\,
            I => \N__5076\
        );

    \I__690\ : Span4Mux_s2_v
    port map (
            O => \N__5076\,
            I => \N__5073\
        );

    \I__689\ : Sp12to4
    port map (
            O => \N__5073\,
            I => \N__5070\
        );

    \I__688\ : Odrv12
    port map (
            O => \N__5070\,
            I => \N_139\
        );

    \I__687\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5064\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5064\,
            I => \N__5061\
        );

    \I__685\ : Span4Mux_v
    port map (
            O => \N__5061\,
            I => \N__5058\
        );

    \I__684\ : Odrv4
    port map (
            O => \N__5058\,
            I => \U409_ADDRESS_DECODE.N_343\
        );

    \I__683\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5051\
        );

    \I__682\ : InMux
    port map (
            O => \N__5054\,
            I => \N__5048\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5051\,
            I => \N__5043\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5048\,
            I => \N__5043\
        );

    \I__679\ : Span4Mux_v
    port map (
            O => \N__5043\,
            I => \N__5039\
        );

    \I__678\ : InMux
    port map (
            O => \N__5042\,
            I => \N__5036\
        );

    \I__677\ : Span4Mux_h
    port map (
            O => \N__5039\,
            I => \N__5033\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__5036\,
            I => \N__5030\
        );

    \I__675\ : Sp12to4
    port map (
            O => \N__5033\,
            I => \N__5027\
        );

    \I__674\ : Span12Mux_h
    port map (
            O => \N__5030\,
            I => \N__5024\
        );

    \I__673\ : Odrv12
    port map (
            O => \N__5027\,
            I => \TM_c_1\
        );

    \I__672\ : Odrv12
    port map (
            O => \N__5024\,
            I => \TM_c_1\
        );

    \I__671\ : InMux
    port map (
            O => \N__5019\,
            I => \N__5015\
        );

    \I__670\ : InMux
    port map (
            O => \N__5018\,
            I => \N__5012\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5015\,
            I => \N__5006\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5012\,
            I => \N__5006\
        );

    \I__667\ : InMux
    port map (
            O => \N__5011\,
            I => \N__5003\
        );

    \I__666\ : Span4Mux_v
    port map (
            O => \N__5006\,
            I => \N__4998\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5003\,
            I => \N__4998\
        );

    \I__664\ : Span4Mux_h
    port map (
            O => \N__4998\,
            I => \N__4995\
        );

    \I__663\ : Sp12to4
    port map (
            O => \N__4995\,
            I => \N__4992\
        );

    \I__662\ : Odrv12
    port map (
            O => \N__4992\,
            I => \TM_c_0\
        );

    \I__661\ : IoInMux
    port map (
            O => \N__4989\,
            I => \N__4986\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4986\,
            I => \N__4983\
        );

    \I__659\ : Span12Mux_s11_v
    port map (
            O => \N__4983\,
            I => \N__4980\
        );

    \I__658\ : Span12Mux_h
    port map (
            O => \N__4980\,
            I => \N__4977\
        );

    \I__657\ : Odrv12
    port map (
            O => \N__4977\,
            I => \N_265_i\
        );

    \I__656\ : CascadeMux
    port map (
            O => \N__4974\,
            I => \N__4969\
        );

    \I__655\ : CascadeMux
    port map (
            O => \N__4973\,
            I => \N__4966\
        );

    \I__654\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4959\
        );

    \I__653\ : InMux
    port map (
            O => \N__4969\,
            I => \N__4959\
        );

    \I__652\ : InMux
    port map (
            O => \N__4966\,
            I => \N__4959\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__4959\,
            I => \N__4956\
        );

    \I__650\ : Odrv12
    port map (
            O => \N__4956\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_o2_4\
        );

    \I__649\ : InMux
    port map (
            O => \N__4953\,
            I => \N__4949\
        );

    \I__648\ : InMux
    port map (
            O => \N__4952\,
            I => \N__4946\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__4949\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_0\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__4946\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_0\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__4941\,
            I => \N__4938\
        );

    \I__644\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4935\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4935\,
            I => \N__4931\
        );

    \I__642\ : InMux
    port map (
            O => \N__4934\,
            I => \N__4928\
        );

    \I__641\ : Odrv4
    port map (
            O => \N__4931\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ1Z_0\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4928\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ1Z_0\
        );

    \I__639\ : IoInMux
    port map (
            O => \N__4923\,
            I => \N__4920\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__4920\,
            I => \N__4917\
        );

    \I__637\ : Span12Mux_s2_v
    port map (
            O => \N__4917\,
            I => \N__4914\
        );

    \I__636\ : Odrv12
    port map (
            O => \N__4914\,
            I => \N_124\
        );

    \I__635\ : CascadeMux
    port map (
            O => \N__4911\,
            I => \N__4908\
        );

    \I__634\ : InMux
    port map (
            O => \N__4908\,
            I => \N__4905\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4905\,
            I => \U409_AUTOCONFIG.un1_STATE_1_0_a2_0Z0Z_2\
        );

    \I__632\ : CascadeMux
    port map (
            O => \N__4902\,
            I => \N__4899\
        );

    \I__631\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4896\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4896\,
            I => \N__4892\
        );

    \I__629\ : InMux
    port map (
            O => \N__4895\,
            I => \N__4889\
        );

    \I__628\ : Sp12to4
    port map (
            O => \N__4892\,
            I => \N__4884\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__4889\,
            I => \N__4884\
        );

    \I__626\ : Span12Mux_v
    port map (
            O => \N__4884\,
            I => \N__4881\
        );

    \I__625\ : Odrv12
    port map (
            O => \N__4881\,
            I => \CPUCONFn_c\
        );

    \I__624\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4874\
        );

    \I__623\ : InMux
    port map (
            O => \N__4877\,
            I => \N__4871\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__4874\,
            I => \U409_AUTOCONFIG.AC_STARTZ0\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__4871\,
            I => \U409_AUTOCONFIG.AC_STARTZ0\
        );

    \I__620\ : CascadeMux
    port map (
            O => \N__4866\,
            I => \N_354_cascade_\
        );

    \I__619\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4860\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__4860\,
            I => \N__4857\
        );

    \I__617\ : Odrv4
    port map (
            O => \N__4857\,
            I => \U409_AUTOCONFIG.N_273\
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__4854\,
            I => \N__4850\
        );

    \I__615\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4845\
        );

    \I__614\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4845\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__4845\,
            I => \U409_AUTOCONFIG.N_400\
        );

    \I__612\ : CascadeMux
    port map (
            O => \N__4842\,
            I => \N__4837\
        );

    \I__611\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4831\
        );

    \I__610\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4827\
        );

    \I__609\ : InMux
    port map (
            O => \N__4837\,
            I => \N__4818\
        );

    \I__608\ : InMux
    port map (
            O => \N__4836\,
            I => \N__4818\
        );

    \I__607\ : InMux
    port map (
            O => \N__4835\,
            I => \N__4818\
        );

    \I__606\ : InMux
    port map (
            O => \N__4834\,
            I => \N__4818\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4831\,
            I => \N__4813\
        );

    \I__604\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4806\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__4827\,
            I => \N__4801\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4818\,
            I => \N__4801\
        );

    \I__601\ : InMux
    port map (
            O => \N__4817\,
            I => \N__4796\
        );

    \I__600\ : InMux
    port map (
            O => \N__4816\,
            I => \N__4796\
        );

    \I__599\ : Span4Mux_v
    port map (
            O => \N__4813\,
            I => \N__4793\
        );

    \I__598\ : InMux
    port map (
            O => \N__4812\,
            I => \N__4786\
        );

    \I__597\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4786\
        );

    \I__596\ : InMux
    port map (
            O => \N__4810\,
            I => \N__4786\
        );

    \I__595\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4783\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__4806\,
            I => \N__4780\
        );

    \I__593\ : Span4Mux_v
    port map (
            O => \N__4801\,
            I => \N__4775\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4796\,
            I => \N__4775\
        );

    \I__591\ : Sp12to4
    port map (
            O => \N__4793\,
            I => \N__4768\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__4786\,
            I => \N__4768\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4783\,
            I => \N__4768\
        );

    \I__588\ : Span4Mux_v
    port map (
            O => \N__4780\,
            I => \N__4765\
        );

    \I__587\ : Span4Mux_v
    port map (
            O => \N__4775\,
            I => \N__4762\
        );

    \I__586\ : Span12Mux_h
    port map (
            O => \N__4768\,
            I => \N__4759\
        );

    \I__585\ : Sp12to4
    port map (
            O => \N__4765\,
            I => \N__4754\
        );

    \I__584\ : Sp12to4
    port map (
            O => \N__4762\,
            I => \N__4754\
        );

    \I__583\ : Span12Mux_v
    port map (
            O => \N__4759\,
            I => \N__4751\
        );

    \I__582\ : Span12Mux_h
    port map (
            O => \N__4754\,
            I => \N__4748\
        );

    \I__581\ : Odrv12
    port map (
            O => \N__4751\,
            I => \A_c_2\
        );

    \I__580\ : Odrv12
    port map (
            O => \N__4748\,
            I => \A_c_2\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__4743\,
            I => \N__4733\
        );

    \I__578\ : CascadeMux
    port map (
            O => \N__4742\,
            I => \N__4729\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__4741\,
            I => \N__4726\
        );

    \I__576\ : CascadeMux
    port map (
            O => \N__4740\,
            I => \N__4722\
        );

    \I__575\ : InMux
    port map (
            O => \N__4739\,
            I => \N__4718\
        );

    \I__574\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4711\
        );

    \I__573\ : InMux
    port map (
            O => \N__4737\,
            I => \N__4711\
        );

    \I__572\ : InMux
    port map (
            O => \N__4736\,
            I => \N__4711\
        );

    \I__571\ : InMux
    port map (
            O => \N__4733\,
            I => \N__4704\
        );

    \I__570\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4704\
        );

    \I__569\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4704\
        );

    \I__568\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4699\
        );

    \I__567\ : InMux
    port map (
            O => \N__4725\,
            I => \N__4699\
        );

    \I__566\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4696\
        );

    \I__565\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4693\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4718\,
            I => \N__4687\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4711\,
            I => \N__4687\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4704\,
            I => \N__4684\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__4699\,
            I => \N__4677\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4696\,
            I => \N__4677\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4693\,
            I => \N__4677\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__4692\,
            I => \N__4673\
        );

    \I__557\ : Span4Mux_v
    port map (
            O => \N__4687\,
            I => \N__4669\
        );

    \I__556\ : Span4Mux_v
    port map (
            O => \N__4684\,
            I => \N__4664\
        );

    \I__555\ : Span4Mux_v
    port map (
            O => \N__4677\,
            I => \N__4664\
        );

    \I__554\ : InMux
    port map (
            O => \N__4676\,
            I => \N__4661\
        );

    \I__553\ : InMux
    port map (
            O => \N__4673\,
            I => \N__4658\
        );

    \I__552\ : InMux
    port map (
            O => \N__4672\,
            I => \N__4655\
        );

    \I__551\ : Sp12to4
    port map (
            O => \N__4669\,
            I => \N__4644\
        );

    \I__550\ : Sp12to4
    port map (
            O => \N__4664\,
            I => \N__4644\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4661\,
            I => \N__4644\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4658\,
            I => \N__4644\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4655\,
            I => \N__4644\
        );

    \I__546\ : Odrv12
    port map (
            O => \N__4644\,
            I => \A_c_4\
        );

    \I__545\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4638\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4638\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_10\
        );

    \I__543\ : InMux
    port map (
            O => \N__4635\,
            I => \N__4632\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4632\,
            I => \N__4629\
        );

    \I__541\ : Span4Mux_h
    port map (
            O => \N__4629\,
            I => \N__4626\
        );

    \I__540\ : Span4Mux_h
    port map (
            O => \N__4626\,
            I => \N__4623\
        );

    \I__539\ : Odrv4
    port map (
            O => \N__4623\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_11\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__4620\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_9_cascade_\
        );

    \I__537\ : CascadeMux
    port map (
            O => \N__4617\,
            I => \N__4613\
        );

    \I__536\ : InMux
    port map (
            O => \N__4616\,
            I => \N__4608\
        );

    \I__535\ : InMux
    port map (
            O => \N__4613\,
            I => \N__4608\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__4608\,
            I => \N__4605\
        );

    \I__533\ : Odrv4
    port map (
            O => \N__4605\,
            I => \N_374\
        );

    \I__532\ : CascadeMux
    port map (
            O => \N__4602\,
            I => \N_401_cascade_\
        );

    \I__531\ : InMux
    port map (
            O => \N__4599\,
            I => \N__4596\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__4596\,
            I => \N_436\
        );

    \I__529\ : InMux
    port map (
            O => \N__4593\,
            I => \N__4590\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__4590\,
            I => \U409_AUTOCONFIG.N_285\
        );

    \I__527\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4584\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4584\,
            I => \U409_AUTOCONFIG.N_9\
        );

    \I__525\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4578\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4578\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0_1\
        );

    \I__523\ : InMux
    port map (
            O => \N__4575\,
            I => \N__4563\
        );

    \I__522\ : InMux
    port map (
            O => \N__4574\,
            I => \N__4563\
        );

    \I__521\ : InMux
    port map (
            O => \N__4573\,
            I => \N__4563\
        );

    \I__520\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4563\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4563\,
            I => \U409_AUTOCONFIG.N_405\
        );

    \I__518\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4557\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4557\,
            I => \N__4554\
        );

    \I__516\ : Odrv4
    port map (
            O => \N__4554\,
            I => \U409_AUTOCONFIG.LIDE_OUTc_0_1\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__4551\,
            I => \N__4548\
        );

    \I__514\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4545\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4545\,
            I => \N__4542\
        );

    \I__512\ : Odrv4
    port map (
            O => \N__4542\,
            I => \U409_AUTOCONFIG.LIDE_OUTc_0_0\
        );

    \I__511\ : InMux
    port map (
            O => \N__4539\,
            I => \N__4536\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__4536\,
            I => \U409_AUTOCONFIG.N_286\
        );

    \I__509\ : InMux
    port map (
            O => \N__4533\,
            I => \N__4521\
        );

    \I__508\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4521\
        );

    \I__507\ : InMux
    port map (
            O => \N__4531\,
            I => \N__4521\
        );

    \I__506\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4521\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4521\,
            I => \U409_AUTOCONFIG.AC_START_RNI3D7VZ0Z2\
        );

    \I__504\ : InMux
    port map (
            O => \N__4518\,
            I => \N__4515\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4515\,
            I => \U409_AUTOCONFIG.N_287\
        );

    \I__502\ : InMux
    port map (
            O => \N__4512\,
            I => \N__4508\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__4511\,
            I => \N__4505\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4508\,
            I => \N__4501\
        );

    \I__499\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4498\
        );

    \I__498\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4495\
        );

    \I__497\ : Span4Mux_v
    port map (
            O => \N__4501\,
            I => \N__4489\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__4498\,
            I => \N__4484\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4495\,
            I => \N__4484\
        );

    \I__494\ : InMux
    port map (
            O => \N__4494\,
            I => \N__4477\
        );

    \I__493\ : InMux
    port map (
            O => \N__4493\,
            I => \N__4477\
        );

    \I__492\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4477\
        );

    \I__491\ : Sp12to4
    port map (
            O => \N__4489\,
            I => \N__4470\
        );

    \I__490\ : Sp12to4
    port map (
            O => \N__4484\,
            I => \N__4470\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4477\,
            I => \N__4470\
        );

    \I__488\ : Odrv12
    port map (
            O => \N__4470\,
            I => \A_c_6\
        );

    \I__487\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4454\
        );

    \I__486\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4454\
        );

    \I__485\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4454\
        );

    \I__484\ : InMux
    port map (
            O => \N__4464\,
            I => \N__4454\
        );

    \I__483\ : InMux
    port map (
            O => \N__4463\,
            I => \N__4451\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4454\,
            I => \N__4448\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4451\,
            I => \N__4444\
        );

    \I__480\ : Span4Mux_v
    port map (
            O => \N__4448\,
            I => \N__4441\
        );

    \I__479\ : InMux
    port map (
            O => \N__4447\,
            I => \N__4438\
        );

    \I__478\ : Span12Mux_v
    port map (
            O => \N__4444\,
            I => \N__4431\
        );

    \I__477\ : Sp12to4
    port map (
            O => \N__4441\,
            I => \N__4431\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4438\,
            I => \N__4431\
        );

    \I__475\ : Odrv12
    port map (
            O => \N__4431\,
            I => \A_c_7\
        );

    \I__474\ : InMux
    port map (
            O => \N__4428\,
            I => \N__4425\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__4425\,
            I => \U409_AUTOCONFIG.N_274\
        );

    \I__472\ : CascadeMux
    port map (
            O => \N__4422\,
            I => \U409_AUTOCONFIG.N_383_cascade_\
        );

    \I__471\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4416\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4416\,
            I => \N__4413\
        );

    \I__469\ : Span4Mux_h
    port map (
            O => \N__4413\,
            I => \N__4410\
        );

    \I__468\ : Sp12to4
    port map (
            O => \N__4410\,
            I => \N__4407\
        );

    \I__467\ : Odrv12
    port map (
            O => \N__4407\,
            I => \TT_c_0\
        );

    \I__466\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4401\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4401\,
            I => \N__4398\
        );

    \I__464\ : Span12Mux_h
    port map (
            O => \N__4398\,
            I => \N__4395\
        );

    \I__463\ : Odrv12
    port map (
            O => \N__4395\,
            I => \TT_c_1\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__4392\,
            I => \N__4389\
        );

    \I__461\ : InMux
    port map (
            O => \N__4389\,
            I => \N__4386\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4386\,
            I => \U409_ADDRESS_DECODE.N_345\
        );

    \I__459\ : InMux
    port map (
            O => \N__4383\,
            I => \N__4380\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4380\,
            I => \U409_ADDRESS_DECODE.N_344\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__4377\,
            I => \U409_AUTOCONFIG.N_288_cascade_\
        );

    \I__456\ : InMux
    port map (
            O => \N__4374\,
            I => \N__4371\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4371\,
            I => \N__4368\
        );

    \I__454\ : Odrv4
    port map (
            O => \N__4368\,
            I => \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_a2Z0Z_1\
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__4365\,
            I => \U409_AUTOCONFIG.N_405_cascade_\
        );

    \I__452\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4354\
        );

    \I__451\ : InMux
    port map (
            O => \N__4361\,
            I => \N__4354\
        );

    \I__450\ : InMux
    port map (
            O => \N__4360\,
            I => \N__4351\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__4359\,
            I => \N__4348\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4354\,
            I => \N__4345\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__4351\,
            I => \N__4342\
        );

    \I__446\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4339\
        );

    \I__445\ : Odrv4
    port map (
            O => \N__4345\,
            I => \U409_AUTOCONFIG.N_414\
        );

    \I__444\ : Odrv4
    port map (
            O => \N__4342\,
            I => \U409_AUTOCONFIG.N_414\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4339\,
            I => \U409_AUTOCONFIG.N_414\
        );

    \I__442\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4328\
        );

    \I__441\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4325\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4328\,
            I => \U409_AUTOCONFIG.N_373\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4325\,
            I => \U409_AUTOCONFIG.N_373\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__4320\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_2_3_0_cascade_\
        );

    \I__437\ : InMux
    port map (
            O => \N__4317\,
            I => \N__4314\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4314\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0_0\
        );

    \I__435\ : InMux
    port map (
            O => \N__4311\,
            I => \N__4305\
        );

    \I__434\ : InMux
    port map (
            O => \N__4310\,
            I => \N__4305\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__4305\,
            I => \U409_AUTOCONFIG.N_269\
        );

    \I__432\ : InMux
    port map (
            O => \N__4302\,
            I => \N__4299\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__4299\,
            I => \N__4295\
        );

    \I__430\ : InMux
    port map (
            O => \N__4298\,
            I => \N__4292\
        );

    \I__429\ : Odrv4
    port map (
            O => \N__4295\,
            I => \U409_AUTOCONFIG.N_370\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__4292\,
            I => \U409_AUTOCONFIG.N_370\
        );

    \I__427\ : CascadeMux
    port map (
            O => \N__4287\,
            I => \U409_AUTOCONFIG.N_195_cascade_\
        );

    \I__426\ : InMux
    port map (
            O => \N__4284\,
            I => \N__4281\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__4281\,
            I => \N__4277\
        );

    \I__424\ : InMux
    port map (
            O => \N__4280\,
            I => \N__4274\
        );

    \I__423\ : Odrv4
    port map (
            O => \N__4277\,
            I => \U409_AUTOCONFIG.N_383\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4274\,
            I => \U409_AUTOCONFIG.N_383\
        );

    \I__421\ : CascadeMux
    port map (
            O => \N__4269\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_8_cascade_\
        );

    \I__420\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4262\
        );

    \I__419\ : InMux
    port map (
            O => \N__4265\,
            I => \N__4259\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__4262\,
            I => \N__4254\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__4259\,
            I => \N__4254\
        );

    \I__416\ : Span4Mux_v
    port map (
            O => \N__4254\,
            I => \N__4251\
        );

    \I__415\ : Span4Mux_v
    port map (
            O => \N__4251\,
            I => \N__4248\
        );

    \I__414\ : Span4Mux_h
    port map (
            O => \N__4248\,
            I => \N__4245\
        );

    \I__413\ : Odrv4
    port map (
            O => \N__4245\,
            I => \A_c_24\
        );

    \I__412\ : CascadeMux
    port map (
            O => \N__4242\,
            I => \N__4239\
        );

    \I__411\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4236\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__4236\,
            I => \U409_AUTOCONFIG.N_270\
        );

    \I__409\ : InMux
    port map (
            O => \N__4233\,
            I => \N__4230\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__4230\,
            I => \U409_AUTOCONFIG.N_271\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__4227\,
            I => \U409_AUTOCONFIG.N_433_cascade_\
        );

    \I__406\ : InMux
    port map (
            O => \N__4224\,
            I => \N__4221\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__4221\,
            I => \U409_AUTOCONFIG.N_433\
        );

    \I__404\ : CascadeMux
    port map (
            O => \N__4218\,
            I => \N__4215\
        );

    \I__403\ : InMux
    port map (
            O => \N__4215\,
            I => \N__4209\
        );

    \I__402\ : InMux
    port map (
            O => \N__4214\,
            I => \N__4209\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__4209\,
            I => \N__4206\
        );

    \I__400\ : Span4Mux_v
    port map (
            O => \N__4206\,
            I => \N__4203\
        );

    \I__399\ : Sp12to4
    port map (
            O => \N__4203\,
            I => \N__4200\
        );

    \I__398\ : Odrv12
    port map (
            O => \N__4200\,
            I => \A_c_25\
        );

    \I__397\ : InMux
    port map (
            O => \N__4197\,
            I => \N__4191\
        );

    \I__396\ : InMux
    port map (
            O => \N__4196\,
            I => \N__4191\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4191\,
            I => \N__4188\
        );

    \I__394\ : Span4Mux_v
    port map (
            O => \N__4188\,
            I => \N__4185\
        );

    \I__393\ : Span4Mux_h
    port map (
            O => \N__4185\,
            I => \N__4182\
        );

    \I__392\ : Odrv4
    port map (
            O => \N__4182\,
            I => \A_c_27\
        );

    \I__391\ : CascadeMux
    port map (
            O => \N__4179\,
            I => \N__4175\
        );

    \I__390\ : InMux
    port map (
            O => \N__4178\,
            I => \N__4170\
        );

    \I__389\ : InMux
    port map (
            O => \N__4175\,
            I => \N__4170\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__4170\,
            I => \N__4167\
        );

    \I__387\ : Span4Mux_v
    port map (
            O => \N__4167\,
            I => \N__4164\
        );

    \I__386\ : Span4Mux_v
    port map (
            O => \N__4164\,
            I => \N__4161\
        );

    \I__385\ : Sp12to4
    port map (
            O => \N__4161\,
            I => \N__4158\
        );

    \I__384\ : Odrv12
    port map (
            O => \N__4158\,
            I => \A_c_26\
        );

    \I__383\ : IoInMux
    port map (
            O => \N__4155\,
            I => \N__4152\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__4152\,
            I => \N__4149\
        );

    \I__381\ : Span4Mux_s2_h
    port map (
            O => \N__4149\,
            I => \N__4146\
        );

    \I__380\ : Sp12to4
    port map (
            O => \N__4146\,
            I => \N__4143\
        );

    \I__379\ : Span12Mux_v
    port map (
            O => \N__4143\,
            I => \N__4140\
        );

    \I__378\ : Span12Mux_v
    port map (
            O => \N__4140\,
            I => \N__4137\
        );

    \I__377\ : Odrv12
    port map (
            O => \N__4137\,
            I => \PIO_P0_c\
        );

    \I__376\ : IoInMux
    port map (
            O => \N__4134\,
            I => \N__4131\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__4131\,
            I => \N__4128\
        );

    \I__374\ : IoSpan4Mux
    port map (
            O => \N__4128\,
            I => \N__4125\
        );

    \I__373\ : Span4Mux_s2_h
    port map (
            O => \N__4125\,
            I => \N__4122\
        );

    \I__372\ : Sp12to4
    port map (
            O => \N__4122\,
            I => \N__4119\
        );

    \I__371\ : Span12Mux_v
    port map (
            O => \N__4119\,
            I => \N__4116\
        );

    \I__370\ : Span12Mux_v
    port map (
            O => \N__4116\,
            I => \N__4113\
        );

    \I__369\ : Odrv12
    port map (
            O => \N__4113\,
            I => \PIO_S0_c\
        );

    \I__368\ : ClkMux
    port map (
            O => \N__4110\,
            I => \N__4077\
        );

    \I__367\ : ClkMux
    port map (
            O => \N__4109\,
            I => \N__4077\
        );

    \I__366\ : ClkMux
    port map (
            O => \N__4108\,
            I => \N__4077\
        );

    \I__365\ : ClkMux
    port map (
            O => \N__4107\,
            I => \N__4077\
        );

    \I__364\ : ClkMux
    port map (
            O => \N__4106\,
            I => \N__4077\
        );

    \I__363\ : ClkMux
    port map (
            O => \N__4105\,
            I => \N__4077\
        );

    \I__362\ : ClkMux
    port map (
            O => \N__4104\,
            I => \N__4077\
        );

    \I__361\ : ClkMux
    port map (
            O => \N__4103\,
            I => \N__4077\
        );

    \I__360\ : ClkMux
    port map (
            O => \N__4102\,
            I => \N__4077\
        );

    \I__359\ : ClkMux
    port map (
            O => \N__4101\,
            I => \N__4077\
        );

    \I__358\ : ClkMux
    port map (
            O => \N__4100\,
            I => \N__4077\
        );

    \I__357\ : GlobalMux
    port map (
            O => \N__4077\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            I => \N__4101\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__4100\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            I => \N__4107\
        );

    \INVU409_TRANSFER_ACK.TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            I => \N__4104\
        );

    \INVU409_TRANSFER_ACK.TACK_OUTnC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            I => \N__4102\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\,
            I => \N__4106\
        );

    \INVU409_AUTOCONFIG.CONFIGENnC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            I => \N__8329\
        );

    \INVU409_TRANSFER_ACK.CIA_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            I => \N__4103\
        );

    \INVU409_AUTOCONFIG.ATA_BASE_ness_3C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.ATA_BASE_ness_3C_net\,
            I => \N__8344\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            I => \N__4108\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            I => \N__4105\
        );

    \INVU409_AUTOCONFIG.ATA_BASE_ness_4C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net\,
            I => \N__8346\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            I => \N__4110\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            I => \N__4109\
        );

    \INVU409_AUTOCONFIG.AC_TACKC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.AC_TACKC_net\,
            I => \N__8342\
        );

    \INVU409_AUTOCONFIG.BRIDGE_BASE_3C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net\,
            I => \N__8349\
        );

    \INVU409_AUTOCONFIG.STATE_0C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.STATE_0C_net\,
            I => \N__8345\
        );

    \INVU409_AUTOCONFIG.LIDE_OUT_0C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            I => \N__8347\
        );

    \INVU409_AUTOCONFIG.BRIDGE_OUT_3C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            I => \N__8350\
        );

    \IN_MUX_bfv_13_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_6_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_14_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_5_0_\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_9_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9009\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_o2_4_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4214\,
            in1 => \N__4196\,
            in2 => \N__4179\,
            in3 => \N__4265\,
            lcout => \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_o2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_8_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5684\,
            in1 => \N__5614\,
            in2 => \N__4218\,
            in3 => \N__5397\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_11_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4197\,
            in1 => \N__4178\,
            in2 => \N__4269\,
            in3 => \N__4266\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__4233\,
            in1 => \N__9169\,
            in2 => \N__4242\,
            in3 => \N__4317\,
            lcout => \U409_AUTOCONFIG.N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4725\,
            in1 => \N__4840\,
            in2 => \_gnd_net_\,
            in3 => \N__4360\,
            lcout => \U409_AUTOCONFIG.N_270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4302\,
            in1 => \N__4332\,
            in2 => \N__4741\,
            in3 => \N__7280\,
            lcout => \U409_AUTOCONFIG.N_271\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__4310\,
            in1 => \N__4834\,
            in2 => \N__4359\,
            in3 => \N__7329\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_5_0_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__4835\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5166\,
            lcout => \U409_AUTOCONFIG.N_373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_7_0_71_i_i_0_a2_1_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__5167\,
            in1 => \N__4836\,
            in2 => \N__4742\,
            in3 => \N__7331\,
            lcout => \U409_AUTOCONFIG.N_433\,
            ltout => \U409_AUTOCONFIG.N_433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__4298\,
            in1 => \_gnd_net_\,
            in2 => \N__4227\,
            in3 => \N__4284\,
            lcout => \U409_AUTOCONFIG.N_285\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__5248\,
            in1 => \N__4224\,
            in2 => \N__4743\,
            in3 => \N__7333\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTc_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_4_0_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7330\,
            in1 => \N__4447\,
            in2 => \N__4740\,
            in3 => \N__5247\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_2_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__4311\,
            in1 => \N__4331\,
            in2 => \N__4320\,
            in3 => \N__4512\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__7332\,
            in1 => \N__4732\,
            in2 => \N__4842\,
            in3 => \N__5168\,
            lcout => \U409_AUTOCONFIG.N_286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_0_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4280\,
            in1 => \N__4464\,
            in2 => \N__5227\,
            in3 => \N__4492\,
            lcout => \U409_AUTOCONFIG.N_269\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_7_0_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5154\,
            in1 => \N__4466\,
            in2 => \N__5228\,
            in3 => \N__4494\,
            lcout => \U409_AUTOCONFIG.N_414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_4_0_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5204\,
            in1 => \N__4465\,
            in2 => \_gnd_net_\,
            in3 => \N__4493\,
            lcout => \U409_AUTOCONFIG.N_370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_o2_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110001"
        )
    port map (
            in0 => \N__4809\,
            in1 => \N__7328\,
            in2 => \N__5229\,
            in3 => \N__4721\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.N_195_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_a2_1_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__4467\,
            in1 => \_gnd_net_\,
            in2 => \N__4287\,
            in3 => \N__4504\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_0_0_a2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__7327\,
            in1 => \N__4817\,
            in2 => \N__4692\,
            in3 => \N__5152\,
            lcout => \U409_AUTOCONFIG.N_274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_6_0_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7326\,
            in1 => \N__4816\,
            in2 => \_gnd_net_\,
            in3 => \N__4672\,
            lcout => \U409_AUTOCONFIG.N_383\,
            ltout => \U409_AUTOCONFIG.N_383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__5151\,
            in1 => \N__4428\,
            in2 => \N__4422\,
            in3 => \N__5249\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTc_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_4_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__6723\,
            in1 => \N__6921\,
            in2 => \N__7700\,
            in3 => \N__7804\,
            lcout => \U409_ADDRESS_DECODE.N_344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_2_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__6722\,
            in1 => \N__6920\,
            in2 => \N__7699\,
            in3 => \N__6117\,
            lcout => \U409_ADDRESS_DECODE.N_345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_10_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4419\,
            in1 => \N__4404\,
            in2 => \N__9177\,
            in3 => \N__6615\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_1_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__7937\,
            in1 => \N__5067\,
            in2 => \N__4392\,
            in3 => \N__4383\,
            lcout => \N_434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000100000"
        )
    port map (
            in0 => \N__4362\,
            in1 => \N__4841\,
            in2 => \N__7325\,
            in3 => \N__4739\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.N_288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110000001000"
        )
    port map (
            in0 => \N__4575\,
            in1 => \N__9170\,
            in2 => \N__4377\,
            in3 => \N__5918\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_RNIJJLA1_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7121\,
            in1 => \N__5556\,
            in2 => \N__4902\,
            in3 => \N__4877\,
            lcout => \U409_AUTOCONFIG.N_405\,
            ltout => \U409_AUTOCONFIG.N_405_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_RNI3D7V2_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111010101"
        )
    port map (
            in0 => \N__9163\,
            in1 => \N__4374\,
            in2 => \N__4365\,
            in3 => \N__4361\,
            lcout => \U409_AUTOCONFIG.AC_START_RNI3D7VZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011000000"
        )
    port map (
            in0 => \N__4593\,
            in1 => \N__9168\,
            in2 => \N__6410\,
            in3 => \N__4574\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__4573\,
            in1 => \N__4587\,
            in2 => \N__9178\,
            in3 => \N__4952\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011000000"
        )
    port map (
            in0 => \N__4581\,
            in1 => \N__9167\,
            in2 => \N__5525\,
            in3 => \N__4572\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__4560\,
            in1 => \N__4934\,
            in2 => \N__5103\,
            in3 => \N__4530\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            ce => 'H',
            sr => \N__9424\
        );

    \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100000010"
        )
    port map (
            in0 => \N__4531\,
            in1 => \N__4863\,
            in2 => \N__4551\,
            in3 => \N__5498\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            ce => 'H',
            sr => \N__9424\
        );

    \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__4539\,
            in1 => \N__6389\,
            in2 => \N__4854\,
            in3 => \N__4532\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            ce => 'H',
            sr => \N__9424\
        );

    \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__4533\,
            in1 => \N__4518\,
            in2 => \N__5942\,
            in3 => \N__4853\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            ce => 'H',
            sr => \N__9424\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4737\,
            in1 => \N__4811\,
            in2 => \N__7363\,
            in3 => \N__5165\,
            lcout => \U409_AUTOCONFIG.N_287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_STATE_1_0_a2_0_2_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5232\,
            in1 => \N__5262\,
            in2 => \N__4511\,
            in3 => \N__4463\,
            lcout => \U409_AUTOCONFIG.un1_STATE_1_0_a2_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4736\,
            in1 => \N__4810\,
            in2 => \N__7362\,
            in3 => \N__5230\,
            lcout => \U409_AUTOCONFIG.N_273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_129_i_i_0_a2_0_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4738\,
            in1 => \N__4812\,
            in2 => \N__7364\,
            in3 => \N__5231\,
            lcout => \U409_AUTOCONFIG.N_400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_2_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__6112\,
            in1 => \N__6893\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_a2_3_0_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4830\,
            in2 => \_gnd_net_\,
            in3 => \N__4676\,
            lcout => \U409_AUTOCONFIG.N_360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14_9_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6699\,
            in1 => \N__7839\,
            in2 => \N__5451\,
            in3 => \N__4616\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_0_14Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__4641\,
            in1 => \N__4635\,
            in2 => \N__4620\,
            in3 => \N__4599\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_i_a2_1_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5018\,
            in1 => \N__5054\,
            in2 => \N__4617\,
            in3 => \N__9270\,
            lcout => \N_401\,
            ltout => \N_401_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6698\,
            in1 => \N__6735\,
            in2 => \N__4602\,
            in3 => \N__6590\,
            lcout => \N_436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_0_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__9159\,
            in1 => \N__5538\,
            in2 => \_gnd_net_\,
            in3 => \N__4972\,
            lcout => \N_348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.N_265_i_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__5536\,
            in1 => \N__9158\,
            in2 => \N__4973\,
            in3 => \N__6842\,
            lcout => \N_265_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_0_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111011"
        )
    port map (
            in0 => \N__5537\,
            in1 => \N__5011\,
            in2 => \N__4974\,
            in3 => \N__5042\,
            lcout => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__4953\,
            in1 => \N__6376\,
            in2 => \N__4941\,
            in3 => \N__7471\,
            lcout => \N_124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8438\,
            in1 => \N__6318\,
            in2 => \_gnd_net_\,
            in3 => \N__7201\,
            lcout => \U409_AUTOCONFIG.AC_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNI2IAK1_0_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5172\,
            in1 => \N__7140\,
            in2 => \N__4911\,
            in3 => \N__5557\,
            lcout => \U409_AUTOCONFIG.un1_STATE_1_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_0_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5558\,
            in1 => \N__4895\,
            in2 => \N__9179\,
            in3 => \N__4878\,
            lcout => \U409_AUTOCONFIG.STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_5_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6932\,
            in1 => \N__6775\,
            in2 => \_gnd_net_\,
            in3 => \N__6088\,
            lcout => OPEN,
            ltout => \N_354_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_DATA_BUFFERS.un1_BUFENn_i_a2_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9230\,
            in1 => \N__6448\,
            in2 => \N__4866\,
            in3 => \N__9308\,
            lcout => \N_356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_1_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7787\,
            in1 => \N__7936\,
            in2 => \_gnd_net_\,
            in3 => \N__7718\,
            lcout => \N_351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.D_1_i_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6661\,
            in1 => \N__7135\,
            in2 => \N__6606\,
            in3 => \N__7059\,
            lcout => \D_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_1_i_a2_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6662\,
            in1 => \N__6586\,
            in2 => \_gnd_net_\,
            in3 => \N__7060\,
            lcout => \N_357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_DATA_BUFFERS.un1_BUFENn_i_a2_0_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7962\,
            in1 => \N__7802\,
            in2 => \N__6607\,
            in3 => \N__7067\,
            lcout => \N_297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5286\,
            in1 => \N__5261\,
            in2 => \N__5250\,
            in3 => \N__5153\,
            lcout => \U409_AUTOCONFIG.N_276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6006\,
            in2 => \_gnd_net_\,
            in3 => \N__5974\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_i_1_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__6736\,
            in1 => \N__7857\,
            in2 => \N__6694\,
            in3 => \N__8417\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.PORTSIZE_iZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_i_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__6854\,
            in1 => \N__9271\,
            in2 => \N__5088\,
            in3 => \N__8039\,
            lcout => \N_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_3_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6116\,
            in1 => \N__6737\,
            in2 => \N__6931\,
            in3 => \N__6519\,
            lcout => \U409_ADDRESS_DECODE.N_343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_x2_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__5055\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5019\,
            lcout => \N_156_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_o2_5_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5691\,
            in1 => \N__5625\,
            in2 => \N__5395\,
            in3 => \N__5447\,
            lcout => \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_o2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__5526\,
            in1 => \N__5505\,
            in2 => \N__6378\,
            in3 => \N__7470\,
            lcout => \N_126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7646\,
            in1 => \N__5651\,
            in2 => \N__7578\,
            in3 => \N__5574\,
            lcout => \BRIDGE_BASE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net\,
            ce => 'H',
            sr => \N__9425\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__5572\,
            in1 => \N__7644\,
            in2 => \N__5822\,
            in3 => \N__5408\,
            lcout => \BRIDGE_BASE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net\,
            ce => 'H',
            sr => \N__9425\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7643\,
            in1 => \N__5345\,
            in2 => \N__5871\,
            in3 => \N__5571\,
            lcout => \BRIDGE_BASE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net\,
            ce => 'H',
            sr => \N__9425\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7645\,
            in1 => \N__5636\,
            in2 => \N__6191\,
            in3 => \N__5573\,
            lcout => \BRIDGE_BASE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net\,
            ce => 'H',
            sr => \N__9425\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__5334\,
            in1 => \N__5580\,
            in2 => \N__6495\,
            in3 => \N__9247\,
            lcout => \N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__5446\,
            in1 => \N__5409\,
            in2 => \N__5396\,
            in3 => \N__5346\,
            lcout => \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIOE6K2_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011101110"
        )
    port map (
            in0 => \N__7392\,
            in1 => \N__9429\,
            in2 => \N__7464\,
            in3 => \N__7285\,
            lcout => \U409_AUTOCONFIG.un1_STATE_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0_1_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__5683\,
            in1 => \N__5652\,
            in2 => \N__5640\,
            in3 => \N__5624\,
            lcout => \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNI25A42_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__7284\,
            in1 => \N__7443\,
            in2 => \_gnd_net_\,
            in3 => \N__7391\,
            lcout => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_o2dup_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__9136\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7202\,
            lcout => \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_o2dupZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_TACK_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5559\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \AC_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.AC_TACKC_net\,
            ce => 'H',
            sr => \N__9418\
        );

    \U409_AUTOCONFIG.BRIDGE_CONF_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010101010"
        )
    port map (
            in0 => \N__6362\,
            in1 => \N__7393\,
            in2 => \N__7365\,
            in3 => \N__7451\,
            lcout => \U409_AUTOCONFIG.BRIDGE_CONFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.AC_TACKC_net\,
            ce => 'H',
            sr => \N__9418\
        );

    \U409_AUTOCONFIG.LIDE_CONF_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__7346\,
            in1 => \N__7394\,
            in2 => \_gnd_net_\,
            in3 => \N__7450\,
            lcout => \U409_AUTOCONFIG.LIDE_CONFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.AC_TACKC_net\,
            ce => 'H',
            sr => \N__9418\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__7041\,
            in1 => \N__7008\,
            in2 => \_gnd_net_\,
            in3 => \N__6987\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__6810\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__5771\,
            in1 => \N__5790\,
            in2 => \N__5745\,
            in3 => \N__6262\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__6810\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5741\,
            in1 => \N__5789\,
            in2 => \_gnd_net_\,
            in3 => \N__6261\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__6810\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__7035\,
            in1 => \N__6001\,
            in2 => \N__5733\,
            in3 => \N__5796\,
            lcout => \U409_TRANSFER_ACK.N_237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__5969\,
            in1 => \N__5787\,
            in2 => \N__5714\,
            in3 => \N__5767\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5788\,
            in1 => \N__5970\,
            in2 => \N__5772\,
            in3 => \N__5706\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6002\,
            in1 => \N__7036\,
            in2 => \N__5754\,
            in3 => \N__5732\,
            lcout => \U409_TRANSFER_ACK.N_268\,
            ltout => \U409_TRANSFER_ACK.N_268_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011111111"
        )
    port map (
            in0 => \N__8380\,
            in1 => \N__6306\,
            in2 => \N__5751\,
            in3 => \N__6221\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7006\,
            in1 => \N__6011\,
            in2 => \N__5715\,
            in3 => \N__5976\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__7037\,
            in1 => \N__6984\,
            in2 => \N__5748\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7005\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6983\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__6952\,
            in1 => \_gnd_net_\,
            in2 => \N__6012\,
            in3 => \N__6256\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__6808\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__6956\,
            in1 => \N__5721\,
            in2 => \N__6264\,
            in3 => \N__5713\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__6808\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__6007\,
            in1 => \N__5975\,
            in2 => \N__6957\,
            in3 => \N__6260\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__6808\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_i_a2_0_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7952\,
            in1 => \N__6515\,
            in2 => \N__7874\,
            in3 => \N__7835\,
            lcout => \N_339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNISS061_3_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__5946\,
            in1 => \N__5925\,
            in2 => \N__7479\,
            in3 => \N__6377\,
            lcout => \N_130\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_2_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__6783\,
            in1 => \N__5879\,
            in2 => \N__6939\,
            in3 => \N__5888\,
            lcout => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.ATA_BASE_ness_4_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__5889\,
            in1 => \N__5870\,
            in2 => \N__7639\,
            in3 => \N__7491\,
            lcout => \ATA_BASE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net\,
            ce => \N__7505\,
            sr => \N__9420\
        );

    \U409_AUTOCONFIG.ATA_BASE_ness_5_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__7492\,
            in1 => \N__7623\,
            in2 => \N__5835\,
            in3 => \N__5880\,
            lcout => \ATA_BASE_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net\,
            ce => \N__7505\,
            sr => \N__9420\
        );

    \U409_AUTOCONFIG.ATA_BASE_ness_0_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__7367\,
            in1 => \N__5869\,
            in2 => \N__7638\,
            in3 => \N__6138\,
            lcout => \ATA_BASE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net\,
            ce => \N__7505\,
            sr => \N__9420\
        );

    \U409_AUTOCONFIG.ATA_BASE_ness_1_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__5831\,
            in1 => \N__7368\,
            in2 => \N__6153\,
            in3 => \N__7618\,
            lcout => \ATA_BASE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net\,
            ce => \N__7505\,
            sr => \N__9420\
        );

    \U409_AUTOCONFIG.ATA_BASE_ness_6_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__7624\,
            in1 => \N__7493\,
            in2 => \N__6210\,
            in3 => \N__6165\,
            lcout => \ATA_BASE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net\,
            ce => \N__7505\,
            sr => \N__9420\
        );

    \U409_AUTOCONFIG.ATA_BASE_ness_2_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__6063\,
            in1 => \N__7619\,
            in2 => \N__6209\,
            in3 => \N__7369\,
            lcout => \ATA_BASE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net\,
            ce => \N__7505\,
            sr => \N__9420\
        );

    \U409_AUTOCONFIG.ATA_BASE_ness_7_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__7625\,
            in1 => \N__7494\,
            in2 => \N__7577\,
            in3 => \N__7737\,
            lcout => \ATA_BASE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_ness_4C_net\,
            ce => \N__7505\,
            sr => \N__9420\
        );

    \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__7968\,
            in1 => \N__6164\,
            in2 => \N__6608\,
            in3 => \N__6149\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_7_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__6455\,
            in1 => \N__6137\,
            in2 => \N__6126\,
            in3 => \N__6051\,
            lcout => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_7\,
            ltout => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNO_1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6123\,
            in3 => \N__7655\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.ATA_EN_2_0_o2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001010"
        )
    port map (
            in0 => \N__9135\,
            in1 => \N__6476\,
            in2 => \N__6120\,
            in3 => \N__6045\,
            lcout => \U409_ADDRESS_DECODE.ATA_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_ATA_ENn_i_x2_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6111\,
            in2 => \_gnd_net_\,
            in3 => \N__6062\,
            lcout => \U409_ADDRESS_DECODE.N_183_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNO_0_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6029\,
            in1 => \N__6038\,
            in2 => \N__7134\,
            in3 => \N__7182\,
            lcout => \U409_ADDRESS_DECODE.ATA_EN_2_0_o2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_ATA_ENn_i_0_3_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6039\,
            in1 => \N__6030\,
            in2 => \N__6504\,
            in3 => \N__6494\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNIU5437_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111111"
        )
    port map (
            in0 => \N__7656\,
            in1 => \_gnd_net_\,
            in2 => \N__6480\,
            in3 => \N__6477\,
            lcout => \N_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_3_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6782\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6456\,
            lcout => \N_422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_3_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6321\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8382\,
            lcout => \U409_TRANSFER_ACK.N_381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6320\,
            in1 => \N__8381\,
            in2 => \N__8129\,
            in3 => \N__8144\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIQQ061_2_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__6414\,
            in1 => \N__6393\,
            in2 => \N__7469\,
            in3 => \N__6363\,
            lcout => \N_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110000110011"
        )
    port map (
            in0 => \N__6319\,
            in1 => \N__7040\,
            in2 => \N__8385\,
            in3 => \N__6233\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__6809\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7039\,
            in1 => \N__6986\,
            in2 => \_gnd_net_\,
            in3 => \N__6263\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__6809\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__6234\,
            in1 => \N__7161\,
            in2 => \_gnd_net_\,
            in3 => \N__6222\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__6809\
        );

    \U409_ADDRESS_DECODE.D_IN_0_a2_0_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__7139\,
            in1 => \N__6612\,
            in2 => \N__7074\,
            in3 => \N__6695\,
            lcout => \N_361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7038\,
            in1 => \N__7007\,
            in2 => \_gnd_net_\,
            in3 => \N__6985\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__9328\,
            in1 => \N__9380\,
            in2 => \N__6911\,
            in3 => \N__7811\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.N_346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__6900\,
            in1 => \N__6697\,
            in2 => \N__6861\,
            in3 => \N__6774\,
            lcout => \U409_TRANSFER_ACK.N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a2_1_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6764\,
            in1 => \N__7964\,
            in2 => \_gnd_net_\,
            in3 => \N__7711\,
            lcout => \N_429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_DATA_BUFFERS.un1_BUFENn_i_o2_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__6858\,
            in1 => \N__9381\,
            in2 => \N__9335\,
            in3 => \N__9236\,
            lcout => \N_190\,
            ltout => \N_190_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001111111111"
        )
    port map (
            in0 => \N__9302\,
            in1 => \N__9180\,
            in2 => \N__6831\,
            in3 => \N__6828\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.N_436_i_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__6763\,
            in1 => \N__6696\,
            in2 => \N__7881\,
            in3 => \N__6613\,
            lcout => \N_436_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_i_a2_2_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7812\,
            in1 => \N__6614\,
            in2 => \_gnd_net_\,
            in3 => \N__7701\,
            lcout => \N_431\,
            ltout => \N_431_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7963\,
            in1 => \N__7870\,
            in2 => \N__7842\,
            in3 => \N__7828\,
            lcout => \U409_CIA.VMA_3_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2_5_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__7803\,
            in1 => \N__7736\,
            in2 => \N__7725\,
            in3 => \N__7523\,
            lcout => \U409_ADDRESS_DECODE.un1_ATA_ENn_i_o2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.ATA_BASE_ness_3_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__7524\,
            in1 => \N__7370\,
            in2 => \N__7647\,
            in3 => \N__7558\,
            lcout => \ATA_BASE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_ness_3C_net\,
            ce => \N__7515\,
            sr => \N__9419\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNI0JVF_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7371\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7475\,
            lcout => \U409_AUTOCONFIG.N_172\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000101010"
        )
    port map (
            in0 => \N__8091\,
            in1 => \N__8916\,
            in2 => \N__8883\,
            in3 => \N__8268\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__9417\
        );

    \U409_AUTOCONFIG.CONFIGENn_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__7468\,
            in1 => \N__7398\,
            in2 => \N__7366\,
            in3 => \N__7188\,
            lcout => \CONFIGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            ce => 'H',
            sr => \N__9416\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7160\,
            in2 => \_gnd_net_\,
            in3 => \N__8105\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7149\,
            in1 => \N__8078\,
            in2 => \N__8094\,
            in3 => \N__8090\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011010000"
        )
    port map (
            in0 => \N__8520\,
            in1 => \N__8551\,
            in2 => \N__8592\,
            in3 => \N__8632\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__9414\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010111010"
        )
    port map (
            in0 => \N__8079\,
            in1 => \N__8552\,
            in2 => \N__8727\,
            in3 => \N__8633\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__9414\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8067\,
            in1 => \N__9304\,
            in2 => \N__8634\,
            in3 => \N__9246\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9303\,
            in1 => \N__8066\,
            in2 => \N__9249\,
            in3 => \N__8058\,
            lcout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8545\,
            in2 => \_gnd_net_\,
            in3 => \N__8625\,
            lcout => \U409_TRANSFER_ACK.N_380\,
            ltout => \U409_TRANSFER_ACK.N_380_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011101110"
        )
    port map (
            in0 => \N__8702\,
            in1 => \N__8585\,
            in2 => \N__8052\,
            in3 => \N__8517\,
            lcout => \U409_TRANSFER_ACK.ROMENn_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_DATA_BUFFERS.N_94_i_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__8049\,
            in1 => \N__9301\,
            in2 => \_gnd_net_\,
            in3 => \N__8043\,
            lcout => \N_94_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8007\,
            in2 => \_gnd_net_\,
            in3 => \N__8277\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS1n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_3_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8908\,
            in2 => \_gnd_net_\,
            in3 => \N__8873\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8787\,
            in1 => \N__8373\,
            in2 => \N__8271\,
            in3 => \N__8807\,
            lcout => \U409_TRANSFER_ACK.N_293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8806\,
            in1 => \N__8786\,
            in2 => \N__8384\,
            in3 => \N__8909\,
            lcout => \U409_TRANSFER_ACK.N_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100100111"
        )
    port map (
            in0 => \N__8178\,
            in1 => \N__8221\,
            in2 => \N__8206\,
            in3 => \N__8161\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__8222\,
            in1 => \_gnd_net_\,
            in2 => \N__8262\,
            in3 => \N__9107\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001000100"
        )
    port map (
            in0 => \N__8180\,
            in1 => \N__9105\,
            in2 => \N__8208\,
            in3 => \N__8162\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__8179\,
            in1 => \_gnd_net_\,
            in2 => \N__8207\,
            in3 => \N__9106\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000001110001"
        )
    port map (
            in0 => \N__8205\,
            in1 => \N__8181\,
            in2 => \N__8464\,
            in3 => \N__8163\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            ce => 'H',
            sr => \N__9415\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__8698\,
            in1 => \N__8148\,
            in2 => \N__8133\,
            in3 => \N__8106\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            ce => 'H',
            sr => \N__9415\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010010"
        )
    port map (
            in0 => \N__8516\,
            in1 => \N__8626\,
            in2 => \N__8591\,
            in3 => \N__8546\,
            lcout => \U409_TRANSFER_ACK.N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8581\,
            in2 => \_gnd_net_\,
            in3 => \N__8515\,
            lcout => \U409_TRANSFER_ACK.N_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__8718\,
            in1 => \N__8712\,
            in2 => \N__8706\,
            in3 => \N__8518\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__9412\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8547\,
            in2 => \_gnd_net_\,
            in3 => \N__8631\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__9412\
        );

    \U409_TRANSFER_ACK.ROMENn_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011000011111010"
        )
    port map (
            in0 => \N__8586\,
            in1 => \N__8676\,
            in2 => \N__8651\,
            in3 => \N__8670\,
            lcout => \ROMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__9412\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101110100000"
        )
    port map (
            in0 => \N__8630\,
            in1 => \N__8590\,
            in2 => \N__8553\,
            in3 => \N__8519\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__9412\
        );

    \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__8465\,
            in1 => \N__8442\,
            in2 => \_gnd_net_\,
            in3 => \N__8421\,
            lcout => \TCIn_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8383\,
            lcout => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNI692L_0_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9696\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9044\,
            lcout => \CIA_ENABLE\,
            ltout => \CIA_ENABLE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8772\,
            in3 => \N__8769\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS0n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__9878\,
            in1 => \N__9801\,
            in2 => \N__8955\,
            in3 => \N__9849\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__9471\,
            in1 => \N__9504\,
            in2 => \N__9528\,
            in3 => \N__9452\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => \U409_TICK.TICK603_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9877\,
            in1 => \N__9848\,
            in2 => \N__8733\,
            in3 => \N__9438\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9486\,
            in1 => \N__8979\,
            in2 => \N__9000\,
            in3 => \N__9647\,
            lcout => \U409_TICK.TICK603_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8999\,
            in2 => \_gnd_net_\,
            in3 => \N__9978\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_1_1_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8821\,
            in2 => \_gnd_net_\,
            in3 => \N__8844\,
            lcout => \U409_TRANSFER_ACK.N_223\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_4_0_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__8845\,
            in1 => \_gnd_net_\,
            in2 => \N__8828\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.m12_i_a2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_2_0_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__8875\,
            in1 => \N__8934\,
            in2 => \N__8730\,
            in3 => \N__8912\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.m12_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__9070\,
            in1 => \N__8853\,
            in2 => \N__8943\,
            in3 => \N__8940\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8785\,
            in2 => \_gnd_net_\,
            in3 => \N__8805\,
            lcout => \U409_TRANSFER_ACK.N_191\,
            ltout => \U409_TRANSFER_ACK.N_191_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111011001"
        )
    port map (
            in0 => \N__8911\,
            in1 => \N__8876\,
            in2 => \N__8928\,
            in3 => \N__8925\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.i5_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8919\,
            in3 => \N__9071\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__8846\,
            in1 => \N__8910\,
            in2 => \N__8829\,
            in3 => \N__8874\,
            lcout => \U409_TRANSFER_ACK.N_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9072\,
            in2 => \_gnd_net_\,
            in3 => \N__9689\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__9413\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9548\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__9413\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8847\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__9413\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8808\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__9413\
        );

    \U409_ADDRESS_DECODE.N_264_i_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__9365\,
            in1 => \N__9339\,
            in2 => \N__9312\,
            in3 => \N__9248\,
            lcout => \N_264_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9099\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8990\,
            in2 => \N__9977\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_6_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8978\,
            in2 => \_gnd_net_\,
            in3 => \N__8967\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__10648\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9617\,
            in2 => \_gnd_net_\,
            in3 => \N__8964\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__10648\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9944\,
            in2 => \_gnd_net_\,
            in3 => \N__8961\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9728\,
            in2 => \_gnd_net_\,
            in3 => \N__8958\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__10648\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9914\,
            in2 => \_gnd_net_\,
            in3 => \N__8946\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9524\,
            in2 => \_gnd_net_\,
            in3 => \N__9513\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__10648\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9767\,
            in2 => \_gnd_net_\,
            in3 => \N__9510\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9932\,
            in2 => \_gnd_net_\,
            in3 => \N__9507\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9503\,
            in2 => \_gnd_net_\,
            in3 => \N__9492\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__10650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9635\,
            in2 => \_gnd_net_\,
            in3 => \N__9489\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__10650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9485\,
            in2 => \_gnd_net_\,
            in3 => \N__9474\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__10650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9470\,
            in2 => \_gnd_net_\,
            in3 => \N__9459\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__10650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9893\,
            in2 => \_gnd_net_\,
            in3 => \N__9456\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9453\,
            in3 => \N__9432\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9648\,
            in2 => \_gnd_net_\,
            in3 => \N__9651\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__9717\,
            in1 => \N__9636\,
            in2 => \N__9624\,
            in3 => \N__9606\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__9581\,
            in1 => \N__9802\,
            in2 => \N__9600\,
            in3 => \N__9847\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10348\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10283\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_2_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10344\,
            in2 => \_gnd_net_\,
            in3 => \N__10246\,
            lcout => OPEN,
            ltout => \U409_CIA.CLK_CIA6_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_0_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__10319\,
            in1 => \N__10055\,
            in2 => \N__9570\,
            in3 => \N__10371\,
            lcout => OPEN,
            ltout => \U409_CIA.CLK_CIA6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9547\,
            in2 => \N__9567\,
            in3 => \N__10359\,
            lcout => \CLK_CIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10283\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_2_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__10247\,
            in1 => \_gnd_net_\,
            in2 => \N__10353\,
            in3 => \N__10311\,
            lcout => OPEN,
            ltout => \U409_CIA.un1_CIA_CLK_COUNT_3_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_1_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__10056\,
            in1 => \N__10269\,
            in2 => \N__9531\,
            in3 => \N__10224\,
            lcout => OPEN,
            ltout => \U409_CIA.VMA_RNOZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__9711\,
            in1 => \N__9688\,
            in2 => \N__9699\,
            in3 => \N__10312\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10283\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10123\,
            in2 => \N__10527\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_5_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10142\,
            in2 => \_gnd_net_\,
            in3 => \N__9672\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__10649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10538\,
            in2 => \_gnd_net_\,
            in3 => \N__9669\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__10649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10082\,
            in2 => \_gnd_net_\,
            in3 => \N__9666\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__10649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10550\,
            in2 => \_gnd_net_\,
            in3 => \N__9663\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10418\,
            in2 => \_gnd_net_\,
            in3 => \N__9660\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10097\,
            in2 => \_gnd_net_\,
            in3 => \N__9657\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__10649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10154\,
            in2 => \_gnd_net_\,
            in3 => \N__9654\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__10649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10667\,
            in2 => \_gnd_net_\,
            in3 => \N__9753\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10475\,
            in2 => \_gnd_net_\,
            in3 => \N__9750\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__10651\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10385\,
            in2 => \_gnd_net_\,
            in3 => \N__9747\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10499\,
            in2 => \_gnd_net_\,
            in3 => \N__9744\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__10651\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10406\,
            in2 => \_gnd_net_\,
            in3 => \N__9741\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10430\,
            in2 => \_gnd_net_\,
            in3 => \N__9738\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10454\,
            in2 => \_gnd_net_\,
            in3 => \N__9735\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10110\,
            in2 => \_gnd_net_\,
            in3 => \N__9732\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10651\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__9729\,
            in1 => \N__9945\,
            in2 => \_gnd_net_\,
            in3 => \N__9972\,
            lcout => \U409_TICK.TICK603_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__9881\,
            in1 => \N__9984\,
            in2 => \N__9816\,
            in3 => \N__9846\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__9843\,
            in1 => \N__9973\,
            in2 => \N__9882\,
            in3 => \N__9813\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9879\,
            in1 => \N__9844\,
            in2 => \N__9814\,
            in3 => \N__9951\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9933\,
            in1 => \N__9768\,
            in2 => \N__9921\,
            in3 => \N__9894\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9803\,
            in1 => \N__9873\,
            in2 => \N__9903\,
            in3 => \N__9900\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9880\,
            in1 => \N__9845\,
            in2 => \N__9815\,
            in3 => \N__9774\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10349\,
            in2 => \N__10320\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10223\,
            in2 => \_gnd_net_\,
            in3 => \N__9756\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__10284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10043\,
            in1 => \N__9999\,
            in2 => \_gnd_net_\,
            in3 => \N__10071\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \N__10284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10248\,
            in2 => \_gnd_net_\,
            in3 => \N__10068\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__10284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10044\,
            in1 => \N__10268\,
            in2 => \_gnd_net_\,
            in3 => \N__10065\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            clk => \N__10284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_6_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10032\,
            in2 => \_gnd_net_\,
            in3 => \N__10062\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\,
            clk => \N__10284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_7_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10016\,
            in2 => \_gnd_net_\,
            in3 => \N__10059\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIBFRM_2_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__10267\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10222\,
            lcout => \U409_CIA.N_420\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__10012\,
            in1 => \N__10030\,
            in2 => \_gnd_net_\,
            in3 => \N__9997\,
            lcout => \U409_CIA.N_427\,
            ltout => \U409_CIA.N_427_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10316\,
            in1 => \N__10350\,
            in2 => \N__10047\,
            in3 => \N__10203\,
            lcout => \U409_CIA.CIA_CLK_COUNT11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_3_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__10245\,
            in1 => \N__10031\,
            in2 => \N__10017\,
            in3 => \N__9998\,
            lcout => OPEN,
            ltout => \U409_CIA.un1_CIA_CLK_COUNT_2_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_1_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__10317\,
            in1 => \N__10351\,
            in2 => \N__10374\,
            in3 => \N__10370\,
            lcout => \U409_CIA.CLK_CIA_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__10352\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10318\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__10266\,
            in1 => \N__10244\,
            in2 => \_gnd_net_\,
            in3 => \N__10221\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__10746\,
            in1 => \N__10772\,
            in2 => \N__10197\,
            in3 => \N__10712\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__10774\,
            in1 => \N__10172\,
            in2 => \N__10716\,
            in3 => \N__10748\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10131\,
            in3 => \N__10525\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10773\,
            in1 => \N__10747\,
            in2 => \N__10715\,
            in3 => \N__10161\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10155\,
            in1 => \N__10143\,
            in2 => \N__10130\,
            in3 => \N__10109\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__10431\,
            in1 => \N__10098\,
            in2 => \N__10086\,
            in3 => \N__10455\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__10705\,
            in1 => \N__10745\,
            in2 => \N__10554\,
            in3 => \N__10526\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__10551\,
            in1 => \N__10539\,
            in2 => \_gnd_net_\,
            in3 => \N__10524\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__10500\,
            in1 => \N__10488\,
            in2 => \N__10479\,
            in3 => \N__10476\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10778\,
            in1 => \N__10701\,
            in2 => \N__10464\,
            in3 => \N__10461\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10656\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10740\,
            in1 => \N__10776\,
            in2 => \N__10714\,
            in3 => \N__10443\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10656\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10777\,
            in1 => \N__10741\,
            in2 => \N__10713\,
            in3 => \N__10437\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10656\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10386\,
            in1 => \N__10419\,
            in2 => \N__10671\,
            in3 => \N__10407\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10775\,
            in1 => \N__10739\,
            in2 => \N__10395\,
            in3 => \N__10392\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10656\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__10785\,
            in1 => \N__10779\,
            in2 => \N__10749\,
            in3 => \N__10700\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10656\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

module U110_INTERRUPT (

    output INT2n

);

//JUST HOLD INT2 HIGH FOR NOW.

assign INT2n = 1;

endmodule

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 15 2025 11:38:09

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    TM : in std_logic_vector(1 downto 0);
    TT : in std_logic_vector(1 downto 0);
    D : inout std_logic_vector(7 downto 4);
    A : in std_logic_vector(31 downto 1);
    PIO_S0 : out std_logic;
    PORTSIZE : out std_logic;
    TICK60 : out std_logic;
    CIACS0n : out std_logic;
    CPUCONFn : in std_logic;
    CLK6 : in std_logic;
    CLK_CIA : out std_logic;
    BUFENn : out std_logic;
    AUTOBOOT : in std_logic;
    RnW : in std_logic;
    PIO_P2 : out std_logic;
    CIACS1n : out std_logic;
    BRIDGE_ENn : out std_logic;
    PIO_S1 : out std_logic;
    PIO_P0 : out std_logic;
    TICK50 : out std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : out std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    REGSPACEn : out std_logic;
    TSn : in std_logic;
    RTC_ENn : out std_logic;
    PIO_S2 : out std_logic;
    ATA_ENn : out std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    CONFIGENn : out std_logic;
    TACKn : inout std_logic;
    ROMENn : out std_logic;
    PIO_P1 : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__11575\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4115\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_14\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \U409_AUTOCONFIG.N_213_2_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_249_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_250_1\ : std_logic;
signal \U409_AUTOCONFIG.N_249\ : std_logic;
signal \U409_AUTOCONFIG.N_250_1_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.N_167_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_233\ : std_logic;
signal \U409_AUTOCONFIG.N_231_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_a5_0_0\ : std_logic;
signal \U409_AUTOCONFIG.N_212\ : std_logic;
signal \U409_AUTOCONFIG.N_213_2\ : std_logic;
signal \U409_AUTOCONFIG.N_212_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_3_0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_165\ : std_logic;
signal \U409_AUTOCONFIG.un1_A_16Z0Z_2\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_0\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U409_ADDRESS_DECODE.REG_SPACEZ0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_0_0\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_1_0\ : std_logic;
signal \U409_AUTOCONFIG.N_168_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_167\ : std_logic;
signal \U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0\ : std_logic;
signal \U409_AUTOCONFIG.N_166\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\ : std_logic;
signal \U409_AUTOCONFIG.N_173\ : std_logic;
signal \U409_AUTOCONFIG.N_249_1_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_155_0\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U409_AUTOCONFIG.un1_A_19Z0Z_1_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn_i\ : std_logic;
signal \U409_ADDRESS_DECODE.un2_REGSPACEn_0_0\ : std_logic;
signal \U409_ADDRESS_DECODE.REG_SPACEZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U409_AUTOCONFIG.un1_A_11Z0Z_0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.un1_AZ0Z_11\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U409_AUTOCONFIG.N_174\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.REG_SPACE_3\ : std_logic;
signal \A_c_25\ : std_logic;
signal \U409_ADDRESS_DECODE.REG_SPACE_3_cascade_\ : std_logic;
signal \A_c_24\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_26\ : std_logic;
signal \D_1_i\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG_D_OUT_0_i_3\ : std_logic;
signal \AUTOCONFIG_SPACE_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0_a3_0\ : std_logic;
signal \CPUCONFn_c\ : std_logic;
signal \U409_AUTOCONFIG.AC_STARTZ0\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\ : std_logic;
signal \U409_AUTOCONFIG_D_OUT_0_i_0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNO_0Z0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.N_265_0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNO_0Z0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_8_0_0\ : std_logic;
signal \U409_AUTOCONFIG.STATE4\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_8Z0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.N_248_0\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_8Z0Z_0_cascade_\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RTC_ENn_i\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACE_3\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACE_2_0\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOVECTOR_8\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOVECTOR_10_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOVECTOR_9\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG_D_OUT_0_i_1\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2\ : std_logic;
signal \U409_AUTOCONFIG_D_OUT_0_i_2\ : std_logic;
signal \INVU409_AUTOCONFIG.STATE_1C_net\ : std_logic;
signal \U409_AUTOCONFIG.STATE_d_2_cascade_\ : std_logic;
signal \A_c_31\ : std_logic;
signal \A_c_30\ : std_logic;
signal \BRIDGE_BASE_3\ : std_logic;
signal \A_c_29\ : std_logic;
signal \A_c_28\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2Z0Z_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5\ : std_logic;
signal \CONFIGENn_c\ : std_logic;
signal \INVU409_AUTOCONFIG.AC_TACKC_net\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U409_AUTOCONFIG.ATA_BASE11Z0Z_1\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U409_AUTOCONFIG.STATEZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.ATA_BASE11_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.STATEZ0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_6\ : std_logic;
signal \ATA_BASE_6\ : std_logic;
signal \D_in_6\ : std_logic;
signal \BRIDGE_BASE_2\ : std_logic;
signal \A_c_20\ : std_logic;
signal \ATA_BASE_4\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONF_RNIDFPAZ0Z3\ : std_logic;
signal \ATA_BASE_5\ : std_logic;
signal \INVU409_AUTOCONFIG.ATA_BASE_6C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_11_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_5_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_2\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\ : std_logic;
signal \U409_AUTOCONFIG.STATE_d_2\ : std_logic;
signal \U409_AUTOCONFIG.un1_AZ0Z_16\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONFZ0\ : std_logic;
signal \D_in_4\ : std_logic;
signal \BRIDGE_BASE_0\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\ : std_logic;
signal \BRIDGE_BASE_1\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_CONFC_net\ : std_logic;
signal \A_c_19\ : std_logic;
signal \A_c_18\ : std_logic;
signal \ATA_BASE_2\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2_cascade_\ : std_logic;
signal \ATA_BASE_7\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_5_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_6_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U409_ADDRESS_DECODE.un2_ATA_SPACEZ0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RTC_ENn\ : std_logic;
signal \U409_ADDRESS_DECODE_PORTSIZE_0_cascade_\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.un1_AUTOVECTOR_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_17_mux_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_3_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_3_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_6_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_17_mux\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1Z0Z_0\ : std_logic;
signal \A_c_22\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U409_TRANSFER_ACK.N_43\ : std_logic;
signal \ROMENn_c\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROMENnC_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \AC_TACK\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER5_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_1_out\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_OUTnC_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\ : std_logic;
signal \TM_c_0\ : std_logic;
signal \TM_c_1\ : std_logic;
signal \CONFIGURED\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_1\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_2\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i\ : std_logic;
signal \RnW_c\ : std_logic;
signal \D_in_5\ : std_logic;
signal \un1_AUTOCONFIG_SPACE_cascade_\ : std_logic;
signal \ATA_BASE_1\ : std_logic;
signal \U409_AUTOCONFIG.STATE_RNIS3FU2Z0Z_0\ : std_logic;
signal \un1_AUTOCONFIG_SPACE\ : std_logic;
signal \D_in_7\ : std_logic;
signal \ATA_BASE_3\ : std_logic;
signal \INVU409_AUTOCONFIG.ATA_BASE_1C_net\ : std_logic;
signal \CLK40_IN_c_g\ : std_logic;
signal \GB_BUFFER_CLK40_IN_c_g_THRU_CO\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\ : std_logic;
signal \U409_TRANSFER_ACK.N_28\ : std_logic;
signal \U409_TRANSFER_ACK.N_22\ : std_logic;
signal \U409_ADDRESS_DECODE_ROMEN_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_33_1\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_33\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_34\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.N_45\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_ENC_net\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_REGSPACEnZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0\ : std_logic;
signal \A_c_21\ : std_logic;
signal \OVL_c\ : std_logic;
signal \AGNUS_SPACE_0_cascade_\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4\ : std_logic;
signal \BUFENn_c\ : std_logic;
signal \U409_ADDRESS_DECODE_PORTSIZE_0\ : std_logic;
signal \AGNUS_SPACE_0\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \TCIn_1_i\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \bfn_13_6_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_ENZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_ATA_ENn_i\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_\ : std_logic;
signal \CIA_SPACE\ : std_logic;
signal \U409_CIA.VMA_RNOZ0Z_0_cascade_\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.TICK503_8\ : std_logic;
signal \U409_TICK.TICK503_11_cascade_\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.TICK603_11\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.TICK603_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \bfn_15_4_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_5\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_6\ : std_logic;
signal \U409_CIA.CLK_CIA_r_1_0\ : std_logic;
signal \U409_CIA.CLK_CIA6_3_cascade_\ : std_logic;
signal \CLK_CIA_c\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_7\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_6\ : std_logic;
signal \U409_CIA.CLK_CIA6_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_0\ : std_logic;
signal \U409_CIA.CLK_CIA6_4_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \bfn_15_6_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \bfn_15_7_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS1n_i\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \CIA_ENABLE\ : std_logic;
signal \A_c_12\ : std_logic;
signal \CIA_ENABLE_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS0n_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \PIO_P1_wire\ : std_logic;
signal \CPUCONFn_wire\ : std_logic;
signal \RTC_ENn_wire\ : std_logic;
signal \TM_wire\ : std_logic_vector(1 downto 0);
signal \RAMSPACEn_wire\ : std_logic;
signal \ROMENn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \PIO_P2_wire\ : std_logic;
signal \BRIDGE_ENn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CIACS0n_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CONFIGENn_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \PIO_P0_wire\ : std_logic;
signal \ATA_ENn_wire\ : std_logic;
signal \CIACS1n_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \CLK_CIA_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \PIO_S0_wire\ : std_logic;
signal \PIO_S2_wire\ : std_logic;
signal \PIO_S1_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    \CLK40_IN_wire\ <= CLK40_IN;
    \A_wire\ <= A;
    \TT_wire\ <= TT;
    PIO_P1 <= \PIO_P1_wire\;
    \CPUCONFn_wire\ <= CPUCONFn;
    RTC_ENn <= \RTC_ENn_wire\;
    \TM_wire\ <= TM;
    RAMSPACEn <= \RAMSPACEn_wire\;
    ROMENn <= \ROMENn_wire\;
    TBIn <= \TBIn_wire\;
    \TSn_wire\ <= TSn;
    PORTSIZE <= \PORTSIZE_wire\;
    PIO_P2 <= \PIO_P2_wire\;
    BRIDGE_ENn <= \BRIDGE_ENn_wire\;
    \RESETn_wire\ <= RESETn;
    CIACS0n <= \CIACS0n_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TCIn <= \TCIn_wire\;
    \RnW_wire\ <= RnW;
    CONFIGENn <= \CONFIGENn_wire\;
    TICK60 <= \TICK60_wire\;
    PIO_P0 <= \PIO_P0_wire\;
    ATA_ENn <= \ATA_ENn_wire\;
    CIACS1n <= \CIACS1n_wire\;
    REGSPACEn <= \REGSPACEn_wire\;
    CLK_CIA <= \CLK_CIA_wire\;
    BUFENn <= \BUFENn_wire\;
    PIO_S0 <= \PIO_S0_wire\;
    PIO_S2 <= \PIO_S2_wire\;
    PIO_S1 <= \PIO_S1_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__7904\,
            RESETB => \N__10466\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11573\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11575\,
            DIN => \N__11574\,
            DOUT => \N__11573\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11575\,
            PADOUT => \N__11574\,
            PADIN => \N__11573\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11563\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11565\,
            DIN => \N__11564\,
            DOUT => \N__11563\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11565\,
            PADOUT => \N__11564\,
            PADIN => \N__11563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11553\,
            GLOBALBUFFEROUTPUT => \CLK40_IN_c_g\
        );

    \CLK40_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11555\,
            DIN => \N__11554\,
            DOUT => \N__11553\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11555\,
            PADOUT => \N__11554\,
            PADIN => \N__11553\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11544\,
            DIN => \N__11543\,
            DOUT => \N__11542\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11544\,
            PADOUT => \N__11543\,
            PADIN => \N__11542\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11535\,
            DIN => \N__11534\,
            DOUT => \N__11533\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11535\,
            PADOUT => \N__11534\,
            PADIN => \N__11533\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_P1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11526\,
            DIN => \N__11525\,
            DOUT => \N__11524\,
            PACKAGEPIN => \PIO_P1_wire\
        );

    \PIO_P1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11526\,
            PADOUT => \N__11525\,
            PADIN => \N__11524\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10433\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11517\,
            DIN => \N__11516\,
            DOUT => \N__11515\,
            PACKAGEPIN => D(7)
        );

    \D_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11517\,
            PADOUT => \N__11516\,
            PADIN => \N__11515\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5178\,
            DIN0 => \D_in_7\,
            DOUT0 => \N__5114\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11508\,
            DIN => \N__11507\,
            DOUT => \N__11506\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11508\,
            PADOUT => \N__11507\,
            PADIN => \N__11506\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUCONFn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11499\,
            DIN => \N__11498\,
            DOUT => \N__11497\,
            PACKAGEPIN => \CPUCONFn_wire\
        );

    \CPUCONFn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11499\,
            PADOUT => \N__11498\,
            PADIN => \N__11497\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CPUCONFn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RTC_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11490\,
            DIN => \N__11489\,
            DOUT => \N__11488\,
            PACKAGEPIN => \RTC_ENn_wire\
        );

    \RTC_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11490\,
            PADOUT => \N__11489\,
            PADIN => \N__11488\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5237\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11481\,
            DIN => \N__11480\,
            DOUT => \N__11479\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11481\,
            PADOUT => \N__11480\,
            PADIN => \N__11479\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11472\,
            DIN => \N__11471\,
            DOUT => \N__11470\,
            PACKAGEPIN => D(4)
        );

    \D_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11472\,
            PADOUT => \N__11471\,
            PADIN => \N__11470\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5160\,
            DIN0 => \D_in_4\,
            DOUT0 => \N__5036\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11463\,
            DIN => \N__11462\,
            DOUT => \N__11461\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11463\,
            PADOUT => \N__11462\,
            PADIN => \N__11461\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11454\,
            DIN => \N__11453\,
            DOUT => \N__11452\,
            PACKAGEPIN => \TM_wire\(1)
        );

    \TM_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11454\,
            PADOUT => \N__11453\,
            PADIN => \N__11452\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11445\,
            DIN => \N__11444\,
            DOUT => \N__11443\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11445\,
            PADOUT => \N__11444\,
            PADIN => \N__11443\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11436\,
            DIN => \N__11435\,
            DOUT => \N__11434\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11436\,
            PADOUT => \N__11435\,
            PADIN => \N__11434\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8879\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11427\,
            DIN => \N__11426\,
            DOUT => \N__11425\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11427\,
            PADOUT => \N__11426\,
            PADIN => \N__11425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11418\,
            DIN => \N__11417\,
            DOUT => \N__11416\,
            PACKAGEPIN => \ROMENn_wire\
        );

    \ROMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11418\,
            PADOUT => \N__11417\,
            PADIN => \N__11416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7304\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11409\,
            DIN => \N__11408\,
            DOUT => \N__11407\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11409\,
            PADOUT => \N__11408\,
            PADIN => \N__11407\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8969\,
            DIN0 => OPEN,
            DOUT0 => \N__7756\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11400\,
            DIN => \N__11399\,
            DOUT => \N__11398\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11400\,
            PADOUT => \N__11399\,
            PADIN => \N__11398\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11391\,
            DIN => \N__11390\,
            DOUT => \N__11389\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11391\,
            PADOUT => \N__11390\,
            PADIN => \N__11389\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6860\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_P2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11382\,
            DIN => \N__11381\,
            DOUT => \N__11380\,
            PACKAGEPIN => \PIO_P2_wire\
        );

    \PIO_P2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11382\,
            PADOUT => \N__11381\,
            PADIN => \N__11380\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4175\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11373\,
            DIN => \N__11372\,
            DOUT => \N__11371\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11373\,
            PADOUT => \N__11372\,
            PADIN => \N__11371\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BRIDGE_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11364\,
            DIN => \N__11363\,
            DOUT => \N__11362\,
            PACKAGEPIN => \BRIDGE_ENn_wire\
        );

    \BRIDGE_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11364\,
            PADOUT => \N__11363\,
            PADIN => \N__11362\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8276\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11355\,
            DIN => \N__11354\,
            DOUT => \N__11353\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11355\,
            PADOUT => \N__11354\,
            PADIN => \N__11353\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11346\,
            DIN => \N__11345\,
            DOUT => \N__11344\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11346\,
            PADOUT => \N__11345\,
            PADIN => \N__11344\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11337\,
            DIN => \N__11336\,
            DOUT => \N__11335\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11337\,
            PADOUT => \N__11336\,
            PADIN => \N__11335\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11328\,
            DIN => \N__11327\,
            DOUT => \N__11326\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11328\,
            PADOUT => \N__11327\,
            PADIN => \N__11326\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11319\,
            DIN => \N__11318\,
            DOUT => \N__11317\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11319\,
            PADOUT => \N__11318\,
            PADIN => \N__11317\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11310\,
            DIN => \N__11309\,
            DOUT => \N__11308\,
            PACKAGEPIN => \CIACS0n_wire\
        );

    \CIACS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11310\,
            PADOUT => \N__11309\,
            PADIN => \N__11308\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10685\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11301\,
            DIN => \N__11300\,
            DOUT => \N__11299\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11301\,
            PADOUT => \N__11300\,
            PADIN => \N__11299\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7859\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11292\,
            DIN => \N__11291\,
            DOUT => \N__11290\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11292\,
            PADOUT => \N__11291\,
            PADIN => \N__11290\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11283\,
            DIN => \N__11282\,
            DOUT => \N__11281\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11283\,
            PADOUT => \N__11282\,
            PADIN => \N__11281\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11274\,
            DIN => \N__11273\,
            DOUT => \N__11272\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11274\,
            PADOUT => \N__11273\,
            PADIN => \N__11272\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11265\,
            DIN => \N__11264\,
            DOUT => \N__11263\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11265\,
            PADOUT => \N__11264\,
            PADIN => \N__11263\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11256\,
            DIN => \N__11255\,
            DOUT => \N__11254\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11256\,
            PADOUT => \N__11255\,
            PADIN => \N__11254\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8921\,
            DIN0 => OPEN,
            DOUT0 => \N__7757\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11247\,
            DIN => \N__11246\,
            DOUT => \N__11245\,
            PACKAGEPIN => D(5)
        );

    \D_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11247\,
            PADOUT => \N__11246\,
            PADIN => \N__11245\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5179\,
            DIN0 => \D_in_5\,
            DOUT0 => \N__5369\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11238\,
            DIN => \N__11237\,
            DOUT => \N__11236\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11238\,
            PADOUT => \N__11237\,
            PADIN => \N__11236\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11229\,
            DIN => \N__11228\,
            DOUT => \N__11227\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11229\,
            PADOUT => \N__11228\,
            PADIN => \N__11227\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11220\,
            DIN => \N__11219\,
            DOUT => \N__11218\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11220\,
            PADOUT => \N__11219\,
            PADIN => \N__11218\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CONFIGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11211\,
            DIN => \N__11210\,
            DOUT => \N__11209\,
            PACKAGEPIN => \CONFIGENn_wire\
        );

    \CONFIGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11211\,
            PADOUT => \N__11210\,
            PADIN => \N__11209\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5681\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11202\,
            DIN => \N__11201\,
            DOUT => \N__11200\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11202\,
            PADOUT => \N__11201\,
            PADIN => \N__11200\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9365\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11193\,
            DIN => \N__11192\,
            DOUT => \N__11191\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11193\,
            PADOUT => \N__11192\,
            PADIN => \N__11191\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_P0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11184\,
            DIN => \N__11183\,
            DOUT => \N__11182\,
            PACKAGEPIN => \PIO_P0_wire\
        );

    \PIO_P0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11184\,
            PADOUT => \N__11183\,
            PADIN => \N__11182\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10730\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11175\,
            DIN => \N__11174\,
            DOUT => \N__11173\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11175\,
            PADOUT => \N__11174\,
            PADIN => \N__11173\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11166\,
            DIN => \N__11165\,
            DOUT => \N__11164\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11166\,
            PADOUT => \N__11165\,
            PADIN => \N__11164\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ATA_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11157\,
            DIN => \N__11156\,
            DOUT => \N__11155\,
            PACKAGEPIN => \ATA_ENn_wire\
        );

    \ATA_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11157\,
            PADOUT => \N__11156\,
            PADIN => \N__11155\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9197\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11148\,
            DIN => \N__11147\,
            DOUT => \N__11146\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11148\,
            PADOUT => \N__11147\,
            PADIN => \N__11146\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11139\,
            DIN => \N__11138\,
            DOUT => \N__11137\,
            PACKAGEPIN => \CIACS1n_wire\
        );

    \CIACS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11139\,
            PADOUT => \N__11138\,
            PADIN => \N__11137\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10397\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11130\,
            DIN => \N__11129\,
            DOUT => \N__11128\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11130\,
            PADOUT => \N__11129\,
            PADIN => \N__11128\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4460\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11121\,
            DIN => \N__11120\,
            DOUT => \N__11119\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11121\,
            PADOUT => \N__11120\,
            PADIN => \N__11119\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_CIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11112\,
            DIN => \N__11111\,
            DOUT => \N__11110\,
            PACKAGEPIN => \CLK_CIA_wire\
        );

    \CLK_CIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11112\,
            PADOUT => \N__11111\,
            PADIN => \N__11110\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10193\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11103\,
            DIN => \N__11102\,
            DOUT => \N__11101\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11103\,
            PADOUT => \N__11102\,
            PADIN => \N__11101\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11094\,
            DIN => \N__11093\,
            DOUT => \N__11092\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11094\,
            PADOUT => \N__11093\,
            PADIN => \N__11092\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8959\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__7749\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11085\,
            DIN => \N__11084\,
            DOUT => \N__11083\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11085\,
            PADOUT => \N__11084\,
            PADIN => \N__11083\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11076\,
            DIN => \N__11075\,
            DOUT => \N__11074\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11076\,
            PADOUT => \N__11075\,
            PADIN => \N__11074\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9011\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_S0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11067\,
            DIN => \N__11066\,
            DOUT => \N__11065\,
            PACKAGEPIN => \PIO_S0_wire\
        );

    \PIO_S0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11067\,
            PADOUT => \N__11066\,
            PADIN => \N__11065\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4199\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11058\,
            DIN => \N__11057\,
            DOUT => \N__11056\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11058\,
            PADOUT => \N__11057\,
            PADIN => \N__11056\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_S2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11049\,
            DIN => \N__11048\,
            DOUT => \N__11047\,
            PACKAGEPIN => \PIO_S2_wire\
        );

    \PIO_S2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11049\,
            PADOUT => \N__11048\,
            PADIN => \N__11047\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10462\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11040\,
            DIN => \N__11039\,
            DOUT => \N__11038\,
            PACKAGEPIN => D(6)
        );

    \D_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11040\,
            PADOUT => \N__11039\,
            PADIN => \N__11038\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5180\,
            DIN0 => \D_in_6\,
            DOUT0 => \N__5330\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11031\,
            DIN => \N__11030\,
            DOUT => \N__11029\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11031\,
            PADOUT => \N__11030\,
            PADIN => \N__11029\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11022\,
            DIN => \N__11021\,
            DOUT => \N__11020\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11022\,
            PADOUT => \N__11021\,
            PADIN => \N__11020\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_S1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11013\,
            DIN => \N__11012\,
            DOUT => \N__11011\,
            PACKAGEPIN => \PIO_S1_wire\
        );

    \PIO_S1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11013\,
            PADOUT => \N__11012\,
            PADIN => \N__11011\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4316\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11004\,
            DIN => \N__11003\,
            DOUT => \N__11002\,
            PACKAGEPIN => \TM_wire\(0)
        );

    \TM_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11004\,
            PADOUT => \N__11003\,
            PADIN => \N__11002\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10995\,
            DIN => \N__10994\,
            DOUT => \N__10993\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10995\,
            PADOUT => \N__10994\,
            PADIN => \N__10993\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10986\,
            DIN => \N__10985\,
            DOUT => \N__10984\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10986\,
            PADOUT => \N__10985\,
            PADIN => \N__10984\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2644\ : InMux
    port map (
            O => \N__10967\,
            I => \N__10964\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__10964\,
            I => \N__10960\
        );

    \I__2642\ : InMux
    port map (
            O => \N__10963\,
            I => \N__10957\
        );

    \I__2641\ : Span4Mux_v
    port map (
            O => \N__10960\,
            I => \N__10954\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__10957\,
            I => \N__10951\
        );

    \I__2639\ : Sp12to4
    port map (
            O => \N__10954\,
            I => \N__10947\
        );

    \I__2638\ : Span4Mux_v
    port map (
            O => \N__10951\,
            I => \N__10944\
        );

    \I__2637\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10941\
        );

    \I__2636\ : Odrv12
    port map (
            O => \N__10947\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2635\ : Odrv4
    port map (
            O => \N__10944\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__10941\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__10934\,
            I => \N__10930\
        );

    \I__2632\ : InMux
    port map (
            O => \N__10933\,
            I => \N__10926\
        );

    \I__2631\ : InMux
    port map (
            O => \N__10930\,
            I => \N__10923\
        );

    \I__2630\ : CascadeMux
    port map (
            O => \N__10929\,
            I => \N__10920\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__10926\,
            I => \N__10908\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__10923\,
            I => \N__10908\
        );

    \I__2627\ : InMux
    port map (
            O => \N__10920\,
            I => \N__10905\
        );

    \I__2626\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10900\
        );

    \I__2625\ : InMux
    port map (
            O => \N__10918\,
            I => \N__10900\
        );

    \I__2624\ : InMux
    port map (
            O => \N__10917\,
            I => \N__10897\
        );

    \I__2623\ : CascadeMux
    port map (
            O => \N__10916\,
            I => \N__10894\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__10915\,
            I => \N__10890\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__10914\,
            I => \N__10885\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__10913\,
            I => \N__10881\
        );

    \I__2619\ : Span4Mux_v
    port map (
            O => \N__10908\,
            I => \N__10872\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__10905\,
            I => \N__10872\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__10900\,
            I => \N__10872\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__10897\,
            I => \N__10868\
        );

    \I__2615\ : InMux
    port map (
            O => \N__10894\,
            I => \N__10859\
        );

    \I__2614\ : InMux
    port map (
            O => \N__10893\,
            I => \N__10859\
        );

    \I__2613\ : InMux
    port map (
            O => \N__10890\,
            I => \N__10859\
        );

    \I__2612\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10859\
        );

    \I__2611\ : InMux
    port map (
            O => \N__10888\,
            I => \N__10856\
        );

    \I__2610\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10853\
        );

    \I__2609\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10850\
        );

    \I__2608\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10847\
        );

    \I__2607\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10842\
        );

    \I__2606\ : InMux
    port map (
            O => \N__10879\,
            I => \N__10842\
        );

    \I__2605\ : Span4Mux_v
    port map (
            O => \N__10872\,
            I => \N__10839\
        );

    \I__2604\ : InMux
    port map (
            O => \N__10871\,
            I => \N__10836\
        );

    \I__2603\ : Span4Mux_h
    port map (
            O => \N__10868\,
            I => \N__10827\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__10859\,
            I => \N__10827\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__10856\,
            I => \N__10827\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__10853\,
            I => \N__10827\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__10850\,
            I => \N__10818\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__10847\,
            I => \N__10818\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__10842\,
            I => \N__10818\
        );

    \I__2596\ : Span4Mux_h
    port map (
            O => \N__10839\,
            I => \N__10811\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__10836\,
            I => \N__10811\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__10827\,
            I => \N__10808\
        );

    \I__2593\ : InMux
    port map (
            O => \N__10826\,
            I => \N__10805\
        );

    \I__2592\ : InMux
    port map (
            O => \N__10825\,
            I => \N__10802\
        );

    \I__2591\ : Span4Mux_v
    port map (
            O => \N__10818\,
            I => \N__10799\
        );

    \I__2590\ : InMux
    port map (
            O => \N__10817\,
            I => \N__10794\
        );

    \I__2589\ : InMux
    port map (
            O => \N__10816\,
            I => \N__10794\
        );

    \I__2588\ : Span4Mux_v
    port map (
            O => \N__10811\,
            I => \N__10790\
        );

    \I__2587\ : Span4Mux_h
    port map (
            O => \N__10808\,
            I => \N__10787\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__10805\,
            I => \N__10782\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__10802\,
            I => \N__10782\
        );

    \I__2584\ : Span4Mux_v
    port map (
            O => \N__10799\,
            I => \N__10777\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__10794\,
            I => \N__10777\
        );

    \I__2582\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10774\
        );

    \I__2581\ : Sp12to4
    port map (
            O => \N__10790\,
            I => \N__10770\
        );

    \I__2580\ : Sp12to4
    port map (
            O => \N__10787\,
            I => \N__10761\
        );

    \I__2579\ : Span12Mux_v
    port map (
            O => \N__10782\,
            I => \N__10761\
        );

    \I__2578\ : Sp12to4
    port map (
            O => \N__10777\,
            I => \N__10761\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__10774\,
            I => \N__10761\
        );

    \I__2576\ : InMux
    port map (
            O => \N__10773\,
            I => \N__10758\
        );

    \I__2575\ : Span12Mux_h
    port map (
            O => \N__10770\,
            I => \N__10755\
        );

    \I__2574\ : Span12Mux_v
    port map (
            O => \N__10761\,
            I => \N__10752\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__10758\,
            I => \N__10749\
        );

    \I__2572\ : Span12Mux_v
    port map (
            O => \N__10755\,
            I => \N__10746\
        );

    \I__2571\ : Span12Mux_h
    port map (
            O => \N__10752\,
            I => \N__10741\
        );

    \I__2570\ : Span12Mux_v
    port map (
            O => \N__10749\,
            I => \N__10741\
        );

    \I__2569\ : Odrv12
    port map (
            O => \N__10746\,
            I => \RESETn_c\
        );

    \I__2568\ : Odrv12
    port map (
            O => \N__10741\,
            I => \RESETn_c\
        );

    \I__2567\ : InMux
    port map (
            O => \N__10736\,
            I => \N__10733\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__10733\,
            I => \CIA_ENABLE\
        );

    \I__2565\ : IoInMux
    port map (
            O => \N__10730\,
            I => \N__10727\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__10727\,
            I => \N__10724\
        );

    \I__2563\ : Span4Mux_s0_h
    port map (
            O => \N__10724\,
            I => \N__10720\
        );

    \I__2562\ : InMux
    port map (
            O => \N__10723\,
            I => \N__10717\
        );

    \I__2561\ : Sp12to4
    port map (
            O => \N__10720\,
            I => \N__10714\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__10717\,
            I => \N__10711\
        );

    \I__2559\ : Span12Mux_s10_v
    port map (
            O => \N__10714\,
            I => \N__10708\
        );

    \I__2558\ : Span12Mux_s10_v
    port map (
            O => \N__10711\,
            I => \N__10705\
        );

    \I__2557\ : Span12Mux_h
    port map (
            O => \N__10708\,
            I => \N__10702\
        );

    \I__2556\ : Span12Mux_h
    port map (
            O => \N__10705\,
            I => \N__10699\
        );

    \I__2555\ : Span12Mux_h
    port map (
            O => \N__10702\,
            I => \N__10696\
        );

    \I__2554\ : Span12Mux_h
    port map (
            O => \N__10699\,
            I => \N__10693\
        );

    \I__2553\ : Odrv12
    port map (
            O => \N__10696\,
            I => \A_c_12\
        );

    \I__2552\ : Odrv12
    port map (
            O => \N__10693\,
            I => \A_c_12\
        );

    \I__2551\ : CascadeMux
    port map (
            O => \N__10688\,
            I => \CIA_ENABLE_cascade_\
        );

    \I__2550\ : IoInMux
    port map (
            O => \N__10685\,
            I => \N__10682\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__10682\,
            I => \N__10679\
        );

    \I__2548\ : Span4Mux_s3_h
    port map (
            O => \N__10679\,
            I => \N__10676\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__10676\,
            I => \N__10673\
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__10673\,
            I => \U409_ADDRESS_DECODE_un1_CIACS0n_i\
        );

    \I__2545\ : InMux
    port map (
            O => \N__10670\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__2544\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10663\
        );

    \I__2543\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10660\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__10663\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__10660\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2540\ : InMux
    port map (
            O => \N__10655\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__2539\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10648\
        );

    \I__2538\ : InMux
    port map (
            O => \N__10651\,
            I => \N__10645\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__10648\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10645\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2535\ : InMux
    port map (
            O => \N__10640\,
            I => \N__10637\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__10637\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__2533\ : InMux
    port map (
            O => \N__10634\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__2532\ : InMux
    port map (
            O => \N__10631\,
            I => \N__10627\
        );

    \I__2531\ : InMux
    port map (
            O => \N__10630\,
            I => \N__10624\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__10627\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__10624\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__2528\ : InMux
    port map (
            O => \N__10619\,
            I => \N__10616\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__10616\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__2526\ : InMux
    port map (
            O => \N__10613\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__2525\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10606\
        );

    \I__2524\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10603\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__10606\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__10603\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__10598\,
            I => \N__10595\
        );

    \I__2520\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10592\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__10592\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__2518\ : InMux
    port map (
            O => \N__10589\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__2517\ : InMux
    port map (
            O => \N__10586\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__2516\ : InMux
    port map (
            O => \N__10583\,
            I => \N__10579\
        );

    \I__2515\ : InMux
    port map (
            O => \N__10582\,
            I => \N__10576\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__10579\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__10576\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__2512\ : ClkMux
    port map (
            O => \N__10571\,
            I => \N__10544\
        );

    \I__2511\ : ClkMux
    port map (
            O => \N__10570\,
            I => \N__10544\
        );

    \I__2510\ : ClkMux
    port map (
            O => \N__10569\,
            I => \N__10544\
        );

    \I__2509\ : ClkMux
    port map (
            O => \N__10568\,
            I => \N__10544\
        );

    \I__2508\ : ClkMux
    port map (
            O => \N__10567\,
            I => \N__10544\
        );

    \I__2507\ : ClkMux
    port map (
            O => \N__10566\,
            I => \N__10544\
        );

    \I__2506\ : ClkMux
    port map (
            O => \N__10565\,
            I => \N__10544\
        );

    \I__2505\ : ClkMux
    port map (
            O => \N__10564\,
            I => \N__10544\
        );

    \I__2504\ : ClkMux
    port map (
            O => \N__10563\,
            I => \N__10544\
        );

    \I__2503\ : GlobalMux
    port map (
            O => \N__10544\,
            I => \N__10541\
        );

    \I__2502\ : gio2CtrlBuf
    port map (
            O => \N__10541\,
            I => \CLK6_c_g\
        );

    \I__2501\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10532\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10537\,
            I => \N__10529\
        );

    \I__2499\ : InMux
    port map (
            O => \N__10536\,
            I => \N__10526\
        );

    \I__2498\ : InMux
    port map (
            O => \N__10535\,
            I => \N__10523\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__10532\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__10529\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__10526\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__10523\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__10514\,
            I => \N__10511\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10511\,
            I => \N__10506\
        );

    \I__2491\ : InMux
    port map (
            O => \N__10510\,
            I => \N__10498\
        );

    \I__2490\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10498\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__10506\,
            I => \N__10495\
        );

    \I__2488\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10492\
        );

    \I__2487\ : InMux
    port map (
            O => \N__10504\,
            I => \N__10487\
        );

    \I__2486\ : InMux
    port map (
            O => \N__10503\,
            I => \N__10487\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__10498\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__10495\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__10492\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__10487\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2481\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10474\
        );

    \I__2480\ : InMux
    port map (
            O => \N__10477\,
            I => \N__10471\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__10474\,
            I => \U409_CIA.CIA_CLK_COUNT11_2\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__10471\,
            I => \U409_CIA.CIA_CLK_COUNT11_2\
        );

    \I__2477\ : IoInMux
    port map (
            O => \N__10466\,
            I => \N__10463\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__10463\,
            I => \N__10459\
        );

    \I__2475\ : IoInMux
    port map (
            O => \N__10462\,
            I => \N__10456\
        );

    \I__2474\ : Span4Mux_s0_v
    port map (
            O => \N__10459\,
            I => \N__10453\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__10456\,
            I => \N__10450\
        );

    \I__2472\ : Sp12to4
    port map (
            O => \N__10453\,
            I => \N__10447\
        );

    \I__2471\ : Span4Mux_s3_h
    port map (
            O => \N__10450\,
            I => \N__10444\
        );

    \I__2470\ : Span12Mux_h
    port map (
            O => \N__10447\,
            I => \N__10441\
        );

    \I__2469\ : Span4Mux_v
    port map (
            O => \N__10444\,
            I => \N__10438\
        );

    \I__2468\ : Odrv12
    port map (
            O => \N__10441\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__10438\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2466\ : IoInMux
    port map (
            O => \N__10433\,
            I => \N__10430\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__10430\,
            I => \N__10427\
        );

    \I__2464\ : IoSpan4Mux
    port map (
            O => \N__10427\,
            I => \N__10423\
        );

    \I__2463\ : InMux
    port map (
            O => \N__10426\,
            I => \N__10420\
        );

    \I__2462\ : IoSpan4Mux
    port map (
            O => \N__10423\,
            I => \N__10417\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__10420\,
            I => \N__10414\
        );

    \I__2460\ : Span4Mux_s3_h
    port map (
            O => \N__10417\,
            I => \N__10409\
        );

    \I__2459\ : Span4Mux_v
    port map (
            O => \N__10414\,
            I => \N__10409\
        );

    \I__2458\ : Sp12to4
    port map (
            O => \N__10409\,
            I => \N__10406\
        );

    \I__2457\ : Span12Mux_h
    port map (
            O => \N__10406\,
            I => \N__10403\
        );

    \I__2456\ : Span12Mux_h
    port map (
            O => \N__10403\,
            I => \N__10400\
        );

    \I__2455\ : Odrv12
    port map (
            O => \N__10400\,
            I => \A_c_13\
        );

    \I__2454\ : IoInMux
    port map (
            O => \N__10397\,
            I => \N__10394\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__10394\,
            I => \N__10391\
        );

    \I__2452\ : Span4Mux_s3_h
    port map (
            O => \N__10391\,
            I => \N__10388\
        );

    \I__2451\ : Span4Mux_v
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__10385\,
            I => \U409_ADDRESS_DECODE_un1_CIACS1n_i\
        );

    \I__2449\ : InMux
    port map (
            O => \N__10382\,
            I => \N__10378\
        );

    \I__2448\ : InMux
    port map (
            O => \N__10381\,
            I => \N__10375\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__10378\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__10375\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2445\ : InMux
    port map (
            O => \N__10370\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__10367\,
            I => \N__10364\
        );

    \I__2443\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10360\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10363\,
            I => \N__10357\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__10360\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__10357\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2439\ : InMux
    port map (
            O => \N__10352\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__2438\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10345\
        );

    \I__2437\ : InMux
    port map (
            O => \N__10348\,
            I => \N__10342\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__10345\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__10342\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10337\,
            I => \N__10334\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__10334\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__2432\ : InMux
    port map (
            O => \N__10331\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__2431\ : InMux
    port map (
            O => \N__10328\,
            I => \N__10324\
        );

    \I__2430\ : InMux
    port map (
            O => \N__10327\,
            I => \N__10321\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__10324\,
            I => \N__10318\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__10321\,
            I => \N__10315\
        );

    \I__2427\ : Odrv4
    port map (
            O => \N__10318\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2426\ : Odrv4
    port map (
            O => \N__10315\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2425\ : InMux
    port map (
            O => \N__10310\,
            I => \N__10307\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__10307\,
            I => \N__10304\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__10304\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10301\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__2421\ : InMux
    port map (
            O => \N__10298\,
            I => \N__10294\
        );

    \I__2420\ : InMux
    port map (
            O => \N__10297\,
            I => \N__10291\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__10294\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__10291\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10286\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10279\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10282\,
            I => \N__10276\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__10279\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__10276\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2412\ : InMux
    port map (
            O => \N__10271\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__10268\,
            I => \N__10265\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10265\,
            I => \N__10261\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10264\,
            I => \N__10258\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__10261\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__10258\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__10253\,
            I => \N__10250\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10250\,
            I => \N__10247\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10247\,
            I => \N__10244\
        );

    \I__2403\ : Odrv12
    port map (
            O => \N__10244\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__2402\ : InMux
    port map (
            O => \N__10241\,
            I => \bfn_15_7_0_\
        );

    \I__2401\ : InMux
    port map (
            O => \N__10238\,
            I => \N__10234\
        );

    \I__2400\ : InMux
    port map (
            O => \N__10237\,
            I => \N__10231\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__10234\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__10231\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2397\ : InMux
    port map (
            O => \N__10226\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10223\,
            I => \N__10220\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__10220\,
            I => \N__10216\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10219\,
            I => \N__10213\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__10216\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__10213\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10208\,
            I => \N__10205\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__10205\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__2389\ : InMux
    port map (
            O => \N__10202\,
            I => \N__10199\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__10199\,
            I => \U409_CIA.CLK_CIA_r_1_0\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__10196\,
            I => \U409_CIA.CLK_CIA6_3_cascade_\
        );

    \I__2386\ : IoInMux
    port map (
            O => \N__10193\,
            I => \N__10190\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__10190\,
            I => \N__10187\
        );

    \I__2384\ : IoSpan4Mux
    port map (
            O => \N__10187\,
            I => \N__10184\
        );

    \I__2383\ : Span4Mux_s3_v
    port map (
            O => \N__10184\,
            I => \N__10181\
        );

    \I__2382\ : Sp12to4
    port map (
            O => \N__10181\,
            I => \N__10176\
        );

    \I__2381\ : InMux
    port map (
            O => \N__10180\,
            I => \N__10173\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__10179\,
            I => \N__10169\
        );

    \I__2379\ : Span12Mux_s10_v
    port map (
            O => \N__10176\,
            I => \N__10166\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10173\,
            I => \N__10163\
        );

    \I__2377\ : InMux
    port map (
            O => \N__10172\,
            I => \N__10160\
        );

    \I__2376\ : InMux
    port map (
            O => \N__10169\,
            I => \N__10157\
        );

    \I__2375\ : Odrv12
    port map (
            O => \N__10166\,
            I => \CLK_CIA_c\
        );

    \I__2374\ : Odrv12
    port map (
            O => \N__10163\,
            I => \CLK_CIA_c\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__10160\,
            I => \CLK_CIA_c\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10157\,
            I => \CLK_CIA_c\
        );

    \I__2371\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10140\
        );

    \I__2370\ : InMux
    port map (
            O => \N__10147\,
            I => \N__10140\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10137\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10145\,
            I => \N__10134\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10140\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__10137\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__10134\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__10127\,
            I => \N__10119\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10126\,
            I => \N__10116\
        );

    \I__2362\ : InMux
    port map (
            O => \N__10125\,
            I => \N__10109\
        );

    \I__2361\ : InMux
    port map (
            O => \N__10124\,
            I => \N__10109\
        );

    \I__2360\ : InMux
    port map (
            O => \N__10123\,
            I => \N__10109\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10122\,
            I => \N__10104\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10119\,
            I => \N__10104\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__10116\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10109\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__10104\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__10097\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\
        );

    \I__2353\ : InMux
    port map (
            O => \N__10094\,
            I => \N__10091\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__10091\,
            I => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__10088\,
            I => \N__10083\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__10087\,
            I => \N__10079\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10086\,
            I => \N__10074\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10083\,
            I => \N__10074\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10071\
        );

    \I__2346\ : InMux
    port map (
            O => \N__10079\,
            I => \N__10068\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10074\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__10071\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__10068\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10061\,
            I => \N__10056\
        );

    \I__2341\ : InMux
    port map (
            O => \N__10060\,
            I => \N__10051\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10059\,
            I => \N__10051\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__10056\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__10051\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__2337\ : InMux
    port map (
            O => \N__10046\,
            I => \N__10041\
        );

    \I__2336\ : InMux
    port map (
            O => \N__10045\,
            I => \N__10038\
        );

    \I__2335\ : InMux
    port map (
            O => \N__10044\,
            I => \N__10035\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__10041\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__10038\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__10035\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10028\,
            I => \N__10024\
        );

    \I__2330\ : InMux
    port map (
            O => \N__10027\,
            I => \N__10021\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10024\,
            I => \U409_CIA.CLK_CIA6_4\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__10021\,
            I => \U409_CIA.CLK_CIA6_4\
        );

    \I__2327\ : InMux
    port map (
            O => \N__10016\,
            I => \N__10013\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__10013\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__10010\,
            I => \U409_CIA.CLK_CIA6_4_cascade_\
        );

    \I__2324\ : InMux
    port map (
            O => \N__10007\,
            I => \N__10004\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__10004\,
            I => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3\
        );

    \I__2322\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9993\
        );

    \I__2321\ : InMux
    port map (
            O => \N__10000\,
            I => \N__9993\
        );

    \I__2320\ : InMux
    port map (
            O => \N__9999\,
            I => \N__9990\
        );

    \I__2319\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9987\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__9993\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__9990\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__9987\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__2315\ : ClkMux
    port map (
            O => \N__9980\,
            I => \N__9971\
        );

    \I__2314\ : ClkMux
    port map (
            O => \N__9979\,
            I => \N__9971\
        );

    \I__2313\ : ClkMux
    port map (
            O => \N__9978\,
            I => \N__9971\
        );

    \I__2312\ : GlobalMux
    port map (
            O => \N__9971\,
            I => \N__9968\
        );

    \I__2311\ : gio2CtrlBuf
    port map (
            O => \N__9968\,
            I => \CLK28_IN_c_g\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__9965\,
            I => \N__9961\
        );

    \I__2309\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9955\
        );

    \I__2308\ : InMux
    port map (
            O => \N__9961\,
            I => \N__9955\
        );

    \I__2307\ : InMux
    port map (
            O => \N__9960\,
            I => \N__9952\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__9955\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__9952\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__9947\,
            I => \N__9941\
        );

    \I__2303\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9936\
        );

    \I__2302\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9936\
        );

    \I__2301\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9933\
        );

    \I__2300\ : InMux
    port map (
            O => \N__9941\,
            I => \N__9930\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__9936\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__9933\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__9930\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2296\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9919\
        );

    \I__2295\ : InMux
    port map (
            O => \N__9922\,
            I => \N__9916\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__9919\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__9916\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2292\ : InMux
    port map (
            O => \N__9911\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__2291\ : InMux
    port map (
            O => \N__9908\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__2290\ : InMux
    port map (
            O => \N__9905\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__2289\ : InMux
    port map (
            O => \N__9902\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__2288\ : InMux
    port map (
            O => \N__9899\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__2287\ : InMux
    port map (
            O => \N__9896\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\
        );

    \I__2286\ : InMux
    port map (
            O => \N__9893\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\
        );

    \I__2285\ : InMux
    port map (
            O => \N__9890\,
            I => \N__9887\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__9887\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__2283\ : InMux
    port map (
            O => \N__9884\,
            I => \N__9879\
        );

    \I__2282\ : InMux
    port map (
            O => \N__9883\,
            I => \N__9876\
        );

    \I__2281\ : InMux
    port map (
            O => \N__9882\,
            I => \N__9873\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__9879\,
            I => \N__9865\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__9876\,
            I => \N__9862\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__9873\,
            I => \N__9859\
        );

    \I__2277\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9854\
        );

    \I__2276\ : InMux
    port map (
            O => \N__9871\,
            I => \N__9854\
        );

    \I__2275\ : InMux
    port map (
            O => \N__9870\,
            I => \N__9847\
        );

    \I__2274\ : InMux
    port map (
            O => \N__9869\,
            I => \N__9847\
        );

    \I__2273\ : InMux
    port map (
            O => \N__9868\,
            I => \N__9847\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__9865\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__9862\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2270\ : Odrv4
    port map (
            O => \N__9859\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__9854\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__9847\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2267\ : InMux
    port map (
            O => \N__9836\,
            I => \N__9833\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__9833\,
            I => \N__9827\
        );

    \I__2265\ : InMux
    port map (
            O => \N__9832\,
            I => \N__9824\
        );

    \I__2264\ : InMux
    port map (
            O => \N__9831\,
            I => \N__9819\
        );

    \I__2263\ : InMux
    port map (
            O => \N__9830\,
            I => \N__9819\
        );

    \I__2262\ : Span4Mux_h
    port map (
            O => \N__9827\,
            I => \N__9811\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__9824\,
            I => \N__9806\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__9819\,
            I => \N__9806\
        );

    \I__2259\ : InMux
    port map (
            O => \N__9818\,
            I => \N__9803\
        );

    \I__2258\ : InMux
    port map (
            O => \N__9817\,
            I => \N__9800\
        );

    \I__2257\ : InMux
    port map (
            O => \N__9816\,
            I => \N__9793\
        );

    \I__2256\ : InMux
    port map (
            O => \N__9815\,
            I => \N__9793\
        );

    \I__2255\ : InMux
    port map (
            O => \N__9814\,
            I => \N__9793\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__9811\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2253\ : Odrv12
    port map (
            O => \N__9806\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__9803\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__9800\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__9793\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2249\ : CascadeMux
    port map (
            O => \N__9782\,
            I => \N__9778\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__9781\,
            I => \N__9772\
        );

    \I__2247\ : InMux
    port map (
            O => \N__9778\,
            I => \N__9769\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__9777\,
            I => \N__9766\
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__9776\,
            I => \N__9762\
        );

    \I__2244\ : CascadeMux
    port map (
            O => \N__9775\,
            I => \N__9757\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9772\,
            I => \N__9754\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__9769\,
            I => \N__9751\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9766\,
            I => \N__9748\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9765\,
            I => \N__9743\
        );

    \I__2239\ : InMux
    port map (
            O => \N__9762\,
            I => \N__9743\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9761\,
            I => \N__9736\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9760\,
            I => \N__9736\
        );

    \I__2236\ : InMux
    port map (
            O => \N__9757\,
            I => \N__9736\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__9754\,
            I => \N__9733\
        );

    \I__2234\ : Span4Mux_v
    port map (
            O => \N__9751\,
            I => \N__9728\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__9748\,
            I => \N__9728\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__9743\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9736\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__9733\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__9728\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2228\ : InMux
    port map (
            O => \N__9719\,
            I => \N__9715\
        );

    \I__2227\ : InMux
    port map (
            O => \N__9718\,
            I => \N__9712\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__9715\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__9712\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__9707\,
            I => \N__9703\
        );

    \I__2223\ : InMux
    port map (
            O => \N__9706\,
            I => \N__9700\
        );

    \I__2222\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9697\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__9700\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__9697\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__2219\ : CascadeMux
    port map (
            O => \N__9692\,
            I => \N__9689\
        );

    \I__2218\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9685\
        );

    \I__2217\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9682\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__9685\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__9682\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2214\ : InMux
    port map (
            O => \N__9677\,
            I => \N__9674\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__9674\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__9671\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__9668\,
            I => \N__9664\
        );

    \I__2210\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9661\
        );

    \I__2209\ : InMux
    port map (
            O => \N__9664\,
            I => \N__9658\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__9661\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__9658\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__2206\ : InMux
    port map (
            O => \N__9653\,
            I => \N__9650\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__9650\,
            I => \N__9646\
        );

    \I__2204\ : InMux
    port map (
            O => \N__9649\,
            I => \N__9643\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__9646\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__9643\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__9638\,
            I => \N__9633\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__9637\,
            I => \N__9630\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__9636\,
            I => \N__9626\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9633\,
            I => \N__9621\
        );

    \I__2197\ : InMux
    port map (
            O => \N__9630\,
            I => \N__9621\
        );

    \I__2196\ : InMux
    port map (
            O => \N__9629\,
            I => \N__9618\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9626\,
            I => \N__9615\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__9621\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__9618\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__9615\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9608\,
            I => \N__9604\
        );

    \I__2190\ : InMux
    port map (
            O => \N__9607\,
            I => \N__9601\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__9604\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__9601\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9596\,
            I => \N__9593\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9593\,
            I => \U409_TICK.TICK603_11\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9586\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9583\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__9586\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__9583\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__9578\,
            I => \U409_TICK.TICK603_8_cascade_\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9572\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9572\,
            I => \N__9568\
        );

    \I__2178\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9565\
        );

    \I__2177\ : Odrv4
    port map (
            O => \N__9568\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9565\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__9560\,
            I => \N__9557\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9557\,
            I => \N__9548\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9556\,
            I => \N__9539\
        );

    \I__2172\ : InMux
    port map (
            O => \N__9555\,
            I => \N__9539\
        );

    \I__2171\ : InMux
    port map (
            O => \N__9554\,
            I => \N__9539\
        );

    \I__2170\ : InMux
    port map (
            O => \N__9553\,
            I => \N__9539\
        );

    \I__2169\ : InMux
    port map (
            O => \N__9552\,
            I => \N__9534\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9551\,
            I => \N__9534\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9548\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__9539\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9534\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__9527\,
            I => \N__9519\
        );

    \I__2163\ : InMux
    port map (
            O => \N__9526\,
            I => \N__9508\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9525\,
            I => \N__9508\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9508\
        );

    \I__2160\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9508\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9499\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9519\,
            I => \N__9499\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9518\,
            I => \N__9499\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9517\,
            I => \N__9499\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9508\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9499\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__9494\,
            I => \N__9489\
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__9493\,
            I => \N__9486\
        );

    \I__2151\ : CascadeMux
    port map (
            O => \N__9492\,
            I => \N__9483\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9489\,
            I => \N__9470\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9470\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9470\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9470\
        );

    \I__2146\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9463\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9480\,
            I => \N__9463\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9479\,
            I => \N__9463\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9470\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9463\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__9458\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__9452\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9445\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9448\,
            I => \N__9442\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9445\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__9442\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2134\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9434\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__9434\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__2132\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__9428\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9421\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9424\,
            I => \N__9418\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__9421\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__9418\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9409\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9406\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9409\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__9406\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9401\,
            I => \N__9397\
        );

    \I__2121\ : InMux
    port map (
            O => \N__9400\,
            I => \N__9394\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9397\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__9394\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__2118\ : InMux
    port map (
            O => \N__9389\,
            I => \N__9386\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9386\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__9383\,
            I => \N__9379\
        );

    \I__2115\ : InMux
    port map (
            O => \N__9382\,
            I => \N__9373\
        );

    \I__2114\ : InMux
    port map (
            O => \N__9379\,
            I => \N__9373\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9378\,
            I => \N__9370\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__9373\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__9370\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__2110\ : IoInMux
    port map (
            O => \N__9365\,
            I => \N__9362\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__9362\,
            I => \N__9359\
        );

    \I__2108\ : Span4Mux_s3_v
    port map (
            O => \N__9359\,
            I => \N__9356\
        );

    \I__2107\ : Span4Mux_h
    port map (
            O => \N__9356\,
            I => \N__9353\
        );

    \I__2106\ : Sp12to4
    port map (
            O => \N__9353\,
            I => \N__9349\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9352\,
            I => \N__9346\
        );

    \I__2104\ : Odrv12
    port map (
            O => \N__9349\,
            I => \TICK60_c\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__9346\,
            I => \TICK60_c\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9341\,
            I => \N__9338\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9338\,
            I => \N__9335\
        );

    \I__2100\ : Span4Mux_h
    port map (
            O => \N__9335\,
            I => \N__9332\
        );

    \I__2099\ : Span4Mux_v
    port map (
            O => \N__9332\,
            I => \N__9329\
        );

    \I__2098\ : Span4Mux_v
    port map (
            O => \N__9329\,
            I => \N__9325\
        );

    \I__2097\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9322\
        );

    \I__2096\ : Sp12to4
    port map (
            O => \N__9325\,
            I => \N__9317\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__9322\,
            I => \N__9317\
        );

    \I__2094\ : Odrv12
    port map (
            O => \N__9317\,
            I => \CIA_SPACE\
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__9314\,
            I => \U409_CIA.VMA_RNOZ0Z_0_cascade_\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__9311\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9305\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9305\,
            I => \U409_TICK.TICK503_8\
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__9302\,
            I => \U409_TICK.TICK503_11_cascade_\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__9299\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9296\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__2086\ : InMux
    port map (
            O => \N__9293\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__2085\ : InMux
    port map (
            O => \N__9290\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__2084\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9283\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9286\,
            I => \N__9280\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__9283\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__9280\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__2080\ : InMux
    port map (
            O => \N__9275\,
            I => \N__9271\
        );

    \I__2079\ : InMux
    port map (
            O => \N__9274\,
            I => \N__9268\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__9271\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__9268\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__2076\ : CascadeMux
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9257\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__9257\,
            I => \N__9253\
        );

    \I__2073\ : InMux
    port map (
            O => \N__9256\,
            I => \N__9250\
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__9253\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__9250\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__2070\ : InMux
    port map (
            O => \N__9245\,
            I => \N__9242\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__9242\,
            I => \N__9237\
        );

    \I__2068\ : InMux
    port map (
            O => \N__9241\,
            I => \N__9234\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9240\,
            I => \N__9231\
        );

    \I__2066\ : Odrv12
    port map (
            O => \N__9237\,
            I => \U409_ADDRESS_DECODE.ATA_ENZ0\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9234\,
            I => \U409_ADDRESS_DECODE.ATA_ENZ0\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__9231\,
            I => \U409_ADDRESS_DECODE.ATA_ENZ0\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9221\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9221\,
            I => \N__9217\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9214\
        );

    \I__2060\ : Span4Mux_v
    port map (
            O => \N__9217\,
            I => \N__9210\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__9214\,
            I => \N__9207\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9213\,
            I => \N__9204\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__9210\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__9207\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__9204\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0\
        );

    \I__2054\ : IoInMux
    port map (
            O => \N__9197\,
            I => \N__9194\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9194\,
            I => \N__9191\
        );

    \I__2052\ : IoSpan4Mux
    port map (
            O => \N__9191\,
            I => \N__9188\
        );

    \I__2051\ : Sp12to4
    port map (
            O => \N__9188\,
            I => \N__9185\
        );

    \I__2050\ : Span12Mux_s7_h
    port map (
            O => \N__9185\,
            I => \N__9182\
        );

    \I__2049\ : Odrv12
    port map (
            O => \N__9182\,
            I => \U409_ADDRESS_DECODE_un1_ATA_ENn_i\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__9179\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9176\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9173\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9170\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9167\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9164\,
            I => \bfn_13_7_0_\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9161\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9158\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9155\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9152\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__9149\,
            I => \AGNUS_SPACE_0_cascade_\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9146\,
            I => \N__9143\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9143\,
            I => \N__9140\
        );

    \I__2035\ : Span12Mux_v
    port map (
            O => \N__9140\,
            I => \N__9137\
        );

    \I__2034\ : Span12Mux_h
    port map (
            O => \N__9137\,
            I => \N__9134\
        );

    \I__2033\ : Odrv12
    port map (
            O => \N__9134\,
            I => \TACKn_in\
        );

    \I__2032\ : SRMux
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9128\,
            I => \N__9122\
        );

    \I__2030\ : SRMux
    port map (
            O => \N__9127\,
            I => \N__9119\
        );

    \I__2029\ : SRMux
    port map (
            O => \N__9126\,
            I => \N__9116\
        );

    \I__2028\ : SRMux
    port map (
            O => \N__9125\,
            I => \N__9113\
        );

    \I__2027\ : Span4Mux_v
    port map (
            O => \N__9122\,
            I => \N__9108\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__9119\,
            I => \N__9108\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__9116\,
            I => \N__9105\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9113\,
            I => \N__9100\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__9108\,
            I => \N__9100\
        );

    \I__2022\ : Span4Mux_v
    port map (
            O => \N__9105\,
            I => \N__9095\
        );

    \I__2021\ : Span4Mux_v
    port map (
            O => \N__9100\,
            I => \N__9095\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__9095\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9088\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9085\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__9088\,
            I => \N__9079\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9085\,
            I => \N__9079\
        );

    \I__2015\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9076\
        );

    \I__2014\ : Span4Mux_h
    port map (
            O => \N__9079\,
            I => \N__9071\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__9076\,
            I => \N__9071\
        );

    \I__2012\ : Span4Mux_v
    port map (
            O => \N__9071\,
            I => \N__9066\
        );

    \I__2011\ : InMux
    port map (
            O => \N__9070\,
            I => \N__9063\
        );

    \I__2010\ : InMux
    port map (
            O => \N__9069\,
            I => \N__9060\
        );

    \I__2009\ : Odrv4
    port map (
            O => \N__9066\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__9063\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__9060\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__9053\,
            I => \N__9048\
        );

    \I__2005\ : InMux
    port map (
            O => \N__9052\,
            I => \N__9045\
        );

    \I__2004\ : InMux
    port map (
            O => \N__9051\,
            I => \N__9042\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9048\,
            I => \N__9039\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9045\,
            I => \N__9032\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__9042\,
            I => \N__9032\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9039\,
            I => \N__9032\
        );

    \I__1999\ : Span4Mux_h
    port map (
            O => \N__9032\,
            I => \N__9029\
        );

    \I__1998\ : Span4Mux_v
    port map (
            O => \N__9029\,
            I => \N__9024\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9028\,
            I => \N__9021\
        );

    \I__1996\ : InMux
    port map (
            O => \N__9027\,
            I => \N__9018\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__9024\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__9021\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9018\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4\
        );

    \I__1992\ : IoInMux
    port map (
            O => \N__9011\,
            I => \N__9008\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__9008\,
            I => \N__9005\
        );

    \I__1990\ : IoSpan4Mux
    port map (
            O => \N__9005\,
            I => \N__9002\
        );

    \I__1989\ : Span4Mux_s3_v
    port map (
            O => \N__9002\,
            I => \N__8999\
        );

    \I__1988\ : Sp12to4
    port map (
            O => \N__8999\,
            I => \N__8996\
        );

    \I__1987\ : Span12Mux_h
    port map (
            O => \N__8996\,
            I => \N__8993\
        );

    \I__1986\ : Odrv12
    port map (
            O => \N__8993\,
            I => \BUFENn_c\
        );

    \I__1985\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8987\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__8987\,
            I => \N__8984\
        );

    \I__1983\ : Odrv12
    port map (
            O => \N__8984\,
            I => \U409_ADDRESS_DECODE_PORTSIZE_0\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__8981\,
            I => \N__8977\
        );

    \I__1981\ : InMux
    port map (
            O => \N__8980\,
            I => \N__8972\
        );

    \I__1980\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8972\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__8972\,
            I => \AGNUS_SPACE_0\
        );

    \I__1978\ : IoInMux
    port map (
            O => \N__8969\,
            I => \N__8966\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__8966\,
            I => \N__8963\
        );

    \I__1976\ : IoSpan4Mux
    port map (
            O => \N__8963\,
            I => \N__8960\
        );

    \I__1975\ : Span4Mux_s0_v
    port map (
            O => \N__8960\,
            I => \N__8956\
        );

    \I__1974\ : IoInMux
    port map (
            O => \N__8959\,
            I => \N__8953\
        );

    \I__1973\ : Sp12to4
    port map (
            O => \N__8956\,
            I => \N__8948\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__8953\,
            I => \N__8948\
        );

    \I__1971\ : Span12Mux_s11_v
    port map (
            O => \N__8948\,
            I => \N__8943\
        );

    \I__1970\ : InMux
    port map (
            O => \N__8947\,
            I => \N__8940\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__8946\,
            I => \N__8937\
        );

    \I__1968\ : Span12Mux_h
    port map (
            O => \N__8943\,
            I => \N__8934\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__8940\,
            I => \N__8931\
        );

    \I__1966\ : InMux
    port map (
            O => \N__8937\,
            I => \N__8928\
        );

    \I__1965\ : Odrv12
    port map (
            O => \N__8934\,
            I => \TACK_EN\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__8931\,
            I => \TACK_EN\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__8928\,
            I => \TACK_EN\
        );

    \I__1962\ : IoInMux
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__8918\,
            I => \N__8915\
        );

    \I__1960\ : IoSpan4Mux
    port map (
            O => \N__8915\,
            I => \N__8912\
        );

    \I__1959\ : Span4Mux_s2_v
    port map (
            O => \N__8912\,
            I => \N__8909\
        );

    \I__1958\ : Sp12to4
    port map (
            O => \N__8909\,
            I => \N__8906\
        );

    \I__1957\ : Span12Mux_h
    port map (
            O => \N__8906\,
            I => \N__8903\
        );

    \I__1956\ : Odrv12
    port map (
            O => \N__8903\,
            I => \TCIn_1_i\
        );

    \I__1955\ : IoInMux
    port map (
            O => \N__8900\,
            I => \N__8897\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__8897\,
            I => \N__8894\
        );

    \I__1953\ : Span12Mux_s2_v
    port map (
            O => \N__8894\,
            I => \N__8891\
        );

    \I__1952\ : Odrv12
    port map (
            O => \N__8891\,
            I => \RESETn_c_i\
        );

    \I__1951\ : InMux
    port map (
            O => \N__8888\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8885\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__1949\ : InMux
    port map (
            O => \N__8882\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__1948\ : IoInMux
    port map (
            O => \N__8879\,
            I => \N__8876\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__8876\,
            I => \N__8873\
        );

    \I__1946\ : Span12Mux_s7_v
    port map (
            O => \N__8873\,
            I => \N__8870\
        );

    \I__1945\ : Odrv12
    port map (
            O => \N__8870\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8867\,
            I => \N__8864\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__8864\,
            I => \U409_TRANSFER_ACK.N_28\
        );

    \I__1942\ : InMux
    port map (
            O => \N__8861\,
            I => \N__8858\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__8858\,
            I => \N__8855\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__8855\,
            I => \N__8851\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8854\,
            I => \N__8848\
        );

    \I__1938\ : Odrv4
    port map (
            O => \N__8851\,
            I => \U409_TRANSFER_ACK.N_22\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__8848\,
            I => \U409_TRANSFER_ACK.N_22\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__8843\,
            I => \N__8839\
        );

    \I__1935\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8836\
        );

    \I__1934\ : InMux
    port map (
            O => \N__8839\,
            I => \N__8832\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__8836\,
            I => \N__8829\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8835\,
            I => \N__8826\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__8832\,
            I => \N__8822\
        );

    \I__1930\ : Span4Mux_h
    port map (
            O => \N__8829\,
            I => \N__8817\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__8826\,
            I => \N__8817\
        );

    \I__1928\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8814\
        );

    \I__1927\ : Span12Mux_v
    port map (
            O => \N__8822\,
            I => \N__8811\
        );

    \I__1926\ : Span4Mux_h
    port map (
            O => \N__8817\,
            I => \N__8808\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__8814\,
            I => \N__8805\
        );

    \I__1924\ : Odrv12
    port map (
            O => \N__8811\,
            I => \U409_ADDRESS_DECODE_ROMEN_1\
        );

    \I__1923\ : Odrv4
    port map (
            O => \N__8808\,
            I => \U409_ADDRESS_DECODE_ROMEN_1\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__8805\,
            I => \U409_ADDRESS_DECODE_ROMEN_1\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8798\,
            I => \N__8795\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__8795\,
            I => \N__8791\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__8794\,
            I => \N__8788\
        );

    \I__1918\ : Span4Mux_h
    port map (
            O => \N__8791\,
            I => \N__8785\
        );

    \I__1917\ : InMux
    port map (
            O => \N__8788\,
            I => \N__8782\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__8785\,
            I => \U409_TRANSFER_ACK.N_33_1\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__8782\,
            I => \U409_TRANSFER_ACK.N_33_1\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__8777\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0_cascade_\
        );

    \I__1913\ : InMux
    port map (
            O => \N__8774\,
            I => \N__8771\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__8771\,
            I => \U409_TRANSFER_ACK.N_33\
        );

    \I__1911\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8753\
        );

    \I__1910\ : InMux
    port map (
            O => \N__8767\,
            I => \N__8753\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8766\,
            I => \N__8753\
        );

    \I__1908\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8753\
        );

    \I__1907\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8746\
        );

    \I__1906\ : InMux
    port map (
            O => \N__8763\,
            I => \N__8746\
        );

    \I__1905\ : InMux
    port map (
            O => \N__8762\,
            I => \N__8746\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8753\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__8746\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__8741\,
            I => \N__8734\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__8740\,
            I => \N__8731\
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__8739\,
            I => \N__8727\
        );

    \I__1899\ : InMux
    port map (
            O => \N__8738\,
            I => \N__8715\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8737\,
            I => \N__8715\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8734\,
            I => \N__8715\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8731\,
            I => \N__8715\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8730\,
            I => \N__8715\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8727\,
            I => \N__8710\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8726\,
            I => \N__8710\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__8715\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__8710\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8705\,
            I => \N__8702\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__8702\,
            I => \U409_TRANSFER_ACK.N_34\
        );

    \I__1888\ : InMux
    port map (
            O => \N__8699\,
            I => \N__8689\
        );

    \I__1887\ : InMux
    port map (
            O => \N__8698\,
            I => \N__8689\
        );

    \I__1886\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8680\
        );

    \I__1885\ : InMux
    port map (
            O => \N__8696\,
            I => \N__8680\
        );

    \I__1884\ : InMux
    port map (
            O => \N__8695\,
            I => \N__8680\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8680\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__8689\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__8680\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__8675\,
            I => \N__8667\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__8674\,
            I => \N__8664\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8673\,
            I => \N__8658\
        );

    \I__1877\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8658\
        );

    \I__1876\ : InMux
    port map (
            O => \N__8671\,
            I => \N__8655\
        );

    \I__1875\ : InMux
    port map (
            O => \N__8670\,
            I => \N__8646\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8646\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8646\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8646\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8658\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8655\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__8646\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8636\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8636\,
            I => \N__8633\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__8633\,
            I => \U409_TRANSFER_ACK.N_45\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8630\,
            I => \N__8624\
        );

    \I__1864\ : InMux
    port map (
            O => \N__8629\,
            I => \N__8621\
        );

    \I__1863\ : InMux
    port map (
            O => \N__8628\,
            I => \N__8616\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8627\,
            I => \N__8616\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8624\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8621\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__8616\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8605\
        );

    \I__1857\ : InMux
    port map (
            O => \N__8608\,
            I => \N__8602\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8605\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__8602\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1854\ : InMux
    port map (
            O => \N__8597\,
            I => \N__8591\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8596\,
            I => \N__8588\
        );

    \I__1852\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8583\
        );

    \I__1851\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8583\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8591\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8588\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8583\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1847\ : SRMux
    port map (
            O => \N__8576\,
            I => \N__8546\
        );

    \I__1846\ : SRMux
    port map (
            O => \N__8575\,
            I => \N__8546\
        );

    \I__1845\ : SRMux
    port map (
            O => \N__8574\,
            I => \N__8546\
        );

    \I__1844\ : SRMux
    port map (
            O => \N__8573\,
            I => \N__8546\
        );

    \I__1843\ : SRMux
    port map (
            O => \N__8572\,
            I => \N__8546\
        );

    \I__1842\ : SRMux
    port map (
            O => \N__8571\,
            I => \N__8546\
        );

    \I__1841\ : SRMux
    port map (
            O => \N__8570\,
            I => \N__8546\
        );

    \I__1840\ : SRMux
    port map (
            O => \N__8569\,
            I => \N__8546\
        );

    \I__1839\ : SRMux
    port map (
            O => \N__8568\,
            I => \N__8546\
        );

    \I__1838\ : SRMux
    port map (
            O => \N__8567\,
            I => \N__8546\
        );

    \I__1837\ : GlobalMux
    port map (
            O => \N__8546\,
            I => \N__8543\
        );

    \I__1836\ : gio2CtrlBuf
    port map (
            O => \N__8543\,
            I => \RESETn_c_i_g\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8540\,
            I => \N__8536\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8539\,
            I => \N__8533\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__8536\,
            I => \N__8530\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8533\,
            I => \N__8527\
        );

    \I__1831\ : Span4Mux_h
    port map (
            O => \N__8530\,
            I => \N__8522\
        );

    \I__1830\ : Span4Mux_v
    port map (
            O => \N__8527\,
            I => \N__8522\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__8522\,
            I => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8516\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8516\,
            I => \N__8513\
        );

    \I__1826\ : Span4Mux_v
    port map (
            O => \N__8513\,
            I => \N__8509\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8506\
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__8509\,
            I => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8506\,
            I => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8497\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__8500\,
            I => \N__8494\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8497\,
            I => \N__8488\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8494\,
            I => \N__8485\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8493\,
            I => \N__8480\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8480\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8491\,
            I => \N__8476\
        );

    \I__1815\ : Span4Mux_v
    port map (
            O => \N__8488\,
            I => \N__8467\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8485\,
            I => \N__8467\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8480\,
            I => \N__8464\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8479\,
            I => \N__8461\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8476\,
            I => \N__8458\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8451\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8451\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8473\,
            I => \N__8451\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__8472\,
            I => \N__8447\
        );

    \I__1806\ : Span4Mux_v
    port map (
            O => \N__8467\,
            I => \N__8444\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__8464\,
            I => \N__8439\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__8461\,
            I => \N__8439\
        );

    \I__1803\ : Span4Mux_v
    port map (
            O => \N__8458\,
            I => \N__8434\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8451\,
            I => \N__8434\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8431\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8447\,
            I => \N__8428\
        );

    \I__1799\ : Span4Mux_h
    port map (
            O => \N__8444\,
            I => \N__8423\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__8439\,
            I => \N__8423\
        );

    \I__1797\ : Span4Mux_v
    port map (
            O => \N__8434\,
            I => \N__8420\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8431\,
            I => \N__8417\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__8428\,
            I => \N__8414\
        );

    \I__1794\ : Span4Mux_h
    port map (
            O => \N__8423\,
            I => \N__8411\
        );

    \I__1793\ : Span4Mux_h
    port map (
            O => \N__8420\,
            I => \N__8406\
        );

    \I__1792\ : Span4Mux_v
    port map (
            O => \N__8417\,
            I => \N__8406\
        );

    \I__1791\ : Span12Mux_v
    port map (
            O => \N__8414\,
            I => \N__8401\
        );

    \I__1790\ : Sp12to4
    port map (
            O => \N__8411\,
            I => \N__8401\
        );

    \I__1789\ : Span4Mux_h
    port map (
            O => \N__8406\,
            I => \N__8398\
        );

    \I__1788\ : Odrv12
    port map (
            O => \N__8401\,
            I => \A_c_21\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__8398\,
            I => \A_c_21\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__8390\,
            I => \N__8386\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8383\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__8386\,
            I => \N__8377\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8383\,
            I => \N__8377\
        );

    \I__1781\ : InMux
    port map (
            O => \N__8382\,
            I => \N__8374\
        );

    \I__1780\ : Sp12to4
    port map (
            O => \N__8377\,
            I => \N__8369\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8374\,
            I => \N__8369\
        );

    \I__1778\ : Span12Mux_v
    port map (
            O => \N__8369\,
            I => \N__8366\
        );

    \I__1777\ : Span12Mux_h
    port map (
            O => \N__8366\,
            I => \N__8363\
        );

    \I__1776\ : Odrv12
    port map (
            O => \N__8363\,
            I => \OVL_c\
        );

    \I__1775\ : CascadeMux
    port map (
            O => \N__8360\,
            I => \N__8356\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__8359\,
            I => \N__8353\
        );

    \I__1773\ : InMux
    port map (
            O => \N__8356\,
            I => \N__8347\
        );

    \I__1772\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8342\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8352\,
            I => \N__8342\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8351\,
            I => \N__8337\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8337\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8347\,
            I => \N__8334\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__8342\,
            I => \N__8328\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__8337\,
            I => \N__8328\
        );

    \I__1765\ : Span4Mux_v
    port map (
            O => \N__8334\,
            I => \N__8324\
        );

    \I__1764\ : InMux
    port map (
            O => \N__8333\,
            I => \N__8321\
        );

    \I__1763\ : Span4Mux_h
    port map (
            O => \N__8328\,
            I => \N__8318\
        );

    \I__1762\ : InMux
    port map (
            O => \N__8327\,
            I => \N__8315\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__8324\,
            I => \CONFIGURED\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__8321\,
            I => \CONFIGURED\
        );

    \I__1759\ : Odrv4
    port map (
            O => \N__8318\,
            I => \CONFIGURED\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__8315\,
            I => \CONFIGURED\
        );

    \I__1757\ : InMux
    port map (
            O => \N__8306\,
            I => \N__8303\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8303\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8300\,
            I => \N__8297\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8297\,
            I => \N__8294\
        );

    \I__1753\ : Span4Mux_v
    port map (
            O => \N__8294\,
            I => \N__8291\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__8291\,
            I => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_1\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8288\,
            I => \N__8285\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__8285\,
            I => \N__8282\
        );

    \I__1749\ : Odrv4
    port map (
            O => \N__8282\,
            I => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_2\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__8279\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_\
        );

    \I__1747\ : IoInMux
    port map (
            O => \N__8276\,
            I => \N__8273\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__8273\,
            I => \N__8270\
        );

    \I__1745\ : Span12Mux_s5_h
    port map (
            O => \N__8270\,
            I => \N__8267\
        );

    \I__1744\ : Span12Mux_h
    port map (
            O => \N__8267\,
            I => \N__8264\
        );

    \I__1743\ : Odrv12
    port map (
            O => \N__8264\,
            I => \U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8254\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8260\,
            I => \N__8249\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8259\,
            I => \N__8246\
        );

    \I__1739\ : InMux
    port map (
            O => \N__8258\,
            I => \N__8243\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8240\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__8254\,
            I => \N__8237\
        );

    \I__1736\ : InMux
    port map (
            O => \N__8253\,
            I => \N__8234\
        );

    \I__1735\ : InMux
    port map (
            O => \N__8252\,
            I => \N__8231\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__8249\,
            I => \N__8226\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8246\,
            I => \N__8226\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__8243\,
            I => \N__8221\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__8240\,
            I => \N__8221\
        );

    \I__1730\ : Span4Mux_v
    port map (
            O => \N__8237\,
            I => \N__8214\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8234\,
            I => \N__8214\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__8231\,
            I => \N__8214\
        );

    \I__1727\ : Span4Mux_v
    port map (
            O => \N__8226\,
            I => \N__8211\
        );

    \I__1726\ : Span4Mux_v
    port map (
            O => \N__8221\,
            I => \N__8206\
        );

    \I__1725\ : Span4Mux_v
    port map (
            O => \N__8214\,
            I => \N__8206\
        );

    \I__1724\ : Sp12to4
    port map (
            O => \N__8211\,
            I => \N__8201\
        );

    \I__1723\ : Sp12to4
    port map (
            O => \N__8206\,
            I => \N__8201\
        );

    \I__1722\ : Span12Mux_h
    port map (
            O => \N__8201\,
            I => \N__8198\
        );

    \I__1721\ : Span12Mux_v
    port map (
            O => \N__8198\,
            I => \N__8195\
        );

    \I__1720\ : Odrv12
    port map (
            O => \N__8195\,
            I => \RnW_c\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8192\,
            I => \N__8187\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__8191\,
            I => \N__8184\
        );

    \I__1717\ : InMux
    port map (
            O => \N__8190\,
            I => \N__8181\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__8187\,
            I => \N__8178\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8184\,
            I => \N__8175\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8181\,
            I => \N__8172\
        );

    \I__1713\ : Span4Mux_h
    port map (
            O => \N__8178\,
            I => \N__8169\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__8175\,
            I => \N__8164\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__8172\,
            I => \N__8164\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__8169\,
            I => \N__8161\
        );

    \I__1709\ : Sp12to4
    port map (
            O => \N__8164\,
            I => \N__8158\
        );

    \I__1708\ : Sp12to4
    port map (
            O => \N__8161\,
            I => \N__8153\
        );

    \I__1707\ : Span12Mux_h
    port map (
            O => \N__8158\,
            I => \N__8153\
        );

    \I__1706\ : Span12Mux_v
    port map (
            O => \N__8153\,
            I => \N__8150\
        );

    \I__1705\ : Odrv12
    port map (
            O => \N__8150\,
            I => \D_in_5\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__8147\,
            I => \un1_AUTOCONFIG_SPACE_cascade_\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8144\,
            I => \N__8140\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8143\,
            I => \N__8137\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8140\,
            I => \ATA_BASE_1\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8137\,
            I => \ATA_BASE_1\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8132\,
            I => \N__8125\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8125\
        );

    \I__1697\ : InMux
    port map (
            O => \N__8130\,
            I => \N__8122\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__8125\,
            I => \U409_AUTOCONFIG.STATE_RNIS3FU2Z0Z_0\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8122\,
            I => \U409_AUTOCONFIG.STATE_RNIS3FU2Z0Z_0\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8117\,
            I => \N__8108\
        );

    \I__1693\ : InMux
    port map (
            O => \N__8116\,
            I => \N__8108\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__8115\,
            I => \N__8104\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__8114\,
            I => \N__8101\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__8113\,
            I => \N__8098\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__8108\,
            I => \N__8092\
        );

    \I__1688\ : InMux
    port map (
            O => \N__8107\,
            I => \N__8081\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8104\,
            I => \N__8081\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8101\,
            I => \N__8081\
        );

    \I__1685\ : InMux
    port map (
            O => \N__8098\,
            I => \N__8081\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8081\
        );

    \I__1683\ : InMux
    port map (
            O => \N__8096\,
            I => \N__8076\
        );

    \I__1682\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8076\
        );

    \I__1681\ : Span4Mux_h
    port map (
            O => \N__8092\,
            I => \N__8071\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__8081\,
            I => \N__8071\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8076\,
            I => \N__8067\
        );

    \I__1678\ : Span4Mux_h
    port map (
            O => \N__8071\,
            I => \N__8064\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8070\,
            I => \N__8061\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__8067\,
            I => \un1_AUTOCONFIG_SPACE\
        );

    \I__1675\ : Odrv4
    port map (
            O => \N__8064\,
            I => \un1_AUTOCONFIG_SPACE\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8061\,
            I => \un1_AUTOCONFIG_SPACE\
        );

    \I__1673\ : CascadeMux
    port map (
            O => \N__8054\,
            I => \N__8050\
        );

    \I__1672\ : InMux
    port map (
            O => \N__8053\,
            I => \N__8047\
        );

    \I__1671\ : InMux
    port map (
            O => \N__8050\,
            I => \N__8044\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8047\,
            I => \N__8039\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8044\,
            I => \N__8039\
        );

    \I__1668\ : Span4Mux_v
    port map (
            O => \N__8039\,
            I => \N__8035\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__8038\,
            I => \N__8032\
        );

    \I__1666\ : Span4Mux_h
    port map (
            O => \N__8035\,
            I => \N__8029\
        );

    \I__1665\ : InMux
    port map (
            O => \N__8032\,
            I => \N__8026\
        );

    \I__1664\ : Sp12to4
    port map (
            O => \N__8029\,
            I => \N__8021\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__8026\,
            I => \N__8021\
        );

    \I__1662\ : Span12Mux_v
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__1661\ : Odrv12
    port map (
            O => \N__8018\,
            I => \D_in_7\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8015\,
            I => \N__8011\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8014\,
            I => \N__8008\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__8011\,
            I => \ATA_BASE_3\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__8008\,
            I => \ATA_BASE_3\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__8003\,
            I => \N__7994\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__8002\,
            I => \N__7991\
        );

    \I__1654\ : InMux
    port map (
            O => \N__8001\,
            I => \N__7988\
        );

    \I__1653\ : InMux
    port map (
            O => \N__8000\,
            I => \N__7985\
        );

    \I__1652\ : InMux
    port map (
            O => \N__7999\,
            I => \N__7982\
        );

    \I__1651\ : InMux
    port map (
            O => \N__7998\,
            I => \N__7979\
        );

    \I__1650\ : InMux
    port map (
            O => \N__7997\,
            I => \N__7976\
        );

    \I__1649\ : InMux
    port map (
            O => \N__7994\,
            I => \N__7971\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7991\,
            I => \N__7971\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__7988\,
            I => \N__7968\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__7985\,
            I => \N__7965\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__7982\,
            I => \N__7960\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7979\,
            I => \N__7957\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7976\,
            I => \N__7952\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__7971\,
            I => \N__7944\
        );

    \I__1641\ : Glb2LocalMux
    port map (
            O => \N__7968\,
            I => \N__7910\
        );

    \I__1640\ : Glb2LocalMux
    port map (
            O => \N__7965\,
            I => \N__7910\
        );

    \I__1639\ : ClkMux
    port map (
            O => \N__7964\,
            I => \N__7910\
        );

    \I__1638\ : ClkMux
    port map (
            O => \N__7963\,
            I => \N__7910\
        );

    \I__1637\ : Glb2LocalMux
    port map (
            O => \N__7960\,
            I => \N__7910\
        );

    \I__1636\ : Glb2LocalMux
    port map (
            O => \N__7957\,
            I => \N__7910\
        );

    \I__1635\ : ClkMux
    port map (
            O => \N__7956\,
            I => \N__7910\
        );

    \I__1634\ : ClkMux
    port map (
            O => \N__7955\,
            I => \N__7910\
        );

    \I__1633\ : Glb2LocalMux
    port map (
            O => \N__7952\,
            I => \N__7910\
        );

    \I__1632\ : ClkMux
    port map (
            O => \N__7951\,
            I => \N__7910\
        );

    \I__1631\ : ClkMux
    port map (
            O => \N__7950\,
            I => \N__7910\
        );

    \I__1630\ : ClkMux
    port map (
            O => \N__7949\,
            I => \N__7910\
        );

    \I__1629\ : ClkMux
    port map (
            O => \N__7948\,
            I => \N__7910\
        );

    \I__1628\ : ClkMux
    port map (
            O => \N__7947\,
            I => \N__7910\
        );

    \I__1627\ : Glb2LocalMux
    port map (
            O => \N__7944\,
            I => \N__7910\
        );

    \I__1626\ : ClkMux
    port map (
            O => \N__7943\,
            I => \N__7910\
        );

    \I__1625\ : GlobalMux
    port map (
            O => \N__7910\,
            I => \N__7907\
        );

    \I__1624\ : gio2CtrlBuf
    port map (
            O => \N__7907\,
            I => \CLK40_IN_c_g\
        );

    \I__1623\ : IoInMux
    port map (
            O => \N__7904\,
            I => \N__7901\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__7901\,
            I => \N__7898\
        );

    \I__1621\ : Span12Mux_s6_v
    port map (
            O => \N__7898\,
            I => \N__7895\
        );

    \I__1620\ : Odrv12
    port map (
            O => \N__7895\,
            I => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\
        );

    \I__1619\ : InMux
    port map (
            O => \N__7892\,
            I => \N__7886\
        );

    \I__1618\ : InMux
    port map (
            O => \N__7891\,
            I => \N__7879\
        );

    \I__1617\ : InMux
    port map (
            O => \N__7890\,
            I => \N__7879\
        );

    \I__1616\ : InMux
    port map (
            O => \N__7889\,
            I => \N__7879\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__7886\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__7879\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1613\ : InMux
    port map (
            O => \N__7874\,
            I => \N__7869\
        );

    \I__1612\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7864\
        );

    \I__1611\ : InMux
    port map (
            O => \N__7872\,
            I => \N__7864\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__7869\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__7864\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__1608\ : IoInMux
    port map (
            O => \N__7859\,
            I => \N__7856\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__7856\,
            I => \N__7853\
        );

    \I__1606\ : Span4Mux_s3_v
    port map (
            O => \N__7853\,
            I => \N__7850\
        );

    \I__1605\ : Span4Mux_v
    port map (
            O => \N__7850\,
            I => \N__7847\
        );

    \I__1604\ : Span4Mux_v
    port map (
            O => \N__7847\,
            I => \N__7844\
        );

    \I__1603\ : Span4Mux_h
    port map (
            O => \N__7844\,
            I => \N__7840\
        );

    \I__1602\ : InMux
    port map (
            O => \N__7843\,
            I => \N__7837\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__7840\,
            I => \TICK50_c\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7837\,
            I => \TICK50_c\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7832\,
            I => \N__7829\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__7829\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__7826\,
            I => \N__7823\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7819\
        );

    \I__1595\ : InMux
    port map (
            O => \N__7822\,
            I => \N__7816\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__7819\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__7816\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1592\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7807\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7804\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__7807\,
            I => \N__7801\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7804\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1588\ : Odrv12
    port map (
            O => \N__7801\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__7796\,
            I => \N__7793\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7793\,
            I => \N__7789\
        );

    \I__1585\ : CascadeMux
    port map (
            O => \N__7792\,
            I => \N__7786\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7789\,
            I => \N__7783\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7786\,
            I => \N__7780\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__7783\,
            I => \AC_TACK\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__7780\,
            I => \AC_TACK\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7772\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__7772\,
            I => \N__7769\
        );

    \I__1578\ : Span4Mux_h
    port map (
            O => \N__7769\,
            I => \N__7766\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__7766\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER5_1\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__7763\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__7760\,
            I => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\
        );

    \I__1574\ : IoInMux
    port map (
            O => \N__7757\,
            I => \N__7753\
        );

    \I__1573\ : IoInMux
    port map (
            O => \N__7756\,
            I => \N__7750\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__7753\,
            I => \N__7744\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__7750\,
            I => \N__7744\
        );

    \I__1570\ : IoInMux
    port map (
            O => \N__7749\,
            I => \N__7741\
        );

    \I__1569\ : IoSpan4Mux
    port map (
            O => \N__7744\,
            I => \N__7738\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7741\,
            I => \N__7735\
        );

    \I__1567\ : Span4Mux_s2_v
    port map (
            O => \N__7738\,
            I => \N__7730\
        );

    \I__1566\ : Span4Mux_s2_v
    port map (
            O => \N__7735\,
            I => \N__7730\
        );

    \I__1565\ : Span4Mux_v
    port map (
            O => \N__7730\,
            I => \N__7727\
        );

    \I__1564\ : Sp12to4
    port map (
            O => \N__7727\,
            I => \N__7724\
        );

    \I__1563\ : Span12Mux_h
    port map (
            O => \N__7724\,
            I => \N__7719\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7723\,
            I => \N__7714\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7722\,
            I => \N__7714\
        );

    \I__1560\ : Odrv12
    port map (
            O => \N__7719\,
            I => \TACK_OUTn\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7714\,
            I => \TACK_OUTn\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__7709\,
            I => \N__7703\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__7708\,
            I => \N__7699\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7707\,
            I => \N__7695\
        );

    \I__1555\ : InMux
    port map (
            O => \N__7706\,
            I => \N__7692\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7683\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7702\,
            I => \N__7683\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7699\,
            I => \N__7683\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7698\,
            I => \N__7683\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7695\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7692\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7683\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7676\,
            I => \N__7670\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7675\,
            I => \N__7667\
        );

    \I__1545\ : InMux
    port map (
            O => \N__7674\,
            I => \N__7662\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7673\,
            I => \N__7662\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__7670\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__7667\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__7662\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7655\,
            I => \N__7651\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7654\,
            I => \N__7648\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7651\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_1_out\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__7648\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_1_out\
        );

    \I__1536\ : InMux
    port map (
            O => \N__7643\,
            I => \N__7640\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__7640\,
            I => \N__7636\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__7639\,
            I => \N__7633\
        );

    \I__1533\ : Span4Mux_h
    port map (
            O => \N__7636\,
            I => \N__7629\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7633\,
            I => \N__7624\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7632\,
            I => \N__7624\
        );

    \I__1530\ : Span4Mux_h
    port map (
            O => \N__7629\,
            I => \N__7619\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__7624\,
            I => \N__7619\
        );

    \I__1528\ : Span4Mux_h
    port map (
            O => \N__7619\,
            I => \N__7616\
        );

    \I__1527\ : Span4Mux_v
    port map (
            O => \N__7616\,
            I => \N__7613\
        );

    \I__1526\ : Span4Mux_v
    port map (
            O => \N__7613\,
            I => \N__7610\
        );

    \I__1525\ : Span4Mux_v
    port map (
            O => \N__7610\,
            I => \N__7607\
        );

    \I__1524\ : Odrv4
    port map (
            O => \N__7607\,
            I => \TM_c_0\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7604\,
            I => \N__7601\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7601\,
            I => \N__7596\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7600\,
            I => \N__7591\
        );

    \I__1520\ : InMux
    port map (
            O => \N__7599\,
            I => \N__7591\
        );

    \I__1519\ : Span4Mux_v
    port map (
            O => \N__7596\,
            I => \N__7588\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7591\,
            I => \N__7585\
        );

    \I__1517\ : Span4Mux_h
    port map (
            O => \N__7588\,
            I => \N__7580\
        );

    \I__1516\ : Span4Mux_v
    port map (
            O => \N__7585\,
            I => \N__7580\
        );

    \I__1515\ : Span4Mux_h
    port map (
            O => \N__7580\,
            I => \N__7577\
        );

    \I__1514\ : Sp12to4
    port map (
            O => \N__7577\,
            I => \N__7574\
        );

    \I__1513\ : Odrv12
    port map (
            O => \N__7574\,
            I => \TM_c_1\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7566\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7561\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7561\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__7566\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7561\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7556\,
            I => \N__7550\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7555\,
            I => \N__7550\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7550\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__7547\,
            I => \N__7541\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7546\,
            I => \N__7537\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7528\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7544\,
            I => \N__7528\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7541\,
            I => \N__7528\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7540\,
            I => \N__7528\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7537\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7528\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7520\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7520\,
            I => \U409_TRANSFER_ACK.N_17_mux\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__7517\,
            I => \N__7512\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7507\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7515\,
            I => \N__7507\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7504\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__7507\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7504\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7499\,
            I => \N__7496\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7496\,
            I => \N__7493\
        );

    \I__1486\ : Odrv12
    port map (
            O => \N__7493\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1Z0Z_0\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__7490\,
            I => \N__7487\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7487\,
            I => \N__7481\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7486\,
            I => \N__7481\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7481\,
            I => \N__7477\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__7480\,
            I => \N__7473\
        );

    \I__1480\ : Span4Mux_v
    port map (
            O => \N__7477\,
            I => \N__7470\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7476\,
            I => \N__7467\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7473\,
            I => \N__7464\
        );

    \I__1477\ : Span4Mux_h
    port map (
            O => \N__7470\,
            I => \N__7455\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7467\,
            I => \N__7455\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__7464\,
            I => \N__7455\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7463\,
            I => \N__7451\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__7462\,
            I => \N__7448\
        );

    \I__1472\ : Span4Mux_v
    port map (
            O => \N__7455\,
            I => \N__7445\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7454\,
            I => \N__7442\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7451\,
            I => \N__7438\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7448\,
            I => \N__7435\
        );

    \I__1468\ : Span4Mux_v
    port map (
            O => \N__7445\,
            I => \N__7430\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__7442\,
            I => \N__7430\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7427\
        );

    \I__1465\ : Span4Mux_v
    port map (
            O => \N__7438\,
            I => \N__7422\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7435\,
            I => \N__7422\
        );

    \I__1463\ : Span4Mux_h
    port map (
            O => \N__7430\,
            I => \N__7417\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7427\,
            I => \N__7417\
        );

    \I__1461\ : Span4Mux_v
    port map (
            O => \N__7422\,
            I => \N__7414\
        );

    \I__1460\ : Span4Mux_v
    port map (
            O => \N__7417\,
            I => \N__7411\
        );

    \I__1459\ : Sp12to4
    port map (
            O => \N__7414\,
            I => \N__7408\
        );

    \I__1458\ : Span4Mux_v
    port map (
            O => \N__7411\,
            I => \N__7405\
        );

    \I__1457\ : Span12Mux_v
    port map (
            O => \N__7408\,
            I => \N__7402\
        );

    \I__1456\ : Span4Mux_v
    port map (
            O => \N__7405\,
            I => \N__7399\
        );

    \I__1455\ : Span12Mux_h
    port map (
            O => \N__7402\,
            I => \N__7396\
        );

    \I__1454\ : Span4Mux_h
    port map (
            O => \N__7399\,
            I => \N__7393\
        );

    \I__1453\ : Odrv12
    port map (
            O => \N__7396\,
            I => \A_c_22\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__7393\,
            I => \A_c_22\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7388\,
            I => \N__7381\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7387\,
            I => \N__7381\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7377\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7381\,
            I => \N__7374\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7380\,
            I => \N__7371\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7377\,
            I => \N__7367\
        );

    \I__1445\ : Span4Mux_v
    port map (
            O => \N__7374\,
            I => \N__7362\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__7371\,
            I => \N__7362\
        );

    \I__1443\ : InMux
    port map (
            O => \N__7370\,
            I => \N__7359\
        );

    \I__1442\ : Span4Mux_v
    port map (
            O => \N__7367\,
            I => \N__7355\
        );

    \I__1441\ : Span4Mux_v
    port map (
            O => \N__7362\,
            I => \N__7351\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__7359\,
            I => \N__7348\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7358\,
            I => \N__7345\
        );

    \I__1438\ : Span4Mux_v
    port map (
            O => \N__7355\,
            I => \N__7342\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7354\,
            I => \N__7339\
        );

    \I__1436\ : Span4Mux_h
    port map (
            O => \N__7351\,
            I => \N__7334\
        );

    \I__1435\ : Span4Mux_v
    port map (
            O => \N__7348\,
            I => \N__7334\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__7345\,
            I => \N__7331\
        );

    \I__1433\ : Sp12to4
    port map (
            O => \N__7342\,
            I => \N__7326\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7339\,
            I => \N__7326\
        );

    \I__1431\ : Span4Mux_h
    port map (
            O => \N__7334\,
            I => \N__7321\
        );

    \I__1430\ : Span4Mux_v
    port map (
            O => \N__7331\,
            I => \N__7321\
        );

    \I__1429\ : Span12Mux_h
    port map (
            O => \N__7326\,
            I => \N__7316\
        );

    \I__1428\ : Sp12to4
    port map (
            O => \N__7321\,
            I => \N__7316\
        );

    \I__1427\ : Odrv12
    port map (
            O => \N__7316\,
            I => \A_c_23\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7313\,
            I => \N__7310\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7310\,
            I => \N__7307\
        );

    \I__1424\ : Odrv4
    port map (
            O => \N__7307\,
            I => \U409_TRANSFER_ACK.N_43\
        );

    \I__1423\ : IoInMux
    port map (
            O => \N__7304\,
            I => \N__7301\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7301\,
            I => \N__7298\
        );

    \I__1421\ : Span4Mux_s3_v
    port map (
            O => \N__7298\,
            I => \N__7295\
        );

    \I__1420\ : Span4Mux_h
    port map (
            O => \N__7295\,
            I => \N__7292\
        );

    \I__1419\ : Span4Mux_v
    port map (
            O => \N__7292\,
            I => \N__7289\
        );

    \I__1418\ : Span4Mux_v
    port map (
            O => \N__7289\,
            I => \N__7286\
        );

    \I__1417\ : Span4Mux_v
    port map (
            O => \N__7286\,
            I => \N__7282\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7285\,
            I => \N__7279\
        );

    \I__1415\ : Odrv4
    port map (
            O => \N__7282\,
            I => \ROMENn_c\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__7279\,
            I => \ROMENn_c\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7274\,
            I => \N__7271\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__7271\,
            I => \N__7267\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7270\,
            I => \N__7264\
        );

    \I__1410\ : Span4Mux_h
    port map (
            O => \N__7267\,
            I => \N__7259\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__7264\,
            I => \N__7259\
        );

    \I__1408\ : Odrv4
    port map (
            O => \N__7259\,
            I => \U409_TRANSFER_ACK.un1_AUTOVECTOR_0\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7256\,
            I => \N__7253\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7253\,
            I => \N__7249\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7252\,
            I => \N__7246\
        );

    \I__1404\ : Span4Mux_v
    port map (
            O => \N__7249\,
            I => \N__7240\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7246\,
            I => \N__7240\
        );

    \I__1402\ : InMux
    port map (
            O => \N__7245\,
            I => \N__7237\
        );

    \I__1401\ : Span4Mux_h
    port map (
            O => \N__7240\,
            I => \N__7229\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7237\,
            I => \N__7229\
        );

    \I__1399\ : InMux
    port map (
            O => \N__7236\,
            I => \N__7226\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7235\,
            I => \N__7223\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7234\,
            I => \N__7220\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__7229\,
            I => \N__7217\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7226\,
            I => \N__7214\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__7223\,
            I => \N__7211\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7220\,
            I => \N__7208\
        );

    \I__1392\ : Span4Mux_v
    port map (
            O => \N__7217\,
            I => \N__7203\
        );

    \I__1391\ : Span4Mux_v
    port map (
            O => \N__7214\,
            I => \N__7203\
        );

    \I__1390\ : Span4Mux_v
    port map (
            O => \N__7211\,
            I => \N__7200\
        );

    \I__1389\ : Span12Mux_h
    port map (
            O => \N__7208\,
            I => \N__7197\
        );

    \I__1388\ : Sp12to4
    port map (
            O => \N__7203\,
            I => \N__7192\
        );

    \I__1387\ : Sp12to4
    port map (
            O => \N__7200\,
            I => \N__7192\
        );

    \I__1386\ : Span12Mux_v
    port map (
            O => \N__7197\,
            I => \N__7189\
        );

    \I__1385\ : Span12Mux_h
    port map (
            O => \N__7192\,
            I => \N__7186\
        );

    \I__1384\ : Odrv12
    port map (
            O => \N__7189\,
            I => \TSn_c\
        );

    \I__1383\ : Odrv12
    port map (
            O => \N__7186\,
            I => \TSn_c\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7181\,
            I => \N__7178\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__7178\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1\
        );

    \I__1380\ : InMux
    port map (
            O => \N__7175\,
            I => \N__7169\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7174\,
            I => \N__7169\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__7169\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__1377\ : InMux
    port map (
            O => \N__7166\,
            I => \N__7162\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7165\,
            I => \N__7159\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__7162\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7159\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__7154\,
            I => \U409_TRANSFER_ACK.N_17_mux_cascade_\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__7151\,
            I => \U409_TRANSFER_ACK.N_3_0_cascade_\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__7148\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0_cascade_\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7142\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__7142\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7136\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7136\,
            I => \U409_TRANSFER_ACK.N_3_0\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__7133\,
            I => \U409_TRANSFER_ACK.N_6_0_cascade_\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7126\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7129\,
            I => \N__7123\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__7126\,
            I => \ATA_BASE_2\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__7123\,
            I => \ATA_BASE_2\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__7118\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2_cascade_\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7115\,
            I => \N__7111\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7114\,
            I => \N__7108\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__7111\,
            I => \N__7105\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7108\,
            I => \ATA_BASE_7\
        );

    \I__1356\ : Odrv4
    port map (
            O => \N__7105\,
            I => \ATA_BASE_7\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7097\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7097\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7094\,
            I => \N__7091\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__7091\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_0\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__7088\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_5_cascade_\
        );

    \I__1350\ : CascadeMux
    port map (
            O => \N__7085\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7082\,
            I => \N__7078\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7081\,
            I => \N__7075\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__7078\,
            I => \U409_AUTOCONFIG.un1_STATE_6_0\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7075\,
            I => \U409_AUTOCONFIG.un1_STATE_6_0\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7057\
        );

    \I__1344\ : InMux
    port map (
            O => \N__7069\,
            I => \N__7054\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7068\,
            I => \N__7051\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7067\,
            I => \N__7046\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7066\,
            I => \N__7046\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7065\,
            I => \N__7039\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7064\,
            I => \N__7039\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7063\,
            I => \N__7039\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7062\,
            I => \N__7036\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__7061\,
            I => \N__7033\
        );

    \I__1335\ : InMux
    port map (
            O => \N__7060\,
            I => \N__7028\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7057\,
            I => \N__7025\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__7054\,
            I => \N__7017\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__7051\,
            I => \N__7017\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__7046\,
            I => \N__7017\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__7039\,
            I => \N__7011\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__7036\,
            I => \N__7011\
        );

    \I__1328\ : InMux
    port map (
            O => \N__7033\,
            I => \N__7004\
        );

    \I__1327\ : InMux
    port map (
            O => \N__7032\,
            I => \N__7004\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7004\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__7028\,
            I => \N__7001\
        );

    \I__1324\ : Span4Mux_v
    port map (
            O => \N__7025\,
            I => \N__6998\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7024\,
            I => \N__6995\
        );

    \I__1322\ : Span4Mux_v
    port map (
            O => \N__7017\,
            I => \N__6992\
        );

    \I__1321\ : InMux
    port map (
            O => \N__7016\,
            I => \N__6989\
        );

    \I__1320\ : Span4Mux_h
    port map (
            O => \N__7011\,
            I => \N__6984\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__7004\,
            I => \N__6984\
        );

    \I__1318\ : Sp12to4
    port map (
            O => \N__7001\,
            I => \N__6981\
        );

    \I__1317\ : Sp12to4
    port map (
            O => \N__6998\,
            I => \N__6972\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6995\,
            I => \N__6972\
        );

    \I__1315\ : Sp12to4
    port map (
            O => \N__6992\,
            I => \N__6972\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__6989\,
            I => \N__6972\
        );

    \I__1313\ : Span4Mux_v
    port map (
            O => \N__6984\,
            I => \N__6969\
        );

    \I__1312\ : Span12Mux_v
    port map (
            O => \N__6981\,
            I => \N__6966\
        );

    \I__1311\ : Span12Mux_h
    port map (
            O => \N__6972\,
            I => \N__6963\
        );

    \I__1310\ : Span4Mux_h
    port map (
            O => \N__6969\,
            I => \N__6960\
        );

    \I__1309\ : Span12Mux_h
    port map (
            O => \N__6966\,
            I => \N__6955\
        );

    \I__1308\ : Span12Mux_v
    port map (
            O => \N__6963\,
            I => \N__6955\
        );

    \I__1307\ : Sp12to4
    port map (
            O => \N__6960\,
            I => \N__6952\
        );

    \I__1306\ : Odrv12
    port map (
            O => \N__6955\,
            I => \A_c_1\
        );

    \I__1305\ : Odrv12
    port map (
            O => \N__6952\,
            I => \A_c_1\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6947\,
            I => \N__6944\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6944\,
            I => \N__6940\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6943\,
            I => \N__6937\
        );

    \I__1301\ : Span4Mux_v
    port map (
            O => \N__6940\,
            I => \N__6933\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6937\,
            I => \N__6930\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6936\,
            I => \N__6927\
        );

    \I__1298\ : Span4Mux_h
    port map (
            O => \N__6933\,
            I => \N__6919\
        );

    \I__1297\ : Span4Mux_v
    port map (
            O => \N__6930\,
            I => \N__6919\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__6927\,
            I => \N__6919\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6926\,
            I => \N__6916\
        );

    \I__1294\ : Span4Mux_v
    port map (
            O => \N__6919\,
            I => \N__6912\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6916\,
            I => \N__6909\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6915\,
            I => \N__6906\
        );

    \I__1291\ : Span4Mux_v
    port map (
            O => \N__6912\,
            I => \N__6903\
        );

    \I__1290\ : Span4Mux_v
    port map (
            O => \N__6909\,
            I => \N__6898\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6906\,
            I => \N__6898\
        );

    \I__1288\ : Span4Mux_v
    port map (
            O => \N__6903\,
            I => \N__6895\
        );

    \I__1287\ : Sp12to4
    port map (
            O => \N__6898\,
            I => \N__6892\
        );

    \I__1286\ : Sp12to4
    port map (
            O => \N__6895\,
            I => \N__6887\
        );

    \I__1285\ : Span12Mux_v
    port map (
            O => \N__6892\,
            I => \N__6887\
        );

    \I__1284\ : Odrv12
    port map (
            O => \N__6887\,
            I => \A_c_17\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6884\,
            I => \N__6881\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__6881\,
            I => \U409_ADDRESS_DECODE.un2_ATA_SPACEZ0Z_0\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6878\,
            I => \N__6875\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__6875\,
            I => \N__6871\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6874\,
            I => \N__6868\
        );

    \I__1278\ : Odrv12
    port map (
            O => \N__6871\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6868\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__6863\,
            I => \U409_ADDRESS_DECODE_PORTSIZE_0_cascade_\
        );

    \I__1275\ : IoInMux
    port map (
            O => \N__6860\,
            I => \N__6857\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__6857\,
            I => \N__6854\
        );

    \I__1273\ : Span4Mux_s3_v
    port map (
            O => \N__6854\,
            I => \N__6851\
        );

    \I__1272\ : Span4Mux_h
    port map (
            O => \N__6851\,
            I => \N__6848\
        );

    \I__1271\ : Sp12to4
    port map (
            O => \N__6848\,
            I => \N__6845\
        );

    \I__1270\ : Span12Mux_v
    port map (
            O => \N__6845\,
            I => \N__6842\
        );

    \I__1269\ : Odrv12
    port map (
            O => \N__6842\,
            I => \PORTSIZE_0_i\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__6839\,
            I => \N__6835\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6838\,
            I => \N__6832\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6829\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6832\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6829\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__6824\,
            I => \N__6819\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__6823\,
            I => \N__6815\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__6822\,
            I => \N__6812\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6819\,
            I => \N__6806\
        );

    \I__1259\ : InMux
    port map (
            O => \N__6818\,
            I => \N__6806\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6815\,
            I => \N__6799\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6812\,
            I => \N__6799\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6811\,
            I => \N__6799\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__6806\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6799\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__6794\,
            I => \N__6791\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6785\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6790\,
            I => \N__6780\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6789\,
            I => \N__6780\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6777\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6785\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6780\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6777\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__6770\,
            I => \N__6762\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6755\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6755\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6767\,
            I => \N__6755\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6766\,
            I => \N__6752\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6747\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6762\,
            I => \N__6747\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6755\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6752\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6747\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6740\,
            I => \N__6735\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6739\,
            I => \N__6730\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6738\,
            I => \N__6730\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6735\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__6730\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6725\,
            I => \N__6722\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__6722\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_2\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6715\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6718\,
            I => \N__6710\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6715\,
            I => \N__6707\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6714\,
            I => \N__6702\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6713\,
            I => \N__6702\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6710\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__6707\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__6702\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6695\,
            I => \N__6692\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6692\,
            I => \N__6689\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__6689\,
            I => \U409_AUTOCONFIG.STATE_d_2\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6686\,
            I => \N__6683\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__6683\,
            I => \N__6678\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6682\,
            I => \N__6675\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6681\,
            I => \N__6672\
        );

    \I__1213\ : Span4Mux_v
    port map (
            O => \N__6678\,
            I => \N__6669\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6675\,
            I => \N__6664\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6672\,
            I => \N__6664\
        );

    \I__1210\ : Sp12to4
    port map (
            O => \N__6669\,
            I => \N__6661\
        );

    \I__1209\ : Span4Mux_v
    port map (
            O => \N__6664\,
            I => \N__6658\
        );

    \I__1208\ : Odrv12
    port map (
            O => \N__6661\,
            I => \U409_AUTOCONFIG.un1_AZ0Z_16\
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__6658\,
            I => \U409_AUTOCONFIG.un1_AZ0Z_16\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6647\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6652\,
            I => \N__6643\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6638\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6650\,
            I => \N__6638\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__6647\,
            I => \N__6635\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6646\,
            I => \N__6632\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6643\,
            I => \N__6625\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6638\,
            I => \N__6625\
        );

    \I__1198\ : Span4Mux_v
    port map (
            O => \N__6635\,
            I => \N__6620\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6632\,
            I => \N__6620\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6631\,
            I => \N__6617\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6630\,
            I => \N__6613\
        );

    \I__1194\ : Span4Mux_v
    port map (
            O => \N__6625\,
            I => \N__6606\
        );

    \I__1193\ : Span4Mux_v
    port map (
            O => \N__6620\,
            I => \N__6606\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6617\,
            I => \N__6606\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6616\,
            I => \N__6603\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__6613\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1189\ : Odrv4
    port map (
            O => \N__6606\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6603\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__6596\,
            I => \N__6593\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6593\,
            I => \N__6589\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6592\,
            I => \N__6586\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6589\,
            I => \N__6581\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6586\,
            I => \N__6581\
        );

    \I__1182\ : Span4Mux_v
    port map (
            O => \N__6581\,
            I => \N__6578\
        );

    \I__1181\ : Sp12to4
    port map (
            O => \N__6578\,
            I => \N__6575\
        );

    \I__1180\ : Span12Mux_h
    port map (
            O => \N__6575\,
            I => \N__6572\
        );

    \I__1179\ : Span12Mux_v
    port map (
            O => \N__6572\,
            I => \N__6569\
        );

    \I__1178\ : Odrv12
    port map (
            O => \N__6569\,
            I => \D_in_4\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6566\,
            I => \N__6563\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__6563\,
            I => \N__6560\
        );

    \I__1175\ : Span4Mux_v
    port map (
            O => \N__6560\,
            I => \N__6556\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6559\,
            I => \N__6553\
        );

    \I__1173\ : Odrv4
    port map (
            O => \N__6556\,
            I => \BRIDGE_BASE_0\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6553\,
            I => \BRIDGE_BASE_0\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6548\,
            I => \N__6536\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6536\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6546\,
            I => \N__6536\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6545\,
            I => \N__6533\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6544\,
            I => \N__6530\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6543\,
            I => \N__6527\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6536\,
            I => \N__6524\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__6533\,
            I => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6530\,
            I => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__6527\,
            I => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\
        );

    \I__1161\ : Odrv12
    port map (
            O => \N__6524\,
            I => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6515\,
            I => \N__6512\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6512\,
            I => \N__6509\
        );

    \I__1158\ : Span4Mux_v
    port map (
            O => \N__6509\,
            I => \N__6505\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6508\,
            I => \N__6502\
        );

    \I__1156\ : Odrv4
    port map (
            O => \N__6505\,
            I => \BRIDGE_BASE_1\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6502\,
            I => \BRIDGE_BASE_1\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6497\,
            I => \N__6493\
        );

    \I__1153\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6488\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6493\,
            I => \N__6485\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6482\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6479\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6488\,
            I => \N__6472\
        );

    \I__1148\ : Span4Mux_h
    port map (
            O => \N__6485\,
            I => \N__6467\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6482\,
            I => \N__6467\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6479\,
            I => \N__6464\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6459\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6477\,
            I => \N__6459\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6476\,
            I => \N__6456\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6453\
        );

    \I__1141\ : Span4Mux_h
    port map (
            O => \N__6472\,
            I => \N__6448\
        );

    \I__1140\ : Span4Mux_v
    port map (
            O => \N__6467\,
            I => \N__6448\
        );

    \I__1139\ : Span4Mux_v
    port map (
            O => \N__6464\,
            I => \N__6445\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__6459\,
            I => \N__6442\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6456\,
            I => \N__6437\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6453\,
            I => \N__6437\
        );

    \I__1135\ : Span4Mux_h
    port map (
            O => \N__6448\,
            I => \N__6434\
        );

    \I__1134\ : Span4Mux_v
    port map (
            O => \N__6445\,
            I => \N__6431\
        );

    \I__1133\ : Span4Mux_v
    port map (
            O => \N__6442\,
            I => \N__6428\
        );

    \I__1132\ : Span4Mux_v
    port map (
            O => \N__6437\,
            I => \N__6425\
        );

    \I__1131\ : Span4Mux_v
    port map (
            O => \N__6434\,
            I => \N__6422\
        );

    \I__1130\ : Sp12to4
    port map (
            O => \N__6431\,
            I => \N__6415\
        );

    \I__1129\ : Sp12to4
    port map (
            O => \N__6428\,
            I => \N__6415\
        );

    \I__1128\ : Sp12to4
    port map (
            O => \N__6425\,
            I => \N__6415\
        );

    \I__1127\ : Sp12to4
    port map (
            O => \N__6422\,
            I => \N__6410\
        );

    \I__1126\ : Span12Mux_h
    port map (
            O => \N__6415\,
            I => \N__6410\
        );

    \I__1125\ : Span12Mux_v
    port map (
            O => \N__6410\,
            I => \N__6407\
        );

    \I__1124\ : Odrv12
    port map (
            O => \N__6407\,
            I => \A_c_19\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__6404\,
            I => \N__6399\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6403\,
            I => \N__6395\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__6402\,
            I => \N__6392\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6399\,
            I => \N__6388\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6398\,
            I => \N__6385\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6395\,
            I => \N__6382\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6392\,
            I => \N__6379\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6391\,
            I => \N__6376\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__6388\,
            I => \N__6373\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6385\,
            I => \N__6370\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__6382\,
            I => \N__6363\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6379\,
            I => \N__6363\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__6376\,
            I => \N__6363\
        );

    \I__1110\ : Span4Mux_v
    port map (
            O => \N__6373\,
            I => \N__6359\
        );

    \I__1109\ : Span4Mux_v
    port map (
            O => \N__6370\,
            I => \N__6354\
        );

    \I__1108\ : Span4Mux_v
    port map (
            O => \N__6363\,
            I => \N__6354\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6362\,
            I => \N__6351\
        );

    \I__1106\ : Sp12to4
    port map (
            O => \N__6359\,
            I => \N__6344\
        );

    \I__1105\ : Sp12to4
    port map (
            O => \N__6354\,
            I => \N__6344\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6351\,
            I => \N__6344\
        );

    \I__1103\ : Span12Mux_h
    port map (
            O => \N__6344\,
            I => \N__6341\
        );

    \I__1102\ : Span12Mux_v
    port map (
            O => \N__6341\,
            I => \N__6338\
        );

    \I__1101\ : Odrv12
    port map (
            O => \N__6338\,
            I => \A_c_18\
        );

    \I__1100\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6332\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6332\,
            I => \N__6329\
        );

    \I__1098\ : Odrv12
    port map (
            O => \N__6329\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6323\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__6323\,
            I => \N__6320\
        );

    \I__1095\ : Odrv4
    port map (
            O => \N__6320\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_11_0\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6317\,
            I => \N__6310\
        );

    \I__1093\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6303\
        );

    \I__1092\ : InMux
    port map (
            O => \N__6315\,
            I => \N__6303\
        );

    \I__1091\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6303\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6300\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__6310\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__6303\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__6300\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6287\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6292\,
            I => \N__6282\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6282\
        );

    \I__1083\ : InMux
    port map (
            O => \N__6290\,
            I => \N__6279\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__6287\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__6282\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__6279\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1079\ : CascadeMux
    port map (
            O => \N__6272\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_5_cascade_\
        );

    \I__1078\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6266\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__6266\,
            I => \N__6263\
        );

    \I__1076\ : Span4Mux_v
    port map (
            O => \N__6263\,
            I => \N__6259\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6262\,
            I => \N__6256\
        );

    \I__1074\ : Odrv4
    port map (
            O => \N__6259\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__6256\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__6251\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_cascade_\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__6248\,
            I => \N__6245\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6245\,
            I => \N__6242\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6242\,
            I => \N__6238\
        );

    \I__1068\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6235\
        );

    \I__1067\ : Odrv12
    port map (
            O => \N__6238\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6235\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6230\,
            I => \N__6227\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__6227\,
            I => \N__6218\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6226\,
            I => \N__6213\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6213\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6224\,
            I => \N__6208\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6223\,
            I => \N__6208\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6222\,
            I => \N__6205\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6221\,
            I => \N__6202\
        );

    \I__1057\ : Span4Mux_v
    port map (
            O => \N__6218\,
            I => \N__6199\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6213\,
            I => \N__6196\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__6208\,
            I => \N__6189\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__6205\,
            I => \N__6189\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__6202\,
            I => \N__6189\
        );

    \I__1052\ : Span4Mux_h
    port map (
            O => \N__6199\,
            I => \N__6184\
        );

    \I__1051\ : Span4Mux_v
    port map (
            O => \N__6196\,
            I => \N__6184\
        );

    \I__1050\ : Span12Mux_v
    port map (
            O => \N__6189\,
            I => \N__6179\
        );

    \I__1049\ : Sp12to4
    port map (
            O => \N__6184\,
            I => \N__6179\
        );

    \I__1048\ : Odrv12
    port map (
            O => \N__6179\,
            I => \A_c_7\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6176\,
            I => \N__6173\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6173\,
            I => \N__6170\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__6170\,
            I => \U409_AUTOCONFIG.ATA_BASE11Z0Z_1\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__6167\,
            I => \N__6162\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6166\,
            I => \N__6153\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6165\,
            I => \N__6153\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6162\,
            I => \N__6150\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6145\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6160\,
            I => \N__6140\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6159\,
            I => \N__6140\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6137\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6153\,
            I => \N__6134\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6150\,
            I => \N__6131\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6149\,
            I => \N__6128\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__6148\,
            I => \N__6125\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6145\,
            I => \N__6121\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6140\,
            I => \N__6115\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6137\,
            I => \N__6115\
        );

    \I__1029\ : Span4Mux_v
    port map (
            O => \N__6134\,
            I => \N__6112\
        );

    \I__1028\ : Span4Mux_h
    port map (
            O => \N__6131\,
            I => \N__6107\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__6128\,
            I => \N__6107\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6125\,
            I => \N__6102\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6124\,
            I => \N__6102\
        );

    \I__1024\ : Span4Mux_v
    port map (
            O => \N__6121\,
            I => \N__6099\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6120\,
            I => \N__6096\
        );

    \I__1022\ : Span12Mux_v
    port map (
            O => \N__6115\,
            I => \N__6083\
        );

    \I__1021\ : Sp12to4
    port map (
            O => \N__6112\,
            I => \N__6083\
        );

    \I__1020\ : Sp12to4
    port map (
            O => \N__6107\,
            I => \N__6083\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6102\,
            I => \N__6083\
        );

    \I__1018\ : Sp12to4
    port map (
            O => \N__6099\,
            I => \N__6083\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__6096\,
            I => \N__6083\
        );

    \I__1016\ : Odrv12
    port map (
            O => \N__6083\,
            I => \A_c_5\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6080\,
            I => \N__6071\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6079\,
            I => \N__6068\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6063\
        );

    \I__1012\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6063\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6060\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6075\,
            I => \N__6057\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6074\,
            I => \N__6054\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6071\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6068\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6063\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__6060\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6057\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6054\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1002\ : CascadeMux
    port map (
            O => \N__6041\,
            I => \U409_AUTOCONFIG.ATA_BASE11_cascade_\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6034\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__6037\,
            I => \N__6028\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__6034\,
            I => \N__6023\
        );

    \I__998\ : InMux
    port map (
            O => \N__6033\,
            I => \N__6020\
        );

    \I__997\ : InMux
    port map (
            O => \N__6032\,
            I => \N__6017\
        );

    \I__996\ : InMux
    port map (
            O => \N__6031\,
            I => \N__6012\
        );

    \I__995\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6012\
        );

    \I__994\ : InMux
    port map (
            O => \N__6027\,
            I => \N__6009\
        );

    \I__993\ : InMux
    port map (
            O => \N__6026\,
            I => \N__6006\
        );

    \I__992\ : Span4Mux_v
    port map (
            O => \N__6023\,
            I => \N__6001\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__6020\,
            I => \N__6001\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__6017\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__6012\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__6009\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__6006\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__6001\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__985\ : InMux
    port map (
            O => \N__5990\,
            I => \N__5986\
        );

    \I__984\ : CascadeMux
    port map (
            O => \N__5989\,
            I => \N__5983\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5986\,
            I => \N__5976\
        );

    \I__982\ : InMux
    port map (
            O => \N__5983\,
            I => \N__5973\
        );

    \I__981\ : InMux
    port map (
            O => \N__5982\,
            I => \N__5963\
        );

    \I__980\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5963\
        );

    \I__979\ : InMux
    port map (
            O => \N__5980\,
            I => \N__5963\
        );

    \I__978\ : InMux
    port map (
            O => \N__5979\,
            I => \N__5963\
        );

    \I__977\ : Span4Mux_v
    port map (
            O => \N__5976\,
            I => \N__5960\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5973\,
            I => \N__5957\
        );

    \I__975\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5954\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__5963\,
            I => \N__5951\
        );

    \I__973\ : Odrv4
    port map (
            O => \N__5960\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\
        );

    \I__972\ : Odrv4
    port map (
            O => \N__5957\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__5954\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\
        );

    \I__970\ : Odrv4
    port map (
            O => \N__5951\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\
        );

    \I__969\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5936\
        );

    \I__968\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5933\
        );

    \I__967\ : InMux
    port map (
            O => \N__5940\,
            I => \N__5930\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__5939\,
            I => \N__5927\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__5936\,
            I => \N__5921\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5933\,
            I => \N__5916\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__5930\,
            I => \N__5916\
        );

    \I__962\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5909\
        );

    \I__961\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5909\
        );

    \I__960\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5909\
        );

    \I__959\ : InMux
    port map (
            O => \N__5924\,
            I => \N__5906\
        );

    \I__958\ : Span4Mux_v
    port map (
            O => \N__5921\,
            I => \N__5903\
        );

    \I__957\ : Span4Mux_v
    port map (
            O => \N__5916\,
            I => \N__5900\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__5909\,
            I => \N__5895\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5906\,
            I => \N__5895\
        );

    \I__954\ : Odrv4
    port map (
            O => \N__5903\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_6\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__5900\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_6\
        );

    \I__952\ : Odrv4
    port map (
            O => \N__5895\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_6\
        );

    \I__951\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5882\
        );

    \I__950\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5882\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5882\,
            I => \ATA_BASE_6\
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__5879\,
            I => \N__5874\
        );

    \I__947\ : InMux
    port map (
            O => \N__5878\,
            I => \N__5869\
        );

    \I__946\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5869\
        );

    \I__945\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5866\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5869\,
            I => \N__5861\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__5866\,
            I => \N__5861\
        );

    \I__942\ : Span4Mux_v
    port map (
            O => \N__5861\,
            I => \N__5858\
        );

    \I__941\ : Sp12to4
    port map (
            O => \N__5858\,
            I => \N__5855\
        );

    \I__940\ : Span12Mux_h
    port map (
            O => \N__5855\,
            I => \N__5852\
        );

    \I__939\ : Span12Mux_v
    port map (
            O => \N__5852\,
            I => \N__5849\
        );

    \I__938\ : Odrv12
    port map (
            O => \N__5849\,
            I => \D_in_6\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__5846\,
            I => \N__5842\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__5845\,
            I => \N__5839\
        );

    \I__935\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5836\
        );

    \I__934\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5833\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__5836\,
            I => \N__5830\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__5833\,
            I => \BRIDGE_BASE_2\
        );

    \I__931\ : Odrv4
    port map (
            O => \N__5830\,
            I => \BRIDGE_BASE_2\
        );

    \I__930\ : InMux
    port map (
            O => \N__5825\,
            I => \N__5819\
        );

    \I__929\ : InMux
    port map (
            O => \N__5824\,
            I => \N__5819\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5819\,
            I => \N__5814\
        );

    \I__927\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5811\
        );

    \I__926\ : CascadeMux
    port map (
            O => \N__5817\,
            I => \N__5805\
        );

    \I__925\ : Span4Mux_h
    port map (
            O => \N__5814\,
            I => \N__5800\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5811\,
            I => \N__5800\
        );

    \I__923\ : InMux
    port map (
            O => \N__5810\,
            I => \N__5797\
        );

    \I__922\ : InMux
    port map (
            O => \N__5809\,
            I => \N__5792\
        );

    \I__921\ : InMux
    port map (
            O => \N__5808\,
            I => \N__5792\
        );

    \I__920\ : InMux
    port map (
            O => \N__5805\,
            I => \N__5787\
        );

    \I__919\ : Span4Mux_h
    port map (
            O => \N__5800\,
            I => \N__5782\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5797\,
            I => \N__5782\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__5792\,
            I => \N__5779\
        );

    \I__916\ : InMux
    port map (
            O => \N__5791\,
            I => \N__5776\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__5790\,
            I => \N__5773\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__5787\,
            I => \N__5770\
        );

    \I__913\ : Span4Mux_v
    port map (
            O => \N__5782\,
            I => \N__5765\
        );

    \I__912\ : Span4Mux_v
    port map (
            O => \N__5779\,
            I => \N__5765\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__5776\,
            I => \N__5762\
        );

    \I__910\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5759\
        );

    \I__909\ : Span12Mux_h
    port map (
            O => \N__5770\,
            I => \N__5750\
        );

    \I__908\ : Sp12to4
    port map (
            O => \N__5765\,
            I => \N__5750\
        );

    \I__907\ : Span12Mux_v
    port map (
            O => \N__5762\,
            I => \N__5750\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5759\,
            I => \N__5750\
        );

    \I__905\ : Odrv12
    port map (
            O => \N__5750\,
            I => \A_c_20\
        );

    \I__904\ : InMux
    port map (
            O => \N__5747\,
            I => \N__5741\
        );

    \I__903\ : InMux
    port map (
            O => \N__5746\,
            I => \N__5741\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5741\,
            I => \ATA_BASE_4\
        );

    \I__901\ : InMux
    port map (
            O => \N__5738\,
            I => \N__5732\
        );

    \I__900\ : InMux
    port map (
            O => \N__5737\,
            I => \N__5725\
        );

    \I__899\ : InMux
    port map (
            O => \N__5736\,
            I => \N__5725\
        );

    \I__898\ : InMux
    port map (
            O => \N__5735\,
            I => \N__5725\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5732\,
            I => \U409_AUTOCONFIG.LIDE_CONF_RNIDFPAZ0Z3\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5725\,
            I => \U409_AUTOCONFIG.LIDE_CONF_RNIDFPAZ0Z3\
        );

    \I__895\ : InMux
    port map (
            O => \N__5720\,
            I => \N__5714\
        );

    \I__894\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5714\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5714\,
            I => \ATA_BASE_5\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__5711\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__5708\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__890\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5698\
        );

    \I__889\ : InMux
    port map (
            O => \N__5704\,
            I => \N__5698\
        );

    \I__888\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5695\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5698\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5695\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__5690\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_\
        );

    \I__884\ : InMux
    port map (
            O => \N__5687\,
            I => \N__5684\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__5684\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5\
        );

    \I__882\ : IoInMux
    port map (
            O => \N__5681\,
            I => \N__5678\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5678\,
            I => \N__5675\
        );

    \I__880\ : Span12Mux_s8_v
    port map (
            O => \N__5675\,
            I => \N__5672\
        );

    \I__879\ : Span12Mux_h
    port map (
            O => \N__5672\,
            I => \N__5668\
        );

    \I__878\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5665\
        );

    \I__877\ : Odrv12
    port map (
            O => \N__5668\,
            I => \CONFIGENn_c\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5665\,
            I => \CONFIGENn_c\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__5660\,
            I => \U409_AUTOCONFIG.STATE_d_2_cascade_\
        );

    \I__874\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5653\
        );

    \I__873\ : InMux
    port map (
            O => \N__5656\,
            I => \N__5650\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5653\,
            I => \N__5646\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5650\,
            I => \N__5643\
        );

    \I__870\ : InMux
    port map (
            O => \N__5649\,
            I => \N__5640\
        );

    \I__869\ : Span4Mux_v
    port map (
            O => \N__5646\,
            I => \N__5637\
        );

    \I__868\ : Span4Mux_v
    port map (
            O => \N__5643\,
            I => \N__5634\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5640\,
            I => \N__5631\
        );

    \I__866\ : Span4Mux_v
    port map (
            O => \N__5637\,
            I => \N__5628\
        );

    \I__865\ : Span4Mux_v
    port map (
            O => \N__5634\,
            I => \N__5625\
        );

    \I__864\ : Span12Mux_v
    port map (
            O => \N__5631\,
            I => \N__5618\
        );

    \I__863\ : Sp12to4
    port map (
            O => \N__5628\,
            I => \N__5618\
        );

    \I__862\ : Sp12to4
    port map (
            O => \N__5625\,
            I => \N__5618\
        );

    \I__861\ : Odrv12
    port map (
            O => \N__5618\,
            I => \A_c_31\
        );

    \I__860\ : InMux
    port map (
            O => \N__5615\,
            I => \N__5611\
        );

    \I__859\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5608\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5611\,
            I => \N__5605\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__5608\,
            I => \N__5602\
        );

    \I__856\ : Span4Mux_v
    port map (
            O => \N__5605\,
            I => \N__5598\
        );

    \I__855\ : Span4Mux_v
    port map (
            O => \N__5602\,
            I => \N__5595\
        );

    \I__854\ : InMux
    port map (
            O => \N__5601\,
            I => \N__5592\
        );

    \I__853\ : Span4Mux_v
    port map (
            O => \N__5598\,
            I => \N__5589\
        );

    \I__852\ : Span4Mux_v
    port map (
            O => \N__5595\,
            I => \N__5586\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5592\,
            I => \N__5583\
        );

    \I__850\ : Span4Mux_h
    port map (
            O => \N__5589\,
            I => \N__5580\
        );

    \I__849\ : Span4Mux_h
    port map (
            O => \N__5586\,
            I => \N__5577\
        );

    \I__848\ : Sp12to4
    port map (
            O => \N__5583\,
            I => \N__5574\
        );

    \I__847\ : Sp12to4
    port map (
            O => \N__5580\,
            I => \N__5567\
        );

    \I__846\ : Sp12to4
    port map (
            O => \N__5577\,
            I => \N__5567\
        );

    \I__845\ : Span12Mux_v
    port map (
            O => \N__5574\,
            I => \N__5567\
        );

    \I__844\ : Odrv12
    port map (
            O => \N__5567\,
            I => \A_c_30\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__5564\,
            I => \N__5560\
        );

    \I__842\ : InMux
    port map (
            O => \N__5563\,
            I => \N__5557\
        );

    \I__841\ : InMux
    port map (
            O => \N__5560\,
            I => \N__5554\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5557\,
            I => \BRIDGE_BASE_3\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5554\,
            I => \BRIDGE_BASE_3\
        );

    \I__838\ : InMux
    port map (
            O => \N__5549\,
            I => \N__5546\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5546\,
            I => \N__5541\
        );

    \I__836\ : InMux
    port map (
            O => \N__5545\,
            I => \N__5538\
        );

    \I__835\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5535\
        );

    \I__834\ : Span4Mux_h
    port map (
            O => \N__5541\,
            I => \N__5530\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__5538\,
            I => \N__5530\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5535\,
            I => \N__5525\
        );

    \I__831\ : Sp12to4
    port map (
            O => \N__5530\,
            I => \N__5525\
        );

    \I__830\ : Span12Mux_v
    port map (
            O => \N__5525\,
            I => \N__5522\
        );

    \I__829\ : Odrv12
    port map (
            O => \N__5522\,
            I => \A_c_29\
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__5519\,
            I => \N__5515\
        );

    \I__827\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5511\
        );

    \I__826\ : InMux
    port map (
            O => \N__5515\,
            I => \N__5508\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__5514\,
            I => \N__5505\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5511\,
            I => \N__5500\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__5508\,
            I => \N__5500\
        );

    \I__822\ : InMux
    port map (
            O => \N__5505\,
            I => \N__5497\
        );

    \I__821\ : Span4Mux_h
    port map (
            O => \N__5500\,
            I => \N__5494\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5497\,
            I => \N__5491\
        );

    \I__819\ : Sp12to4
    port map (
            O => \N__5494\,
            I => \N__5488\
        );

    \I__818\ : Span12Mux_v
    port map (
            O => \N__5491\,
            I => \N__5485\
        );

    \I__817\ : Span12Mux_v
    port map (
            O => \N__5488\,
            I => \N__5482\
        );

    \I__816\ : Odrv12
    port map (
            O => \N__5485\,
            I => \A_c_28\
        );

    \I__815\ : Odrv12
    port map (
            O => \N__5482\,
            I => \A_c_28\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__5477\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2Z0Z_0_cascade_\
        );

    \I__813\ : InMux
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5471\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_3\
        );

    \I__811\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5465\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__5465\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0\
        );

    \I__809\ : InMux
    port map (
            O => \N__5462\,
            I => \N__5458\
        );

    \I__808\ : InMux
    port map (
            O => \N__5461\,
            I => \N__5455\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__5458\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_4\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5455\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_4\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__5450\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_\
        );

    \I__804\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5444\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5444\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_2_0\
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__5441\,
            I => \N__5438\
        );

    \I__801\ : InMux
    port map (
            O => \N__5438\,
            I => \N__5434\
        );

    \I__800\ : InMux
    port map (
            O => \N__5437\,
            I => \N__5431\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__5434\,
            I => \N__5426\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5431\,
            I => \N__5426\
        );

    \I__797\ : Span4Mux_v
    port map (
            O => \N__5426\,
            I => \N__5423\
        );

    \I__796\ : Odrv4
    port map (
            O => \N__5423\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6\
        );

    \I__795\ : InMux
    port map (
            O => \N__5420\,
            I => \N__5417\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__5417\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7\
        );

    \I__793\ : InMux
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5411\,
            I => \U409_ADDRESS_DECODE_AUTOVECTOR_8\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__5408\,
            I => \U409_ADDRESS_DECODE_AUTOVECTOR_10_cascade_\
        );

    \I__790\ : InMux
    port map (
            O => \N__5405\,
            I => \N__5402\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5402\,
            I => \U409_ADDRESS_DECODE_AUTOVECTOR_9\
        );

    \I__788\ : InMux
    port map (
            O => \N__5399\,
            I => \N__5396\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5396\,
            I => \N__5392\
        );

    \I__786\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5389\
        );

    \I__785\ : Odrv4
    port map (
            O => \N__5392\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__5389\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__5384\,
            I => \N__5381\
        );

    \I__782\ : InMux
    port map (
            O => \N__5381\,
            I => \N__5377\
        );

    \I__781\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5374\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5377\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5374\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\
        );

    \I__778\ : IoInMux
    port map (
            O => \N__5369\,
            I => \N__5366\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__776\ : Span12Mux_s6_v
    port map (
            O => \N__5363\,
            I => \N__5360\
        );

    \I__775\ : Odrv12
    port map (
            O => \N__5360\,
            I => \U409_AUTOCONFIG_D_OUT_0_i_1\
        );

    \I__774\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5353\
        );

    \I__773\ : InMux
    port map (
            O => \N__5356\,
            I => \N__5350\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5353\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5350\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\
        );

    \I__770\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5342\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5342\,
            I => \N__5338\
        );

    \I__768\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5335\
        );

    \I__767\ : Odrv4
    port map (
            O => \N__5338\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5335\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2\
        );

    \I__765\ : IoInMux
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5327\,
            I => \N__5324\
        );

    \I__763\ : Span12Mux_s7_v
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__762\ : Odrv12
    port map (
            O => \N__5321\,
            I => \U409_AUTOCONFIG_D_OUT_0_i_2\
        );

    \I__761\ : InMux
    port map (
            O => \N__5318\,
            I => \N__5315\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__5315\,
            I => \N__5311\
        );

    \I__759\ : InMux
    port map (
            O => \N__5314\,
            I => \N__5308\
        );

    \I__758\ : Odrv4
    port map (
            O => \N__5311\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__5308\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\
        );

    \I__756\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5300\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__754\ : Odrv12
    port map (
            O => \N__5297\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNO_0Z0Z_0\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__5294\,
            I => \N__5290\
        );

    \I__752\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5287\
        );

    \I__751\ : InMux
    port map (
            O => \N__5290\,
            I => \N__5284\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__5287\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__5284\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\
        );

    \I__748\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5276\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__5276\,
            I => \U409_AUTOCONFIG.un1_STATE_8_0_0\
        );

    \I__746\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5267\
        );

    \I__745\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5267\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5267\,
            I => \U409_AUTOCONFIG.STATE4\
        );

    \I__743\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5255\
        );

    \I__742\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5255\
        );

    \I__741\ : InMux
    port map (
            O => \N__5262\,
            I => \N__5255\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5255\,
            I => \U409_AUTOCONFIG.un1_STATE_8Z0Z_0\
        );

    \I__739\ : InMux
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__5249\,
            I => \N__5246\
        );

    \I__737\ : Span4Mux_h
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__736\ : Odrv4
    port map (
            O => \N__5243\,
            I => \U409_AUTOCONFIG.N_248_0\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__5240\,
            I => \U409_AUTOCONFIG.un1_STATE_8Z0Z_0_cascade_\
        );

    \I__734\ : IoInMux
    port map (
            O => \N__5237\,
            I => \N__5234\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5234\,
            I => \N__5231\
        );

    \I__732\ : IoSpan4Mux
    port map (
            O => \N__5231\,
            I => \N__5228\
        );

    \I__731\ : Span4Mux_s2_h
    port map (
            O => \N__5228\,
            I => \N__5225\
        );

    \I__730\ : Sp12to4
    port map (
            O => \N__5225\,
            I => \N__5222\
        );

    \I__729\ : Span12Mux_s10_h
    port map (
            O => \N__5222\,
            I => \N__5219\
        );

    \I__728\ : Span12Mux_v
    port map (
            O => \N__5219\,
            I => \N__5216\
        );

    \I__727\ : Odrv12
    port map (
            O => \N__5216\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn_i\
        );

    \I__726\ : InMux
    port map (
            O => \N__5213\,
            I => \N__5210\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5210\,
            I => \N__5207\
        );

    \I__724\ : Span4Mux_v
    port map (
            O => \N__5207\,
            I => \N__5204\
        );

    \I__723\ : Sp12to4
    port map (
            O => \N__5204\,
            I => \N__5201\
        );

    \I__722\ : Span12Mux_h
    port map (
            O => \N__5201\,
            I => \N__5198\
        );

    \I__721\ : Odrv12
    port map (
            O => \N__5198\,
            I => \TT_c_1\
        );

    \I__720\ : InMux
    port map (
            O => \N__5195\,
            I => \N__5192\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__5192\,
            I => \N__5189\
        );

    \I__718\ : Span12Mux_h
    port map (
            O => \N__5189\,
            I => \N__5186\
        );

    \I__717\ : Span12Mux_v
    port map (
            O => \N__5186\,
            I => \N__5183\
        );

    \I__716\ : Odrv12
    port map (
            O => \N__5183\,
            I => \TT_c_0\
        );

    \I__715\ : IoInMux
    port map (
            O => \N__5180\,
            I => \N__5175\
        );

    \I__714\ : IoInMux
    port map (
            O => \N__5179\,
            I => \N__5172\
        );

    \I__713\ : IoInMux
    port map (
            O => \N__5178\,
            I => \N__5169\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__5175\,
            I => \N__5164\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__5172\,
            I => \N__5164\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5169\,
            I => \N__5161\
        );

    \I__709\ : Span4Mux_s2_v
    port map (
            O => \N__5164\,
            I => \N__5157\
        );

    \I__708\ : Span4Mux_s3_v
    port map (
            O => \N__5161\,
            I => \N__5154\
        );

    \I__707\ : IoInMux
    port map (
            O => \N__5160\,
            I => \N__5151\
        );

    \I__706\ : Span4Mux_v
    port map (
            O => \N__5157\,
            I => \N__5148\
        );

    \I__705\ : Span4Mux_h
    port map (
            O => \N__5154\,
            I => \N__5145\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5151\,
            I => \N__5142\
        );

    \I__703\ : Span4Mux_v
    port map (
            O => \N__5148\,
            I => \N__5139\
        );

    \I__702\ : Sp12to4
    port map (
            O => \N__5145\,
            I => \N__5134\
        );

    \I__701\ : Span12Mux_s4_v
    port map (
            O => \N__5142\,
            I => \N__5134\
        );

    \I__700\ : Odrv4
    port map (
            O => \N__5139\,
            I => \D_1_i\
        );

    \I__699\ : Odrv12
    port map (
            O => \N__5134\,
            I => \D_1_i\
        );

    \I__698\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5126\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5126\,
            I => \N__5122\
        );

    \I__696\ : InMux
    port map (
            O => \N__5125\,
            I => \N__5119\
        );

    \I__695\ : Odrv4
    port map (
            O => \N__5122\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__5119\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\
        );

    \I__693\ : IoInMux
    port map (
            O => \N__5114\,
            I => \N__5111\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5111\,
            I => \N__5108\
        );

    \I__691\ : Sp12to4
    port map (
            O => \N__5108\,
            I => \N__5105\
        );

    \I__690\ : Span12Mux_v
    port map (
            O => \N__5105\,
            I => \N__5102\
        );

    \I__689\ : Odrv12
    port map (
            O => \N__5102\,
            I => \U409_AUTOCONFIG_D_OUT_0_i_3\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__5099\,
            I => \AUTOCONFIG_SPACE_cascade_\
        );

    \I__687\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5093\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5093\,
            I => \U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0_a3_0\
        );

    \I__685\ : CascadeMux
    port map (
            O => \N__5090\,
            I => \N__5087\
        );

    \I__684\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5084\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__5084\,
            I => \N__5081\
        );

    \I__682\ : Span4Mux_v
    port map (
            O => \N__5081\,
            I => \N__5077\
        );

    \I__681\ : InMux
    port map (
            O => \N__5080\,
            I => \N__5074\
        );

    \I__680\ : Sp12to4
    port map (
            O => \N__5077\,
            I => \N__5069\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5074\,
            I => \N__5069\
        );

    \I__678\ : Span12Mux_v
    port map (
            O => \N__5069\,
            I => \N__5066\
        );

    \I__677\ : Odrv12
    port map (
            O => \N__5066\,
            I => \CPUCONFn_c\
        );

    \I__676\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5059\
        );

    \I__675\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5056\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__5059\,
            I => \U409_AUTOCONFIG.AC_STARTZ0\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__5056\,
            I => \U409_AUTOCONFIG.AC_STARTZ0\
        );

    \I__672\ : CascadeMux
    port map (
            O => \N__5051\,
            I => \N__5048\
        );

    \I__671\ : InMux
    port map (
            O => \N__5048\,
            I => \N__5044\
        );

    \I__670\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5041\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5044\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5041\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\
        );

    \I__667\ : IoInMux
    port map (
            O => \N__5036\,
            I => \N__5033\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__5033\,
            I => \N__5030\
        );

    \I__665\ : Span12Mux_s10_v
    port map (
            O => \N__5030\,
            I => \N__5027\
        );

    \I__664\ : Odrv12
    port map (
            O => \N__5027\,
            I => \U409_AUTOCONFIG_D_OUT_0_i_0\
        );

    \I__663\ : InMux
    port map (
            O => \N__5024\,
            I => \N__5021\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__5021\,
            I => \N__5018\
        );

    \I__661\ : Odrv4
    port map (
            O => \N__5018\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNO_0Z0Z_1\
        );

    \I__660\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5012\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__5012\,
            I => \N__5009\
        );

    \I__658\ : Span4Mux_v
    port map (
            O => \N__5009\,
            I => \N__5006\
        );

    \I__657\ : Odrv4
    port map (
            O => \N__5006\,
            I => \U409_AUTOCONFIG.N_265_0\
        );

    \I__656\ : InMux
    port map (
            O => \N__5003\,
            I => \N__4991\
        );

    \I__655\ : InMux
    port map (
            O => \N__5002\,
            I => \N__4991\
        );

    \I__654\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4984\
        );

    \I__653\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4984\
        );

    \I__652\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4984\
        );

    \I__651\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4978\
        );

    \I__650\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4978\
        );

    \I__649\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4974\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4991\,
            I => \N__4966\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__4984\,
            I => \N__4966\
        );

    \I__646\ : InMux
    port map (
            O => \N__4983\,
            I => \N__4963\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4978\,
            I => \N__4958\
        );

    \I__644\ : InMux
    port map (
            O => \N__4977\,
            I => \N__4955\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4974\,
            I => \N__4952\
        );

    \I__642\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4945\
        );

    \I__641\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4945\
        );

    \I__640\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4945\
        );

    \I__639\ : Span4Mux_h
    port map (
            O => \N__4966\,
            I => \N__4940\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__4963\,
            I => \N__4940\
        );

    \I__637\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4935\
        );

    \I__636\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4935\
        );

    \I__635\ : Span4Mux_v
    port map (
            O => \N__4958\,
            I => \N__4930\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__4955\,
            I => \N__4930\
        );

    \I__633\ : Span4Mux_v
    port map (
            O => \N__4952\,
            I => \N__4925\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__4945\,
            I => \N__4925\
        );

    \I__631\ : Span4Mux_h
    port map (
            O => \N__4940\,
            I => \N__4920\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4935\,
            I => \N__4920\
        );

    \I__629\ : Span4Mux_v
    port map (
            O => \N__4930\,
            I => \N__4917\
        );

    \I__628\ : Span4Mux_v
    port map (
            O => \N__4925\,
            I => \N__4914\
        );

    \I__627\ : Span4Mux_v
    port map (
            O => \N__4920\,
            I => \N__4911\
        );

    \I__626\ : Sp12to4
    port map (
            O => \N__4917\,
            I => \N__4906\
        );

    \I__625\ : Sp12to4
    port map (
            O => \N__4914\,
            I => \N__4906\
        );

    \I__624\ : Span4Mux_h
    port map (
            O => \N__4911\,
            I => \N__4903\
        );

    \I__623\ : Span12Mux_h
    port map (
            O => \N__4906\,
            I => \N__4898\
        );

    \I__622\ : Sp12to4
    port map (
            O => \N__4903\,
            I => \N__4898\
        );

    \I__621\ : Odrv12
    port map (
            O => \N__4898\,
            I => \A_c_2\
        );

    \I__620\ : CascadeMux
    port map (
            O => \N__4895\,
            I => \U409_AUTOCONFIG.un1_A_11Z0Z_0_cascade_\
        );

    \I__619\ : InMux
    port map (
            O => \N__4892\,
            I => \N__4889\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__4889\,
            I => \U409_AUTOCONFIG.un1_AZ0Z_11\
        );

    \I__617\ : InMux
    port map (
            O => \N__4886\,
            I => \N__4877\
        );

    \I__616\ : InMux
    port map (
            O => \N__4885\,
            I => \N__4877\
        );

    \I__615\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4874\
        );

    \I__614\ : InMux
    port map (
            O => \N__4883\,
            I => \N__4871\
        );

    \I__613\ : InMux
    port map (
            O => \N__4882\,
            I => \N__4868\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4877\,
            I => \N__4863\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__4874\,
            I => \N__4863\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4871\,
            I => \N__4858\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__4868\,
            I => \N__4858\
        );

    \I__608\ : Span4Mux_v
    port map (
            O => \N__4863\,
            I => \N__4853\
        );

    \I__607\ : Span4Mux_v
    port map (
            O => \N__4858\,
            I => \N__4850\
        );

    \I__606\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4845\
        );

    \I__605\ : InMux
    port map (
            O => \N__4856\,
            I => \N__4845\
        );

    \I__604\ : Sp12to4
    port map (
            O => \N__4853\,
            I => \N__4838\
        );

    \I__603\ : Sp12to4
    port map (
            O => \N__4850\,
            I => \N__4838\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4845\,
            I => \N__4838\
        );

    \I__601\ : Odrv12
    port map (
            O => \N__4838\,
            I => \A_c_6\
        );

    \I__600\ : CascadeMux
    port map (
            O => \N__4835\,
            I => \N__4831\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__4834\,
            I => \N__4827\
        );

    \I__598\ : InMux
    port map (
            O => \N__4831\,
            I => \N__4820\
        );

    \I__597\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4815\
        );

    \I__596\ : InMux
    port map (
            O => \N__4827\,
            I => \N__4815\
        );

    \I__595\ : InMux
    port map (
            O => \N__4826\,
            I => \N__4809\
        );

    \I__594\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4809\
        );

    \I__593\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4806\
        );

    \I__592\ : InMux
    port map (
            O => \N__4823\,
            I => \N__4803\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4820\,
            I => \N__4800\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__4815\,
            I => \N__4797\
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__4814\,
            I => \N__4794\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4809\,
            I => \N__4791\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4806\,
            I => \N__4788\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4803\,
            I => \N__4785\
        );

    \I__585\ : Span4Mux_v
    port map (
            O => \N__4800\,
            I => \N__4778\
        );

    \I__584\ : Span4Mux_v
    port map (
            O => \N__4797\,
            I => \N__4778\
        );

    \I__583\ : InMux
    port map (
            O => \N__4794\,
            I => \N__4775\
        );

    \I__582\ : Span4Mux_v
    port map (
            O => \N__4791\,
            I => \N__4770\
        );

    \I__581\ : Span4Mux_v
    port map (
            O => \N__4788\,
            I => \N__4770\
        );

    \I__580\ : Span4Mux_v
    port map (
            O => \N__4785\,
            I => \N__4767\
        );

    \I__579\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4762\
        );

    \I__578\ : InMux
    port map (
            O => \N__4783\,
            I => \N__4762\
        );

    \I__577\ : Sp12to4
    port map (
            O => \N__4778\,
            I => \N__4751\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__4775\,
            I => \N__4751\
        );

    \I__575\ : Sp12to4
    port map (
            O => \N__4770\,
            I => \N__4751\
        );

    \I__574\ : Sp12to4
    port map (
            O => \N__4767\,
            I => \N__4751\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4762\,
            I => \N__4751\
        );

    \I__572\ : Span12Mux_h
    port map (
            O => \N__4751\,
            I => \N__4748\
        );

    \I__571\ : Span12Mux_v
    port map (
            O => \N__4748\,
            I => \N__4745\
        );

    \I__570\ : Odrv12
    port map (
            O => \N__4745\,
            I => \A_c_3\
        );

    \I__569\ : InMux
    port map (
            O => \N__4742\,
            I => \N__4737\
        );

    \I__568\ : InMux
    port map (
            O => \N__4741\,
            I => \N__4732\
        );

    \I__567\ : InMux
    port map (
            O => \N__4740\,
            I => \N__4732\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4737\,
            I => \N__4727\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__4732\,
            I => \N__4724\
        );

    \I__564\ : InMux
    port map (
            O => \N__4731\,
            I => \N__4721\
        );

    \I__563\ : InMux
    port map (
            O => \N__4730\,
            I => \N__4718\
        );

    \I__562\ : Odrv4
    port map (
            O => \N__4727\,
            I => \U409_AUTOCONFIG.N_174\
        );

    \I__561\ : Odrv12
    port map (
            O => \N__4724\,
            I => \U409_AUTOCONFIG.N_174\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4721\,
            I => \U409_AUTOCONFIG.N_174\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4718\,
            I => \U409_AUTOCONFIG.N_174\
        );

    \I__558\ : InMux
    port map (
            O => \N__4709\,
            I => \N__4706\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__4706\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\
        );

    \I__556\ : InMux
    port map (
            O => \N__4703\,
            I => \N__4697\
        );

    \I__555\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4697\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__4697\,
            I => \N__4694\
        );

    \I__553\ : Odrv12
    port map (
            O => \N__4694\,
            I => \U409_ADDRESS_DECODE.REG_SPACE_3\
        );

    \I__552\ : InMux
    port map (
            O => \N__4691\,
            I => \N__4685\
        );

    \I__551\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4685\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4685\,
            I => \N__4682\
        );

    \I__549\ : Span4Mux_v
    port map (
            O => \N__4682\,
            I => \N__4679\
        );

    \I__548\ : Sp12to4
    port map (
            O => \N__4679\,
            I => \N__4676\
        );

    \I__547\ : Odrv12
    port map (
            O => \N__4676\,
            I => \A_c_25\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__4673\,
            I => \U409_ADDRESS_DECODE.REG_SPACE_3_cascade_\
        );

    \I__545\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4666\
        );

    \I__544\ : InMux
    port map (
            O => \N__4669\,
            I => \N__4663\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4666\,
            I => \N__4660\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4663\,
            I => \N__4657\
        );

    \I__541\ : Span4Mux_v
    port map (
            O => \N__4660\,
            I => \N__4654\
        );

    \I__540\ : Span4Mux_v
    port map (
            O => \N__4657\,
            I => \N__4651\
        );

    \I__539\ : Span4Mux_v
    port map (
            O => \N__4654\,
            I => \N__4648\
        );

    \I__538\ : Span4Mux_v
    port map (
            O => \N__4651\,
            I => \N__4645\
        );

    \I__537\ : Sp12to4
    port map (
            O => \N__4648\,
            I => \N__4640\
        );

    \I__536\ : Sp12to4
    port map (
            O => \N__4645\,
            I => \N__4640\
        );

    \I__535\ : Odrv12
    port map (
            O => \N__4640\,
            I => \A_c_24\
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__4637\,
            I => \N__4633\
        );

    \I__533\ : InMux
    port map (
            O => \N__4636\,
            I => \N__4628\
        );

    \I__532\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4628\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__4628\,
            I => \N__4625\
        );

    \I__530\ : Span12Mux_v
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__529\ : Odrv12
    port map (
            O => \N__4622\,
            I => \A_c_27\
        );

    \I__528\ : CascadeMux
    port map (
            O => \N__4619\,
            I => \N__4616\
        );

    \I__527\ : InMux
    port map (
            O => \N__4616\,
            I => \N__4610\
        );

    \I__526\ : InMux
    port map (
            O => \N__4615\,
            I => \N__4610\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__524\ : Span4Mux_h
    port map (
            O => \N__4607\,
            I => \N__4604\
        );

    \I__523\ : Sp12to4
    port map (
            O => \N__4604\,
            I => \N__4601\
        );

    \I__522\ : Span12Mux_v
    port map (
            O => \N__4601\,
            I => \N__4598\
        );

    \I__521\ : Odrv12
    port map (
            O => \N__4598\,
            I => \A_c_26\
        );

    \I__520\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4592\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4592\,
            I => \U409_AUTOCONFIG.N_173\
        );

    \I__518\ : CascadeMux
    port map (
            O => \N__4589\,
            I => \U409_AUTOCONFIG.N_249_1_cascade_\
        );

    \I__517\ : InMux
    port map (
            O => \N__4586\,
            I => \N__4581\
        );

    \I__516\ : InMux
    port map (
            O => \N__4585\,
            I => \N__4576\
        );

    \I__515\ : InMux
    port map (
            O => \N__4584\,
            I => \N__4576\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__4581\,
            I => \U409_AUTOCONFIG.N_155_0\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4576\,
            I => \U409_AUTOCONFIG.N_155_0\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__4571\,
            I => \N__4566\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__4570\,
            I => \N__4563\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__4569\,
            I => \N__4557\
        );

    \I__509\ : InMux
    port map (
            O => \N__4566\,
            I => \N__4548\
        );

    \I__508\ : InMux
    port map (
            O => \N__4563\,
            I => \N__4548\
        );

    \I__507\ : InMux
    port map (
            O => \N__4562\,
            I => \N__4543\
        );

    \I__506\ : InMux
    port map (
            O => \N__4561\,
            I => \N__4543\
        );

    \I__505\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4540\
        );

    \I__504\ : InMux
    port map (
            O => \N__4557\,
            I => \N__4531\
        );

    \I__503\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4531\
        );

    \I__502\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4531\
        );

    \I__501\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4531\
        );

    \I__500\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4526\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4548\,
            I => \N__4521\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4543\,
            I => \N__4521\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4540\,
            I => \N__4516\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__4531\,
            I => \N__4516\
        );

    \I__495\ : CascadeMux
    port map (
            O => \N__4530\,
            I => \N__4513\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__4529\,
            I => \N__4510\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__4526\,
            I => \N__4506\
        );

    \I__492\ : Span4Mux_v
    port map (
            O => \N__4521\,
            I => \N__4501\
        );

    \I__491\ : Span4Mux_v
    port map (
            O => \N__4516\,
            I => \N__4498\
        );

    \I__490\ : InMux
    port map (
            O => \N__4513\,
            I => \N__4495\
        );

    \I__489\ : InMux
    port map (
            O => \N__4510\,
            I => \N__4492\
        );

    \I__488\ : InMux
    port map (
            O => \N__4509\,
            I => \N__4489\
        );

    \I__487\ : Span4Mux_v
    port map (
            O => \N__4506\,
            I => \N__4486\
        );

    \I__486\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4481\
        );

    \I__485\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4481\
        );

    \I__484\ : Sp12to4
    port map (
            O => \N__4501\,
            I => \N__4466\
        );

    \I__483\ : Sp12to4
    port map (
            O => \N__4498\,
            I => \N__4466\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4495\,
            I => \N__4466\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4492\,
            I => \N__4466\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__4489\,
            I => \N__4466\
        );

    \I__479\ : Sp12to4
    port map (
            O => \N__4486\,
            I => \N__4466\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4481\,
            I => \N__4466\
        );

    \I__477\ : Odrv12
    port map (
            O => \N__4466\,
            I => \A_c_4\
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__4463\,
            I => \U409_AUTOCONFIG.un1_A_19Z0Z_1_cascade_\
        );

    \I__475\ : IoInMux
    port map (
            O => \N__4460\,
            I => \N__4457\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4457\,
            I => \N__4454\
        );

    \I__473\ : Span12Mux_s2_v
    port map (
            O => \N__4454\,
            I => \N__4451\
        );

    \I__472\ : Span12Mux_v
    port map (
            O => \N__4451\,
            I => \N__4448\
        );

    \I__471\ : Span12Mux_h
    port map (
            O => \N__4448\,
            I => \N__4445\
        );

    \I__470\ : Odrv12
    port map (
            O => \N__4445\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\
        );

    \I__469\ : InMux
    port map (
            O => \N__4442\,
            I => \N__4436\
        );

    \I__468\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4436\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4436\,
            I => \N__4433\
        );

    \I__466\ : Odrv12
    port map (
            O => \N__4433\,
            I => \U409_ADDRESS_DECODE.un2_REGSPACEn_0_0\
        );

    \I__465\ : CascadeMux
    port map (
            O => \N__4430\,
            I => \N__4426\
        );

    \I__464\ : InMux
    port map (
            O => \N__4429\,
            I => \N__4421\
        );

    \I__463\ : InMux
    port map (
            O => \N__4426\,
            I => \N__4421\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4421\,
            I => \N__4418\
        );

    \I__461\ : Odrv4
    port map (
            O => \N__4418\,
            I => \U409_ADDRESS_DECODE.REG_SPACEZ0\
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__4415\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_\
        );

    \I__459\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4409\,
            I => \U409_ADDRESS_DECODE.REG_SPACEZ0Z_0\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__4406\,
            I => \N__4403\
        );

    \I__456\ : InMux
    port map (
            O => \N__4403\,
            I => \N__4400\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4400\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_0_0\
        );

    \I__454\ : InMux
    port map (
            O => \N__4397\,
            I => \N__4394\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__4394\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_1_0\
        );

    \I__452\ : CascadeMux
    port map (
            O => \N__4391\,
            I => \U409_AUTOCONFIG.N_168_cascade_\
        );

    \I__451\ : InMux
    port map (
            O => \N__4388\,
            I => \N__4385\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4385\,
            I => \U409_AUTOCONFIG.N_167\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__4382\,
            I => \U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0_cascade_\
        );

    \I__448\ : InMux
    port map (
            O => \N__4379\,
            I => \N__4370\
        );

    \I__447\ : InMux
    port map (
            O => \N__4378\,
            I => \N__4370\
        );

    \I__446\ : InMux
    port map (
            O => \N__4377\,
            I => \N__4370\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4370\,
            I => \U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__443\ : InMux
    port map (
            O => \N__4364\,
            I => \N__4361\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__441\ : Odrv4
    port map (
            O => \N__4358\,
            I => \U409_AUTOCONFIG.N_166\
        );

    \I__440\ : InMux
    port map (
            O => \N__4355\,
            I => \N__4352\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4352\,
            I => \N__4349\
        );

    \I__438\ : Odrv4
    port map (
            O => \N__4349\,
            I => \U409_AUTOCONFIG.N_213_2\
        );

    \I__437\ : CascadeMux
    port map (
            O => \N__4346\,
            I => \U409_AUTOCONFIG.N_212_cascade_\
        );

    \I__436\ : CascadeMux
    port map (
            O => \N__4343\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_3_0_cascade_\
        );

    \I__435\ : InMux
    port map (
            O => \N__4340\,
            I => \N__4337\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__4337\,
            I => \N__4334\
        );

    \I__433\ : Odrv4
    port map (
            O => \N__4334\,
            I => \U409_AUTOCONFIG.N_165\
        );

    \I__432\ : CascadeMux
    port map (
            O => \N__4331\,
            I => \N__4328\
        );

    \I__431\ : InMux
    port map (
            O => \N__4328\,
            I => \N__4325\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__4325\,
            I => \U409_AUTOCONFIG.un1_A_16Z0Z_2\
        );

    \I__429\ : InMux
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__4319\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_0\
        );

    \I__427\ : IoInMux
    port map (
            O => \N__4316\,
            I => \N__4313\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__4313\,
            I => \N__4309\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__4312\,
            I => \N__4306\
        );

    \I__424\ : IoSpan4Mux
    port map (
            O => \N__4309\,
            I => \N__4302\
        );

    \I__423\ : InMux
    port map (
            O => \N__4306\,
            I => \N__4299\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__4305\,
            I => \N__4296\
        );

    \I__421\ : Span4Mux_s0_h
    port map (
            O => \N__4302\,
            I => \N__4293\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__4299\,
            I => \N__4290\
        );

    \I__419\ : InMux
    port map (
            O => \N__4296\,
            I => \N__4287\
        );

    \I__418\ : Sp12to4
    port map (
            O => \N__4293\,
            I => \N__4284\
        );

    \I__417\ : Span4Mux_v
    port map (
            O => \N__4290\,
            I => \N__4281\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__4287\,
            I => \N__4278\
        );

    \I__415\ : Span12Mux_v
    port map (
            O => \N__4284\,
            I => \N__4275\
        );

    \I__414\ : Sp12to4
    port map (
            O => \N__4281\,
            I => \N__4272\
        );

    \I__413\ : Span4Mux_h
    port map (
            O => \N__4278\,
            I => \N__4269\
        );

    \I__412\ : Span12Mux_h
    port map (
            O => \N__4275\,
            I => \N__4266\
        );

    \I__411\ : Span12Mux_s7_h
    port map (
            O => \N__4272\,
            I => \N__4261\
        );

    \I__410\ : Sp12to4
    port map (
            O => \N__4269\,
            I => \N__4261\
        );

    \I__409\ : Span12Mux_h
    port map (
            O => \N__4266\,
            I => \N__4256\
        );

    \I__408\ : Span12Mux_v
    port map (
            O => \N__4261\,
            I => \N__4256\
        );

    \I__407\ : Odrv12
    port map (
            O => \N__4256\,
            I => \A_c_16\
        );

    \I__406\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__4250\,
            I => \U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0\
        );

    \I__404\ : CascadeMux
    port map (
            O => \N__4247\,
            I => \U409_AUTOCONFIG.N_167_cascade_\
        );

    \I__403\ : InMux
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__4241\,
            I => \N__4238\
        );

    \I__401\ : Odrv4
    port map (
            O => \N__4238\,
            I => \U409_AUTOCONFIG.N_233\
        );

    \I__400\ : CascadeMux
    port map (
            O => \N__4235\,
            I => \U409_AUTOCONFIG.N_231_cascade_\
        );

    \I__399\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4229\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__4229\,
            I => \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_a5_0_0\
        );

    \I__397\ : InMux
    port map (
            O => \N__4226\,
            I => \N__4223\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__4223\,
            I => \U409_AUTOCONFIG.N_212\
        );

    \I__395\ : CascadeMux
    port map (
            O => \N__4220\,
            I => \U409_AUTOCONFIG.N_213_2_cascade_\
        );

    \I__394\ : CascadeMux
    port map (
            O => \N__4217\,
            I => \U409_AUTOCONFIG.N_249_cascade_\
        );

    \I__393\ : InMux
    port map (
            O => \N__4214\,
            I => \N__4211\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__4211\,
            I => \U409_AUTOCONFIG.N_250_1\
        );

    \I__391\ : InMux
    port map (
            O => \N__4208\,
            I => \N__4205\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__4205\,
            I => \U409_AUTOCONFIG.N_249\
        );

    \I__389\ : CascadeMux
    port map (
            O => \N__4202\,
            I => \U409_AUTOCONFIG.N_250_1_cascade_\
        );

    \I__388\ : IoInMux
    port map (
            O => \N__4199\,
            I => \N__4196\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__4196\,
            I => \N__4193\
        );

    \I__386\ : IoSpan4Mux
    port map (
            O => \N__4193\,
            I => \N__4190\
        );

    \I__385\ : Span4Mux_s3_h
    port map (
            O => \N__4190\,
            I => \N__4187\
        );

    \I__384\ : Sp12to4
    port map (
            O => \N__4187\,
            I => \N__4184\
        );

    \I__383\ : Span12Mux_h
    port map (
            O => \N__4184\,
            I => \N__4181\
        );

    \I__382\ : Span12Mux_h
    port map (
            O => \N__4181\,
            I => \N__4178\
        );

    \I__381\ : Odrv12
    port map (
            O => \N__4178\,
            I => \A_c_15\
        );

    \I__380\ : IoInMux
    port map (
            O => \N__4175\,
            I => \N__4172\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__4172\,
            I => \N__4169\
        );

    \I__378\ : Span4Mux_s3_h
    port map (
            O => \N__4169\,
            I => \N__4166\
        );

    \I__377\ : Span4Mux_v
    port map (
            O => \N__4166\,
            I => \N__4163\
        );

    \I__376\ : Sp12to4
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__375\ : Span12Mux_h
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__374\ : Span12Mux_h
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__373\ : Odrv12
    port map (
            O => \N__4154\,
            I => \A_c_14\
        );

    \I__372\ : ClkMux
    port map (
            O => \N__4151\,
            I => \N__4115\
        );

    \I__371\ : ClkMux
    port map (
            O => \N__4150\,
            I => \N__4115\
        );

    \I__370\ : ClkMux
    port map (
            O => \N__4149\,
            I => \N__4115\
        );

    \I__369\ : ClkMux
    port map (
            O => \N__4148\,
            I => \N__4115\
        );

    \I__368\ : ClkMux
    port map (
            O => \N__4147\,
            I => \N__4115\
        );

    \I__367\ : ClkMux
    port map (
            O => \N__4146\,
            I => \N__4115\
        );

    \I__366\ : ClkMux
    port map (
            O => \N__4145\,
            I => \N__4115\
        );

    \I__365\ : ClkMux
    port map (
            O => \N__4144\,
            I => \N__4115\
        );

    \I__364\ : ClkMux
    port map (
            O => \N__4143\,
            I => \N__4115\
        );

    \I__363\ : ClkMux
    port map (
            O => \N__4142\,
            I => \N__4115\
        );

    \I__362\ : ClkMux
    port map (
            O => \N__4141\,
            I => \N__4115\
        );

    \I__361\ : ClkMux
    port map (
            O => \N__4140\,
            I => \N__4115\
        );

    \I__360\ : GlobalMux
    port map (
            O => \N__4115\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            I => \N__4143\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            I => \N__4140\
        );

    \INVU409_AUTOCONFIG.ATA_BASE_1C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.ATA_BASE_1C_net\,
            I => \N__7943\
        );

    \INVU409_TRANSFER_ACK.TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            I => \N__4149\
        );

    \INVU409_TRANSFER_ACK.TACK_OUTnC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            I => \N__4146\
        );

    \INVU409_TRANSFER_ACK.ROMENnC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            I => \N__4144\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            I => \N__4142\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__4141\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            I => \N__4151\
        );

    \INVU409_AUTOCONFIG.LIDE_CONFC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            I => \N__7949\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            I => \N__4148\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            I => \N__4145\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            I => \N__4150\
        );

    \INVU409_AUTOCONFIG.ATA_BASE_6C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.ATA_BASE_6C_net\,
            I => \N__7948\
        );

    \INVU409_AUTOCONFIG.AC_TACKC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.AC_TACKC_net\,
            I => \N__7951\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            I => \N__4147\
        );

    \INVU409_AUTOCONFIG.STATE_1C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.STATE_1C_net\,
            I => \N__7956\
        );

    \INVU409_AUTOCONFIG.BRIDGE_BASE_3C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net\,
            I => \N__7950\
        );

    \INVU409_AUTOCONFIG.LIDE_OUT_1C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            I => \N__7955\
        );

    \INVU409_AUTOCONFIG.BRIDGE_OUT_0C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            I => \N__7964\
        );

    \IN_MUX_bfv_13_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_6_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_15_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_6_0_\
        );

    \IN_MUX_bfv_15_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_15_7_0_\
        );

    \IN_MUX_bfv_15_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_4_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8900\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_a5_0_2_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4823\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4983\,
            lcout => \U409_AUTOCONFIG.N_213_2\,
            ltout => \U409_AUTOCONFIG.N_213_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_3_1_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7062\,
            in1 => \N__4553\,
            in2 => \N__4220\,
            in3 => \N__6120\,
            lcout => \U409_AUTOCONFIG.N_233\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_141_i_a4_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6161\,
            in1 => \N__4505\,
            in2 => \N__7061\,
            in3 => \N__4962\,
            lcout => \U409_AUTOCONFIG.N_249\,
            ltout => \U409_AUTOCONFIG.N_249_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__4784\,
            in1 => \N__4214\,
            in2 => \N__4217\,
            in3 => \N__7032\,
            lcout => \U409_AUTOCONFIG.N_265_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_2_0_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4961\,
            in2 => \_gnd_net_\,
            in3 => \N__4504\,
            lcout => \U409_AUTOCONFIG.N_250_1\,
            ltout => \U409_AUTOCONFIG.N_250_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100011"
        )
    port map (
            in0 => \N__4783\,
            in1 => \N__4208\,
            in2 => \N__4202\,
            in3 => \N__7031\,
            lcout => \U409_AUTOCONFIG.N_248_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__4253\,
            in1 => \N__6492\,
            in2 => \N__5790\,
            in3 => \N__6398\,
            lcout => \U409_ADDRESS_DECODE.un2_REGSPACEn_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7441\,
            in1 => \N__7358\,
            in2 => \_gnd_net_\,
            in3 => \N__8450\,
            lcout => \U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.REG_SPACE_0_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6475\,
            in1 => \N__5818\,
            in2 => \_gnd_net_\,
            in3 => \N__6915\,
            lcout => \U409_ADDRESS_DECODE.REG_SPACEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_2_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4742\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4226\,
            lcout => \U409_AUTOCONFIG.N_167\,
            ltout => \U409_AUTOCONFIG.N_167_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__4340\,
            in1 => \N__4560\,
            in2 => \N__4247\,
            in3 => \N__4996\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6476\,
            in1 => \N__6362\,
            in2 => \N__4312\,
            in3 => \N__6926\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4999\,
            in1 => \N__4825\,
            in2 => \_gnd_net_\,
            in3 => \N__4555\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_a5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__4556\,
            in1 => \N__5000\,
            in2 => \N__6148\,
            in3 => \N__7064\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.N_231_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__7063\,
            in1 => \N__4244\,
            in2 => \N__4235\,
            in3 => \N__4232\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_85_i_a4_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__4826\,
            in1 => \N__5001\,
            in2 => \N__4569\,
            in3 => \N__7065\,
            lcout => \U409_AUTOCONFIG.N_212\,
            ltout => \U409_AUTOCONFIG.N_212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001101"
        )
    port map (
            in0 => \N__4355\,
            in1 => \N__6124\,
            in2 => \N__4346\,
            in3 => \N__4554\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__7066\,
            in1 => \N__4731\,
            in2 => \_gnd_net_\,
            in3 => \N__4971\,
            lcout => \U409_AUTOCONFIG.N_166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4972\,
            in1 => \N__6165\,
            in2 => \N__4814\,
            in3 => \N__7067\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4882\,
            in1 => \N__6225\,
            in2 => \N__4343\,
            in3 => \N__4509\,
            lcout => \U409_AUTOCONFIG.N_165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_16_2_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6166\,
            in1 => \N__6226\,
            in2 => \N__4529\,
            in3 => \N__4973\,
            lcout => \U409_AUTOCONFIG.un1_A_16Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_16_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4883\,
            in1 => \N__4824\,
            in2 => \N__4331\,
            in3 => \N__7016\,
            lcout => \U409_AUTOCONFIG.un1_AZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_6_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5545\,
            in1 => \N__4322\,
            in2 => \N__5519\,
            in3 => \N__5601\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5656\,
            in2 => \_gnd_net_\,
            in3 => \N__4669\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__4702\,
            in1 => \N__8825\,
            in2 => \N__4305\,
            in3 => \N__5810\,
            lcout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.REG_SPACE_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4703\,
            in1 => \N__4412\,
            in2 => \N__8472\,
            in3 => \N__6391\,
            lcout => \U409_ADDRESS_DECODE.REG_SPACEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__4397\,
            in1 => \N__5047\,
            in2 => \N__4406\,
            in3 => \N__4377\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__4998\,
            in1 => \N__4741\,
            in2 => \N__4571\,
            in3 => \N__4585\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000000000"
        )
    port map (
            in0 => \N__4997\,
            in1 => \N__4740\,
            in2 => \N__4570\,
            in3 => \N__7069\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.N_168_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000001100"
        )
    port map (
            in0 => \N__5125\,
            in1 => \N__10919\,
            in2 => \N__4391\,
            in3 => \N__4379\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_RNI10V92_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010101010"
        )
    port map (
            in0 => \N__10918\,
            in1 => \N__5096\,
            in2 => \N__5090\,
            in3 => \N__5063\,
            lcout => \U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0\,
            ltout => \U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__4388\,
            in1 => \N__4586\,
            in2 => \N__4382\,
            in3 => \N__5341\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__4378\,
            in1 => \N__4584\,
            in2 => \N__4367\,
            in3 => \N__5395\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_3_0_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6221\,
            in1 => \N__4857\,
            in2 => \_gnd_net_\,
            in3 => \N__6149\,
            lcout => \U409_AUTOCONFIG.N_173\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.ATA_BASE11_1_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4561\,
            in1 => \N__4856\,
            in2 => \N__4835\,
            in3 => \N__5002\,
            lcout => \U409_AUTOCONFIG.ATA_BASE11Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_6_2_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5003\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4562\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.N_249_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_o3_0_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001001100"
        )
    port map (
            in0 => \N__4595\,
            in1 => \N__10917\,
            in2 => \N__4589\,
            in3 => \N__7068\,
            lcout => \U409_AUTOCONFIG.N_155_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_19_1_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101101"
        )
    port map (
            in0 => \N__6158\,
            in1 => \N__6222\,
            in2 => \N__4530\,
            in3 => \N__4884\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.un1_A_19Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_STATE_8_0_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__4892\,
            in1 => \N__4730\,
            in2 => \N__4463\,
            in3 => \N__8252\,
            lcout => \U409_AUTOCONFIG.un1_STATE_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_1_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__5980\,
            in1 => \N__5925\,
            in2 => \N__7639\,
            in3 => \N__7600\,
            lcout => \U409_ADDRESS_DECODE_ROMEN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111110111111"
        )
    port map (
            in0 => \N__4442\,
            in1 => \N__5982\,
            in2 => \N__5939\,
            in3 => \N__4429\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000000000"
        )
    port map (
            in0 => \N__5981\,
            in1 => \N__4441\,
            in2 => \N__4430\,
            in3 => \N__5926\,
            lcout => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__7632\,
            in1 => \N__7370\,
            in2 => \_gnd_net_\,
            in3 => \N__7599\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\,
            ltout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7476\,
            in1 => \N__5924\,
            in2 => \N__4415\,
            in3 => \N__5979\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACE_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_11_0_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4886\,
            in1 => \N__7024\,
            in2 => \_gnd_net_\,
            in3 => \N__6224\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.un1_A_11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_11_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4830\,
            in1 => \N__4977\,
            in2 => \N__4895\,
            in3 => \N__6160\,
            lcout => \U409_AUTOCONFIG.un1_AZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_0_0_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6223\,
            in1 => \N__4885\,
            in2 => \N__4834\,
            in3 => \N__6159\,
            lcout => \U409_AUTOCONFIG.N_174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_4_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5791\,
            in1 => \N__4709\,
            in2 => \N__7480\,
            in3 => \N__6943\,
            lcout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__10933\,
            in1 => \N__4636\,
            in2 => \N__4619\,
            in3 => \N__4691\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7354\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7454\,
            lcout => \U409_ADDRESS_DECODE.REG_SPACE_3\,
            ltout => \U409_ADDRESS_DECODE.REG_SPACE_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5437\,
            in1 => \N__4690\,
            in2 => \N__4673\,
            in3 => \N__4670\,
            lcout => \U409_ADDRESS_DECODE_AUTOVECTOR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5544\,
            in1 => \N__5518\,
            in2 => \N__4637\,
            in3 => \N__4615\,
            lcout => \U409_ADDRESS_DECODE_AUTOVECTOR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.D_1_i_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9070\,
            in1 => \N__9028\,
            in2 => \_gnd_net_\,
            in3 => \N__8261\,
            lcout => \D_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIG8DB1_3_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__5129\,
            in1 => \N__5318\,
            in2 => \N__8360\,
            in3 => \N__6653\,
            lcout => \U409_AUTOCONFIG_D_OUT_0_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8491\,
            in1 => \N__6496\,
            in2 => \N__6402\,
            in3 => \N__6936\,
            lcout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9069\,
            in2 => \_gnd_net_\,
            in3 => \N__9027\,
            lcout => OPEN,
            ltout => \AUTOCONFIG_SPACE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__7245\,
            in1 => \N__10888\,
            in2 => \N__5099\,
            in3 => \N__8350\,
            lcout => \U409_AUTOCONFIG.AC_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIBIND1_0_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__8253\,
            in1 => \N__6076\,
            in2 => \_gnd_net_\,
            in3 => \N__6026\,
            lcout => \U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_RNI04BC_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5080\,
            in2 => \_gnd_net_\,
            in3 => \N__5062\,
            lcout => \U409_AUTOCONFIG.STATE4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIA2DB1_0_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__8351\,
            in1 => \N__5293\,
            in2 => \N__5051\,
            in3 => \N__6652\,
            lcout => \U409_AUTOCONFIG_D_OUT_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_1_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__5024\,
            in1 => \N__5380\,
            in2 => \N__10915\,
            in3 => \N__5263\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__5264\,
            in1 => \N__5015\,
            in2 => \N__10929\,
            in3 => \N__5314\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_0_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__5273\,
            in1 => \N__6031\,
            in2 => \N__10916\,
            in3 => \N__6078\,
            lcout => \U409_AUTOCONFIG.STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_0_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__10889\,
            in1 => \N__5303\,
            in2 => \N__5294\,
            in3 => \N__5262\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIILDD3_0_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6077\,
            in1 => \N__5279\,
            in2 => \N__6037\,
            in3 => \N__5272\,
            lcout => \U409_AUTOCONFIG.un1_STATE_8Z0Z_0\,
            ltout => \U409_AUTOCONFIG.un1_STATE_8Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_2_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__10893\,
            in1 => \N__5252\,
            in2 => \N__5240\,
            in3 => \N__5356\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__8053\,
            in1 => \N__8117\,
            in2 => \N__5564\,
            in3 => \N__6545\,
            lcout => \BRIDGE_BASE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net\,
            ce => 'H',
            sr => \N__8573\
        );

    \U409_AUTOCONFIG.ATA_BASE_7_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__8116\,
            in1 => \N__5738\,
            in2 => \N__8054\,
            in3 => \N__7114\,
            lcout => \ATA_BASE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net\,
            ce => 'H',
            sr => \N__8573\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__5462\,
            in1 => \N__5941\,
            in2 => \N__5989\,
            in3 => \N__5468\,
            lcout => \U409_ADDRESS_DECODE_un1_RTC_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5474\,
            in1 => \N__5213\,
            in2 => \N__10934\,
            in3 => \N__5195\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_3_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5808\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8473\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__8475\,
            in1 => \N__6497\,
            in2 => \_gnd_net_\,
            in3 => \N__6403\,
            lcout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0\,
            ltout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5940\,
            in1 => \N__5461\,
            in2 => \N__5450\,
            in3 => \N__5972\,
            lcout => \U409_ADDRESS_DECODE_un1_RTC_ENn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5809\,
            in1 => \N__5447\,
            in2 => \N__5441\,
            in3 => \N__8474\,
            lcout => \CIA_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5657\,
            in1 => \N__5420\,
            in2 => \_gnd_net_\,
            in3 => \N__5614\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE_AUTOVECTOR_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_AUTOVECTOR_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__5414\,
            in1 => \N__6874\,
            in2 => \N__5408\,
            in3 => \N__5405\,
            lcout => \U409_TRANSFER_ACK.un1_AUTOVECTOR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIC4DB1_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__5399\,
            in1 => \N__6650\,
            in2 => \N__5384\,
            in3 => \N__8352\,
            lcout => \U409_AUTOCONFIG_D_OUT_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIE6DB1_2_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011100100"
        )
    port map (
            in0 => \N__6651\,
            in1 => \N__5357\,
            in2 => \N__8359\,
            in3 => \N__5345\,
            lcout => \U409_AUTOCONFIG_D_OUT_0_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_1_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000011000000"
        )
    port map (
            in0 => \N__8259\,
            in1 => \N__6079\,
            in2 => \N__10914\,
            in3 => \N__6032\,
            lcout => \U409_AUTOCONFIG.STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6074\,
            in2 => \_gnd_net_\,
            in3 => \N__6027\,
            lcout => \U409_AUTOCONFIG.STATE_d_2\,
            ltout => \U409_AUTOCONFIG.STATE_d_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__6681\,
            in1 => \_gnd_net_\,
            in2 => \N__5660\,
            in3 => \N__6631\,
            lcout => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_2_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__5649\,
            in1 => \N__5615\,
            in2 => \N__5845\,
            in3 => \N__5563\,
            lcout => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIDFPA3_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__7070\,
            in1 => \N__7082\,
            in2 => \_gnd_net_\,
            in3 => \N__6646\,
            lcout => \U409_AUTOCONFIG.LIDE_CONF_RNIDFPAZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_1_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__6515\,
            in1 => \N__5549\,
            in2 => \N__5514\,
            in3 => \N__6566\,
            lcout => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_0_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5824\,
            in1 => \N__8492\,
            in2 => \_gnd_net_\,
            in3 => \N__6477\,
            lcout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2_0_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6478\,
            in1 => \N__7463\,
            in2 => \_gnd_net_\,
            in3 => \N__5825\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__7313\,
            in1 => \N__7386\,
            in2 => \N__5477\,
            in3 => \N__8493\,
            lcout => \U409_TRANSFER_ACK.N_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__6292\,
            in1 => \N__5687\,
            in2 => \N__6823\,
            in3 => \N__6316\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__9131\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6314\,
            in1 => \N__6291\,
            in2 => \N__6248\,
            in3 => \N__6725\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_6_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__7999\,
            in1 => \N__7252\,
            in2 => \N__5711\,
            in3 => \N__6262\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__6315\,
            in1 => \N__5704\,
            in2 => \N__5708\,
            in3 => \N__6769\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__9131\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__5705\,
            in1 => \N__6326\,
            in2 => \N__6822\,
            in3 => \N__6740\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__9131\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5703\,
            in1 => \N__6768\,
            in2 => \_gnd_net_\,
            in3 => \N__6811\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__9131\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_1_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6719\,
            in1 => \N__7706\,
            in2 => \N__6794\,
            in3 => \N__7675\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_6_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5690\,
            in3 => \N__6767\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_TACK_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111010100000"
        )
    port map (
            in0 => \N__6080\,
            in1 => \N__8260\,
            in2 => \N__7792\,
            in3 => \N__6038\,
            lcout => \AC_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.AC_TACKC_net\,
            ce => 'H',
            sr => \N__8574\
        );

    \U409_AUTOCONFIG.CONFIGENn_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5671\,
            in2 => \_gnd_net_\,
            in3 => \N__6543\,
            lcout => \CONFIGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.AC_TACKC_net\,
            ce => 'H',
            sr => \N__8574\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNI0EA21_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6230\,
            in1 => \N__6176\,
            in2 => \N__6167\,
            in3 => \N__6616\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.ATA_BASE11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIDSPQ2_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__6682\,
            in1 => \N__6075\,
            in2 => \N__6041\,
            in3 => \N__6033\,
            lcout => \U409_AUTOCONFIG.un1_STATE_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000001000"
        )
    port map (
            in0 => \N__5990\,
            in1 => \N__5942\,
            in2 => \N__7462\,
            in3 => \N__5887\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.ATA_BASE_6_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__5888\,
            in1 => \N__5877\,
            in2 => \N__8115\,
            in3 => \N__5737\,
            lcout => \ATA_BASE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_6C_net\,
            ce => 'H',
            sr => \N__8570\
        );

    \U409_AUTOCONFIG.ATA_BASE_2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__8097\,
            in1 => \N__8130\,
            in2 => \N__5879\,
            in3 => \N__7130\,
            lcout => \ATA_BASE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_6C_net\,
            ce => 'H',
            sr => \N__8570\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__5878\,
            in1 => \N__8107\,
            in2 => \N__5846\,
            in3 => \N__6544\,
            lcout => \BRIDGE_BASE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_6C_net\,
            ce => 'H',
            sr => \N__8570\
        );

    \U409_AUTOCONFIG.ATA_BASE_4_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__5747\,
            in1 => \N__6592\,
            in2 => \N__8113\,
            in3 => \N__5735\,
            lcout => \ATA_BASE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_6C_net\,
            ce => 'H',
            sr => \N__8570\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__8479\,
            in1 => \N__5719\,
            in2 => \N__5817\,
            in3 => \N__5746\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.ATA_BASE_5_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__5720\,
            in1 => \N__8190\,
            in2 => \N__8114\,
            in3 => \N__5736\,
            lcout => \ATA_BASE_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_6C_net\,
            ce => 'H',
            sr => \N__8570\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__6335\,
            in1 => \N__6838\,
            in2 => \_gnd_net_\,
            in3 => \N__6269\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            ce => 'H',
            sr => \N__9127\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7270\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7235\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__7998\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7256\,
            lcout => \U409_TRANSFER_ACK.N_33_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_7_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6293\,
            in1 => \N__6317\,
            in2 => \_gnd_net_\,
            in3 => \N__6766\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8835\,
            in1 => \N__8854\,
            in2 => \_gnd_net_\,
            in3 => \N__8671\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_3_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6789\,
            in1 => \N__6765\,
            in2 => \N__7708\,
            in3 => \N__6313\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_7_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6290\,
            in1 => \N__6739\,
            in2 => \N__6272\,
            in3 => \N__6241\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010100000101"
        )
    port map (
            in0 => \N__7702\,
            in1 => \N__7234\,
            in2 => \N__6251\,
            in3 => \N__7997\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__9126\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_1_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7673\,
            in2 => \_gnd_net_\,
            in3 => \N__6713\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__7674\,
            in1 => \_gnd_net_\,
            in2 => \N__7709\,
            in3 => \N__6818\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__9126\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__7655\,
            in1 => \N__6790\,
            in2 => \N__6824\,
            in3 => \N__6714\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__9126\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_7_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6788\,
            in1 => \N__7698\,
            in2 => \N__6770\,
            in3 => \N__6738\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7654\,
            in2 => \_gnd_net_\,
            in3 => \N__6718\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__9125\
        );

    \U409_AUTOCONFIG.LIDE_CONF_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__6695\,
            in1 => \N__6686\,
            in2 => \_gnd_net_\,
            in3 => \N__6630\,
            lcout => \U409_AUTOCONFIG.LIDE_CONFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__8571\
        );

    \U409_AUTOCONFIG.CONFIGURED_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__6546\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8333\,
            lcout => \CONFIGURED\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__8571\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__6547\,
            in1 => \N__8095\,
            in2 => \N__6596\,
            in3 => \N__6559\,
            lcout => \BRIDGE_BASE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__8571\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__8096\,
            in1 => \N__6548\,
            in2 => \N__8191\,
            in3 => \N__6508\,
            lcout => \BRIDGE_BASE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__8571\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__6491\,
            in1 => \N__8014\,
            in2 => \N__6404\,
            in3 => \N__7129\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_5_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000010000"
        )
    port map (
            in0 => \N__7380\,
            in1 => \N__6884\,
            in2 => \N__7118\,
            in3 => \N__7115\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7100\,
            in1 => \N__7094\,
            in2 => \N__7088\,
            in3 => \N__8306\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0\,
            ltout => \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000100000"
        )
    port map (
            in0 => \N__10871\,
            in1 => \N__8257\,
            in2 => \N__7085\,
            in3 => \N__9240\,
            lcout => \U409_ADDRESS_DECODE.ATA_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7947\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIS3FU2_0_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7081\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7060\,
            lcout => \U409_AUTOCONFIG.STATE_RNIS3FU2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un2_ATA_SPACE_0_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__6947\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8143\,
            lcout => \U409_ADDRESS_DECODE.un2_ATA_SPACEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__9084\,
            in1 => \N__6878\,
            in2 => \N__9053\,
            in3 => \N__9328\,
            lcout => \U409_ADDRESS_DECODE_PORTSIZE_0\,
            ltout => \U409_ADDRESS_DECODE_PORTSIZE_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNI4345U_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111110101111"
        )
    port map (
            in0 => \N__8539\,
            in1 => \N__9213\,
            in2 => \N__6863\,
            in3 => \N__9241\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6839\,
            in3 => \N__7165\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7274\,
            in1 => \N__7236\,
            in2 => \N__8002\,
            in3 => \N__7174\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \N__8567\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__7181\,
            in1 => \N__7175\,
            in2 => \N__8003\,
            in3 => \N__7166\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \N__8567\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__8000\,
            in1 => \N__7569\,
            in2 => \_gnd_net_\,
            in3 => \N__7555\,
            lcout => \U409_TRANSFER_ACK.N_17_mux\,
            ltout => \U409_TRANSFER_ACK.N_17_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101011111"
        )
    port map (
            in0 => \N__7540\,
            in1 => \N__7872\,
            in2 => \N__7154\,
            in3 => \N__7889\,
            lcout => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7570\,
            in2 => \_gnd_net_\,
            in3 => \N__7556\,
            lcout => \U409_TRANSFER_ACK.N_3_0\,
            ltout => \U409_TRANSFER_ACK.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__7544\,
            in1 => \N__7873\,
            in2 => \N__7151\,
            in3 => \N__7891\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000101010"
        )
    port map (
            in0 => \N__10816\,
            in1 => \N__7516\,
            in2 => \N__7148\,
            in3 => \N__7145\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000011111"
        )
    port map (
            in0 => \N__7874\,
            in1 => \N__7890\,
            in2 => \N__7547\,
            in3 => \N__7139\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.N_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101000001000"
        )
    port map (
            in0 => \N__10817\,
            in1 => \N__7515\,
            in2 => \N__7133\,
            in3 => \N__7545\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10180\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__8576\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7571\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__8576\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111100001000"
        )
    port map (
            in0 => \N__7546\,
            in1 => \N__7523\,
            in2 => \N__7517\,
            in3 => \N__7810\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__8576\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_0_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__7387\,
            in1 => \N__8842\,
            in2 => \_gnd_net_\,
            in3 => \N__7486\,
            lcout => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8389\,
            in1 => \N__7499\,
            in2 => \N__7490\,
            in3 => \N__7388\,
            lcout => \U409_TRANSFER_ACK.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__7285\,
            in1 => \N__8705\,
            in2 => \_gnd_net_\,
            in3 => \N__8774\,
            lcout => \ROMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            ce => 'H',
            sr => \N__8572\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8730\,
            in2 => \_gnd_net_\,
            in3 => \N__8765\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            ce => 'H',
            sr => \N__8572\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100011001100"
        )
    port map (
            in0 => \N__8767\,
            in1 => \N__8673\,
            in2 => \N__8741\,
            in3 => \N__8699\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            ce => 'H',
            sr => \N__8572\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011110010"
        )
    port map (
            in0 => \N__8639\,
            in1 => \N__8768\,
            in2 => \N__7826\,
            in3 => \N__8737\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            ce => 'H',
            sr => \N__8572\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101110100000"
        )
    port map (
            in0 => \N__8766\,
            in1 => \N__8672\,
            in2 => \N__8740\,
            in3 => \N__8698\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            ce => 'H',
            sr => \N__8572\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100000"
        )
    port map (
            in0 => \N__7832\,
            in1 => \N__8738\,
            in2 => \N__8794\,
            in3 => \N__8867\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            ce => 'H',
            sr => \N__8572\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__7822\,
            in1 => \N__7811\,
            in2 => \N__7796\,
            in3 => \N__7775\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER6\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111011101"
        )
    port map (
            in0 => \N__8627\,
            in1 => \N__8594\,
            in2 => \N__7763\,
            in3 => \N__7722\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__7723\,
            in1 => \_gnd_net_\,
            in2 => \N__7760\,
            in3 => \N__10880\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI7S9R_1_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7707\,
            in2 => \_gnd_net_\,
            in3 => \N__7676\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_1_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__8595\,
            in1 => \N__10879\,
            in2 => \_gnd_net_\,
            in3 => \N__8628\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000110000"
        )
    port map (
            in0 => \N__8630\,
            in1 => \N__8597\,
            in2 => \N__10913\,
            in3 => \N__8608\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7643\,
            in1 => \N__7604\,
            in2 => \_gnd_net_\,
            in3 => \N__8327\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1\,
            ltout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__8300\,
            in1 => \N__8288\,
            in2 => \N__8279\,
            in3 => \N__10884\,
            lcout => \U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__8258\,
            in1 => \N__9091\,
            in2 => \_gnd_net_\,
            in3 => \N__9051\,
            lcout => \un1_AUTOCONFIG_SPACE\,
            ltout => \un1_AUTOCONFIG_SPACE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.ATA_BASE_1_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__8192\,
            in1 => \N__8131\,
            in2 => \N__8147\,
            in3 => \N__8144\,
            lcout => \ATA_BASE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_1C_net\,
            ce => 'H',
            sr => \N__8568\
        );

    \U409_AUTOCONFIG.ATA_BASE_3_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__8132\,
            in1 => \N__8070\,
            in2 => \N__8038\,
            in3 => \N__8015\,
            lcout => \ATA_BASE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_1C_net\,
            ce => 'H',
            sr => \N__8568\
        );

    \GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8001\,
            lcout => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10963\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10793\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__8575\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7892\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__8575\
        );

    \U409_TICK.TICK50_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__9836\,
            in1 => \N__7843\,
            in2 => \N__9781\,
            in3 => \N__9884\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10566\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__8382\,
            in1 => \N__8512\,
            in2 => \_gnd_net_\,
            in3 => \N__8501\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011010"
        )
    port map (
            in0 => \N__8696\,
            in1 => \_gnd_net_\,
            in2 => \N__8675\,
            in3 => \N__8762\,
            lcout => \U409_TRANSFER_ACK.N_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8861\,
            in1 => \N__8663\,
            in2 => \N__8843\,
            in3 => \N__8694\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8798\,
            in1 => \N__8726\,
            in2 => \N__8777\,
            in3 => \N__8763\,
            lcout => \U409_TRANSFER_ACK.N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__8764\,
            in1 => \N__8670\,
            in2 => \N__8739\,
            in3 => \N__8697\,
            lcout => \U409_TRANSFER_ACK.N_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__8695\,
            in1 => \_gnd_net_\,
            in2 => \N__8674\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011110001"
        )
    port map (
            in0 => \N__8629\,
            in1 => \N__8609\,
            in2 => \N__8946\,
            in3 => \N__8596\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            ce => 'H',
            sr => \N__8569\
        );

    \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010001"
        )
    port map (
            in0 => \N__8540\,
            in1 => \N__8519\,
            in2 => \N__8500\,
            in3 => \N__8393\,
            lcout => \AGNUS_SPACE_0\,
            ltout => \AGNUS_SPACE_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__10825\,
            in1 => \_gnd_net_\,
            in2 => \N__9149\,
            in3 => \N__9146\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.LV_SPACE_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__9092\,
            in1 => \N__9052\,
            in2 => \N__8981\,
            in3 => \N__9224\,
            lcout => \BUFENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_RNI2ED4S_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__8990\,
            in1 => \N__8980\,
            in2 => \_gnd_net_\,
            in3 => \N__8947\,
            lcout => \TCIn_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10826\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9378\,
            in2 => \N__9636\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_6_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9412\,
            in2 => \_gnd_net_\,
            in3 => \N__8888\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__10564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9571\,
            in2 => \_gnd_net_\,
            in3 => \N__8885\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__10564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9607\,
            in2 => \_gnd_net_\,
            in3 => \N__8882\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9649\,
            in2 => \_gnd_net_\,
            in3 => \N__9176\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__10564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9707\,
            in3 => \N__9173\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9256\,
            in2 => \_gnd_net_\,
            in3 => \N__9170\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__10564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9688\,
            in2 => \_gnd_net_\,
            in3 => \N__9167\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9718\,
            in2 => \_gnd_net_\,
            in3 => \N__9164\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9274\,
            in2 => \_gnd_net_\,
            in3 => \N__9161\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__10565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9589\,
            in2 => \_gnd_net_\,
            in3 => \N__9158\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__10565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9424\,
            in2 => \_gnd_net_\,
            in3 => \N__9155\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__10565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9286\,
            in2 => \_gnd_net_\,
            in3 => \N__9152\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__10565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9448\,
            in2 => \_gnd_net_\,
            in3 => \N__9296\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9668\,
            in3 => \N__9293\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9401\,
            in2 => \_gnd_net_\,
            in3 => \N__9290\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__9287\,
            in1 => \N__9275\,
            in2 => \N__9263\,
            in3 => \N__9667\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNI206O6_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__9245\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9220\,
            lcout => \U409_ADDRESS_DECODE_un1_ATA_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9818\,
            in1 => \N__9883\,
            in2 => \N__9777\,
            in3 => \N__10310\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__10298\,
            in1 => \N__10631\,
            in2 => \N__10367\,
            in3 => \N__10610\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_1_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__9999\,
            in1 => \N__10146\,
            in2 => \N__10087\,
            in3 => \N__10126\,
            lcout => OPEN,
            ltout => \U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010000000"
        )
    port map (
            in0 => \N__10027\,
            in1 => \N__10537\,
            in2 => \N__9179\,
            in3 => \N__10509\,
            lcout => OPEN,
            ltout => \U409_CIA.VMA_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__10510\,
            in1 => \N__9341\,
            in2 => \N__9314\,
            in3 => \N__10950\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9979\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__10349\,
            in1 => \N__10382\,
            in2 => \_gnd_net_\,
            in3 => \N__9944\,
            lcout => \U409_TICK.TICK503_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__9869\,
            in1 => \N__9815\,
            in2 => \N__10598\,
            in3 => \N__9761\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9816\,
            in1 => \N__9870\,
            in2 => \N__9775\,
            in3 => \N__10337\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10328\,
            in1 => \N__10223\,
            in2 => \N__10268\,
            in3 => \N__10652\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__9814\,
            in1 => \N__9868\,
            in2 => \N__9311\,
            in3 => \N__9945\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10283\,
            in1 => \N__9923\,
            in2 => \N__9965\,
            in3 => \N__10582\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__9308\,
            in1 => \N__10667\,
            in2 => \N__9302\,
            in3 => \N__10238\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9817\,
            in1 => \N__9760\,
            in2 => \N__9299\,
            in3 => \N__10619\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9964\,
            in2 => \_gnd_net_\,
            in3 => \N__9946\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__9523\,
            in1 => \N__9556\,
            in2 => \N__9637\,
            in3 => \N__9482\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9554\,
            in1 => \N__9525\,
            in2 => \N__9493\,
            in3 => \N__9437\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__9872\,
            in1 => \N__9831\,
            in2 => \N__10253\,
            in3 => \N__9765\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9555\,
            in1 => \N__9526\,
            in2 => \N__9494\,
            in3 => \N__9431\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9425\,
            in1 => \N__9413\,
            in2 => \N__9383\,
            in3 => \N__9400\,
            lcout => \U409_TICK.TICK603_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9553\,
            in1 => \N__9524\,
            in2 => \N__9492\,
            in3 => \N__9389\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__9382\,
            in1 => \_gnd_net_\,
            in2 => \N__9638\,
            in3 => \_gnd_net_\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9830\,
            in1 => \N__9871\,
            in2 => \N__9776\,
            in3 => \N__10640\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__9481\,
            in1 => \N__9352\,
            in2 => \N__9560\,
            in3 => \N__9518\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9551\,
            in1 => \N__9480\,
            in2 => \N__9527\,
            in3 => \N__9890\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9882\,
            in1 => \N__9832\,
            in2 => \N__9782\,
            in3 => \N__10208\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9719\,
            in1 => \N__9706\,
            in2 => \N__9692\,
            in3 => \N__9449\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__9677\,
            in1 => \N__9552\,
            in2 => \N__9671\,
            in3 => \N__9522\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__9653\,
            in1 => \N__9629\,
            in2 => \_gnd_net_\,
            in3 => \N__9608\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__9596\,
            in1 => \N__9590\,
            in2 => \N__9578\,
            in3 => \N__9575\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9517\,
            in1 => \N__9479\,
            in2 => \N__9458\,
            in3 => \N__9455\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10503\,
            in2 => \N__10127\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_4_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10145\,
            in2 => \_gnd_net_\,
            in3 => \N__9908\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__9980\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9998\,
            in2 => \_gnd_net_\,
            in3 => \N__9905\,
            lcout => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10535\,
            in2 => \_gnd_net_\,
            in3 => \N__9902\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__9980\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10082\,
            in2 => \_gnd_net_\,
            in3 => \N__9899\,
            lcout => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_6_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10046\,
            in2 => \_gnd_net_\,
            in3 => \N__9896\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\,
            clk => \N__9980\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_7_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10061\,
            in2 => \_gnd_net_\,
            in3 => \N__9893\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9980\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__10504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10122\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9980\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_1_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000010000"
        )
    port map (
            in0 => \N__10001\,
            in1 => \N__10148\,
            in2 => \N__10179\,
            in3 => \N__10538\,
            lcout => \U409_CIA.CLK_CIA_r_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10125\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9978\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_0_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10045\,
            in1 => \N__10124\,
            in2 => \N__10514\,
            in3 => \N__10060\,
            lcout => OPEN,
            ltout => \U409_CIA.CLK_CIA6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001101010"
        )
    port map (
            in0 => \N__10172\,
            in1 => \N__10202\,
            in2 => \N__10196\,
            in3 => \N__10086\,
            lcout => \CLK_CIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9978\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__10000\,
            in1 => \N__10147\,
            in2 => \N__10088\,
            in3 => \N__10123\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_2_0\,
            ltout => \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10478\,
            in1 => \N__10028\,
            in2 => \N__10097\,
            in3 => \N__10094\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9978\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10059\,
            in2 => \_gnd_net_\,
            in3 => \N__10044\,
            lcout => \U409_CIA.CLK_CIA6_4\,
            ltout => \U409_CIA.CLK_CIA6_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10016\,
            in1 => \N__10477\,
            in2 => \N__10010\,
            in3 => \N__10007\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9978\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9960\,
            in2 => \N__9947\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_6_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9922\,
            in2 => \_gnd_net_\,
            in3 => \N__9911\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__10569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10381\,
            in2 => \_gnd_net_\,
            in3 => \N__10370\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__10569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10363\,
            in2 => \_gnd_net_\,
            in3 => \N__10352\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__10569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10348\,
            in2 => \_gnd_net_\,
            in3 => \N__10331\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10327\,
            in2 => \_gnd_net_\,
            in3 => \N__10301\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10297\,
            in2 => \_gnd_net_\,
            in3 => \N__10286\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__10569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10282\,
            in2 => \_gnd_net_\,
            in3 => \N__10271\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__10569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10264\,
            in2 => \_gnd_net_\,
            in3 => \N__10241\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_15_7_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10237\,
            in2 => \_gnd_net_\,
            in3 => \N__10226\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__10571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10219\,
            in2 => \_gnd_net_\,
            in3 => \N__10670\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10666\,
            in2 => \_gnd_net_\,
            in3 => \N__10655\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__10571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10651\,
            in2 => \_gnd_net_\,
            in3 => \N__10634\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10630\,
            in2 => \_gnd_net_\,
            in3 => \N__10613\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10609\,
            in2 => \_gnd_net_\,
            in3 => \N__10589\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10583\,
            in2 => \_gnd_net_\,
            in3 => \N__10586\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10536\,
            in2 => \_gnd_net_\,
            in3 => \N__10505\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_24_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_24_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__10736\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10426\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS1n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNI692L_0_LC_24_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10967\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10773\,
            lcout => \CIA_ENABLE\,
            ltout => \CIA_ENABLE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_24_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__10723\,
            in1 => \_gnd_net_\,
            in2 => \N__10688\,
            in3 => \_gnd_net_\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS0n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

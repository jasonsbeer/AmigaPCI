// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Feb 2 2025 09:29:49

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    CMA,
    DRA,
    SIZ,
    A,
    TSn,
    DMA_LATCH,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    LDSn,
    LATCH_CLK,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    DBRn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    output [10:0] CMA;
    input [9:0] DRA;
    input [1:0] SIZ;
    input [20:0] A;
    input TSn;
    output DMA_LATCH;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    input DBRn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__11197;
    wire N__11196;
    wire N__11195;
    wire N__11188;
    wire N__11187;
    wire N__11186;
    wire N__11179;
    wire N__11178;
    wire N__11177;
    wire N__11170;
    wire N__11169;
    wire N__11168;
    wire N__11161;
    wire N__11160;
    wire N__11159;
    wire N__11152;
    wire N__11151;
    wire N__11150;
    wire N__11143;
    wire N__11142;
    wire N__11141;
    wire N__11134;
    wire N__11133;
    wire N__11132;
    wire N__11125;
    wire N__11124;
    wire N__11123;
    wire N__11116;
    wire N__11115;
    wire N__11114;
    wire N__11107;
    wire N__11106;
    wire N__11105;
    wire N__11098;
    wire N__11097;
    wire N__11096;
    wire N__11089;
    wire N__11088;
    wire N__11087;
    wire N__11080;
    wire N__11079;
    wire N__11078;
    wire N__11071;
    wire N__11070;
    wire N__11069;
    wire N__11062;
    wire N__11061;
    wire N__11060;
    wire N__11053;
    wire N__11052;
    wire N__11051;
    wire N__11044;
    wire N__11043;
    wire N__11042;
    wire N__11035;
    wire N__11034;
    wire N__11033;
    wire N__11026;
    wire N__11025;
    wire N__11024;
    wire N__11017;
    wire N__11016;
    wire N__11015;
    wire N__11008;
    wire N__11007;
    wire N__11006;
    wire N__10999;
    wire N__10998;
    wire N__10997;
    wire N__10990;
    wire N__10989;
    wire N__10988;
    wire N__10981;
    wire N__10980;
    wire N__10979;
    wire N__10972;
    wire N__10971;
    wire N__10970;
    wire N__10963;
    wire N__10962;
    wire N__10961;
    wire N__10954;
    wire N__10953;
    wire N__10952;
    wire N__10945;
    wire N__10944;
    wire N__10943;
    wire N__10936;
    wire N__10935;
    wire N__10934;
    wire N__10927;
    wire N__10926;
    wire N__10925;
    wire N__10918;
    wire N__10917;
    wire N__10916;
    wire N__10909;
    wire N__10908;
    wire N__10907;
    wire N__10900;
    wire N__10899;
    wire N__10898;
    wire N__10891;
    wire N__10890;
    wire N__10889;
    wire N__10882;
    wire N__10881;
    wire N__10880;
    wire N__10873;
    wire N__10872;
    wire N__10871;
    wire N__10864;
    wire N__10863;
    wire N__10862;
    wire N__10855;
    wire N__10854;
    wire N__10853;
    wire N__10846;
    wire N__10845;
    wire N__10844;
    wire N__10837;
    wire N__10836;
    wire N__10835;
    wire N__10828;
    wire N__10827;
    wire N__10826;
    wire N__10819;
    wire N__10818;
    wire N__10817;
    wire N__10810;
    wire N__10809;
    wire N__10808;
    wire N__10801;
    wire N__10800;
    wire N__10799;
    wire N__10792;
    wire N__10791;
    wire N__10790;
    wire N__10783;
    wire N__10782;
    wire N__10781;
    wire N__10774;
    wire N__10773;
    wire N__10772;
    wire N__10765;
    wire N__10764;
    wire N__10763;
    wire N__10756;
    wire N__10755;
    wire N__10754;
    wire N__10747;
    wire N__10746;
    wire N__10745;
    wire N__10738;
    wire N__10737;
    wire N__10736;
    wire N__10729;
    wire N__10728;
    wire N__10727;
    wire N__10720;
    wire N__10719;
    wire N__10718;
    wire N__10711;
    wire N__10710;
    wire N__10709;
    wire N__10702;
    wire N__10701;
    wire N__10700;
    wire N__10693;
    wire N__10692;
    wire N__10691;
    wire N__10684;
    wire N__10683;
    wire N__10682;
    wire N__10675;
    wire N__10674;
    wire N__10673;
    wire N__10666;
    wire N__10665;
    wire N__10664;
    wire N__10657;
    wire N__10656;
    wire N__10655;
    wire N__10648;
    wire N__10647;
    wire N__10646;
    wire N__10639;
    wire N__10638;
    wire N__10637;
    wire N__10630;
    wire N__10629;
    wire N__10628;
    wire N__10621;
    wire N__10620;
    wire N__10619;
    wire N__10612;
    wire N__10611;
    wire N__10610;
    wire N__10603;
    wire N__10602;
    wire N__10601;
    wire N__10594;
    wire N__10593;
    wire N__10592;
    wire N__10585;
    wire N__10584;
    wire N__10583;
    wire N__10576;
    wire N__10575;
    wire N__10574;
    wire N__10567;
    wire N__10566;
    wire N__10565;
    wire N__10558;
    wire N__10557;
    wire N__10556;
    wire N__10549;
    wire N__10548;
    wire N__10547;
    wire N__10540;
    wire N__10539;
    wire N__10538;
    wire N__10531;
    wire N__10530;
    wire N__10529;
    wire N__10522;
    wire N__10521;
    wire N__10520;
    wire N__10513;
    wire N__10512;
    wire N__10511;
    wire N__10504;
    wire N__10503;
    wire N__10502;
    wire N__10495;
    wire N__10494;
    wire N__10493;
    wire N__10486;
    wire N__10485;
    wire N__10484;
    wire N__10477;
    wire N__10476;
    wire N__10475;
    wire N__10468;
    wire N__10467;
    wire N__10466;
    wire N__10459;
    wire N__10458;
    wire N__10457;
    wire N__10450;
    wire N__10449;
    wire N__10448;
    wire N__10441;
    wire N__10440;
    wire N__10439;
    wire N__10432;
    wire N__10431;
    wire N__10430;
    wire N__10413;
    wire N__10412;
    wire N__10411;
    wire N__10408;
    wire N__10405;
    wire N__10404;
    wire N__10401;
    wire N__10398;
    wire N__10395;
    wire N__10392;
    wire N__10389;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10359;
    wire N__10358;
    wire N__10357;
    wire N__10354;
    wire N__10353;
    wire N__10352;
    wire N__10351;
    wire N__10348;
    wire N__10347;
    wire N__10346;
    wire N__10343;
    wire N__10342;
    wire N__10341;
    wire N__10340;
    wire N__10339;
    wire N__10338;
    wire N__10335;
    wire N__10332;
    wire N__10329;
    wire N__10326;
    wire N__10323;
    wire N__10320;
    wire N__10317;
    wire N__10308;
    wire N__10305;
    wire N__10304;
    wire N__10303;
    wire N__10300;
    wire N__10299;
    wire N__10298;
    wire N__10297;
    wire N__10296;
    wire N__10295;
    wire N__10294;
    wire N__10285;
    wire N__10282;
    wire N__10273;
    wire N__10268;
    wire N__10265;
    wire N__10260;
    wire N__10257;
    wire N__10252;
    wire N__10249;
    wire N__10246;
    wire N__10239;
    wire N__10232;
    wire N__10227;
    wire N__10222;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10208;
    wire N__10205;
    wire N__10200;
    wire N__10199;
    wire N__10198;
    wire N__10195;
    wire N__10192;
    wire N__10189;
    wire N__10188;
    wire N__10183;
    wire N__10180;
    wire N__10177;
    wire N__10174;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10158;
    wire N__10155;
    wire N__10152;
    wire N__10151;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10136;
    wire N__10135;
    wire N__10134;
    wire N__10133;
    wire N__10132;
    wire N__10131;
    wire N__10130;
    wire N__10129;
    wire N__10128;
    wire N__10125;
    wire N__10104;
    wire N__10101;
    wire N__10098;
    wire N__10097;
    wire N__10094;
    wire N__10093;
    wire N__10092;
    wire N__10091;
    wire N__10090;
    wire N__10087;
    wire N__10086;
    wire N__10083;
    wire N__10080;
    wire N__10077;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10064;
    wire N__10059;
    wire N__10056;
    wire N__10053;
    wire N__10046;
    wire N__10043;
    wire N__10038;
    wire N__10035;
    wire N__10032;
    wire N__10029;
    wire N__10020;
    wire N__10019;
    wire N__10018;
    wire N__10017;
    wire N__10016;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__9998;
    wire N__9997;
    wire N__9996;
    wire N__9995;
    wire N__9994;
    wire N__9991;
    wire N__9990;
    wire N__9989;
    wire N__9988;
    wire N__9987;
    wire N__9986;
    wire N__9983;
    wire N__9982;
    wire N__9981;
    wire N__9980;
    wire N__9979;
    wire N__9978;
    wire N__9975;
    wire N__9974;
    wire N__9973;
    wire N__9972;
    wire N__9971;
    wire N__9970;
    wire N__9969;
    wire N__9968;
    wire N__9965;
    wire N__9964;
    wire N__9963;
    wire N__9962;
    wire N__9961;
    wire N__9960;
    wire N__9959;
    wire N__9958;
    wire N__9957;
    wire N__9956;
    wire N__9955;
    wire N__9954;
    wire N__9953;
    wire N__9952;
    wire N__9951;
    wire N__9950;
    wire N__9949;
    wire N__9948;
    wire N__9947;
    wire N__9946;
    wire N__9943;
    wire N__9852;
    wire N__9849;
    wire N__9846;
    wire N__9843;
    wire N__9840;
    wire N__9837;
    wire N__9834;
    wire N__9831;
    wire N__9830;
    wire N__9829;
    wire N__9828;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9809;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9792;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9780;
    wire N__9777;
    wire N__9774;
    wire N__9771;
    wire N__9768;
    wire N__9765;
    wire N__9764;
    wire N__9763;
    wire N__9762;
    wire N__9759;
    wire N__9756;
    wire N__9751;
    wire N__9746;
    wire N__9741;
    wire N__9738;
    wire N__9735;
    wire N__9732;
    wire N__9729;
    wire N__9726;
    wire N__9723;
    wire N__9722;
    wire N__9721;
    wire N__9720;
    wire N__9717;
    wire N__9714;
    wire N__9709;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9684;
    wire N__9681;
    wire N__9678;
    wire N__9675;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9663;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9651;
    wire N__9648;
    wire N__9645;
    wire N__9642;
    wire N__9639;
    wire N__9636;
    wire N__9633;
    wire N__9630;
    wire N__9629;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9619;
    wire N__9618;
    wire N__9615;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9603;
    wire N__9596;
    wire N__9593;
    wire N__9590;
    wire N__9585;
    wire N__9582;
    wire N__9579;
    wire N__9576;
    wire N__9575;
    wire N__9574;
    wire N__9571;
    wire N__9568;
    wire N__9565;
    wire N__9562;
    wire N__9557;
    wire N__9556;
    wire N__9553;
    wire N__9550;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9538;
    wire N__9531;
    wire N__9528;
    wire N__9525;
    wire N__9522;
    wire N__9519;
    wire N__9516;
    wire N__9515;
    wire N__9514;
    wire N__9509;
    wire N__9508;
    wire N__9505;
    wire N__9502;
    wire N__9499;
    wire N__9492;
    wire N__9489;
    wire N__9486;
    wire N__9483;
    wire N__9480;
    wire N__9477;
    wire N__9474;
    wire N__9473;
    wire N__9472;
    wire N__9469;
    wire N__9466;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9453;
    wire N__9450;
    wire N__9447;
    wire N__9442;
    wire N__9439;
    wire N__9436;
    wire N__9433;
    wire N__9430;
    wire N__9425;
    wire N__9420;
    wire N__9419;
    wire N__9414;
    wire N__9411;
    wire N__9408;
    wire N__9405;
    wire N__9402;
    wire N__9399;
    wire N__9396;
    wire N__9393;
    wire N__9390;
    wire N__9387;
    wire N__9384;
    wire N__9381;
    wire N__9378;
    wire N__9375;
    wire N__9372;
    wire N__9369;
    wire N__9366;
    wire N__9363;
    wire N__9360;
    wire N__9357;
    wire N__9354;
    wire N__9351;
    wire N__9348;
    wire N__9345;
    wire N__9342;
    wire N__9339;
    wire N__9336;
    wire N__9333;
    wire N__9330;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9309;
    wire N__9306;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9292;
    wire N__9291;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9264;
    wire N__9261;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9221;
    wire N__9220;
    wire N__9219;
    wire N__9218;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9206;
    wire N__9201;
    wire N__9192;
    wire N__9191;
    wire N__9190;
    wire N__9189;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9178;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9166;
    wire N__9163;
    wire N__9162;
    wire N__9159;
    wire N__9156;
    wire N__9153;
    wire N__9150;
    wire N__9147;
    wire N__9144;
    wire N__9139;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9114;
    wire N__9111;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9101;
    wire N__9100;
    wire N__9099;
    wire N__9098;
    wire N__9097;
    wire N__9096;
    wire N__9095;
    wire N__9094;
    wire N__9093;
    wire N__9092;
    wire N__9091;
    wire N__9090;
    wire N__9089;
    wire N__9088;
    wire N__9087;
    wire N__9086;
    wire N__9085;
    wire N__9084;
    wire N__9083;
    wire N__9082;
    wire N__9081;
    wire N__9080;
    wire N__9079;
    wire N__9078;
    wire N__9077;
    wire N__9076;
    wire N__9075;
    wire N__9072;
    wire N__9071;
    wire N__9070;
    wire N__9069;
    wire N__9068;
    wire N__9067;
    wire N__9066;
    wire N__8997;
    wire N__8994;
    wire N__8993;
    wire N__8990;
    wire N__8989;
    wire N__8988;
    wire N__8985;
    wire N__8984;
    wire N__8983;
    wire N__8980;
    wire N__8977;
    wire N__8974;
    wire N__8971;
    wire N__8968;
    wire N__8965;
    wire N__8952;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8937;
    wire N__8934;
    wire N__8931;
    wire N__8928;
    wire N__8925;
    wire N__8924;
    wire N__8923;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8894;
    wire N__8889;
    wire N__8886;
    wire N__8883;
    wire N__8882;
    wire N__8881;
    wire N__8880;
    wire N__8877;
    wire N__8874;
    wire N__8869;
    wire N__8868;
    wire N__8867;
    wire N__8866;
    wire N__8865;
    wire N__8864;
    wire N__8863;
    wire N__8862;
    wire N__8859;
    wire N__8856;
    wire N__8853;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8825;
    wire N__8822;
    wire N__8821;
    wire N__8818;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8808;
    wire N__8805;
    wire N__8802;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8790;
    wire N__8785;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8769;
    wire N__8766;
    wire N__8763;
    wire N__8762;
    wire N__8761;
    wire N__8758;
    wire N__8755;
    wire N__8752;
    wire N__8749;
    wire N__8746;
    wire N__8743;
    wire N__8740;
    wire N__8737;
    wire N__8734;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8709;
    wire N__8708;
    wire N__8707;
    wire N__8706;
    wire N__8705;
    wire N__8704;
    wire N__8703;
    wire N__8702;
    wire N__8701;
    wire N__8700;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8688;
    wire N__8685;
    wire N__8682;
    wire N__8681;
    wire N__8680;
    wire N__8677;
    wire N__8676;
    wire N__8675;
    wire N__8674;
    wire N__8671;
    wire N__8666;
    wire N__8663;
    wire N__8662;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8644;
    wire N__8641;
    wire N__8636;
    wire N__8633;
    wire N__8628;
    wire N__8625;
    wire N__8622;
    wire N__8617;
    wire N__8614;
    wire N__8611;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8595;
    wire N__8584;
    wire N__8579;
    wire N__8574;
    wire N__8571;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8544;
    wire N__8541;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8517;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8478;
    wire N__8475;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8463;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8455;
    wire N__8454;
    wire N__8453;
    wire N__8448;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8413;
    wire N__8408;
    wire N__8405;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8388;
    wire N__8385;
    wire N__8382;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8355;
    wire N__8352;
    wire N__8349;
    wire N__8346;
    wire N__8343;
    wire N__8340;
    wire N__8337;
    wire N__8334;
    wire N__8331;
    wire N__8328;
    wire N__8325;
    wire N__8322;
    wire N__8319;
    wire N__8316;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8306;
    wire N__8305;
    wire N__8304;
    wire N__8301;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8286;
    wire N__8283;
    wire N__8282;
    wire N__8279;
    wire N__8274;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8257;
    wire N__8250;
    wire N__8247;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8239;
    wire N__8238;
    wire N__8237;
    wire N__8232;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8221;
    wire N__8220;
    wire N__8219;
    wire N__8216;
    wire N__8213;
    wire N__8208;
    wire N__8207;
    wire N__8206;
    wire N__8205;
    wire N__8204;
    wire N__8203;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8193;
    wire N__8192;
    wire N__8191;
    wire N__8188;
    wire N__8187;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8169;
    wire N__8166;
    wire N__8165;
    wire N__8164;
    wire N__8163;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8151;
    wire N__8148;
    wire N__8141;
    wire N__8140;
    wire N__8137;
    wire N__8132;
    wire N__8127;
    wire N__8118;
    wire N__8107;
    wire N__8104;
    wire N__8091;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8080;
    wire N__8075;
    wire N__8072;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8062;
    wire N__8055;
    wire N__8052;
    wire N__8049;
    wire N__8048;
    wire N__8047;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8035;
    wire N__8034;
    wire N__8029;
    wire N__8028;
    wire N__8025;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8013;
    wire N__8010;
    wire N__8001;
    wire N__7998;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7971;
    wire N__7970;
    wire N__7969;
    wire N__7966;
    wire N__7961;
    wire N__7956;
    wire N__7955;
    wire N__7950;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7931;
    wire N__7930;
    wire N__7927;
    wire N__7926;
    wire N__7925;
    wire N__7924;
    wire N__7923;
    wire N__7922;
    wire N__7921;
    wire N__7920;
    wire N__7919;
    wire N__7916;
    wire N__7915;
    wire N__7914;
    wire N__7913;
    wire N__7906;
    wire N__7903;
    wire N__7902;
    wire N__7899;
    wire N__7896;
    wire N__7893;
    wire N__7890;
    wire N__7889;
    wire N__7888;
    wire N__7885;
    wire N__7882;
    wire N__7881;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7869;
    wire N__7864;
    wire N__7861;
    wire N__7858;
    wire N__7857;
    wire N__7856;
    wire N__7849;
    wire N__7846;
    wire N__7845;
    wire N__7844;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7830;
    wire N__7825;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7813;
    wire N__7808;
    wire N__7803;
    wire N__7798;
    wire N__7793;
    wire N__7784;
    wire N__7767;
    wire N__7764;
    wire N__7761;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7751;
    wire N__7748;
    wire N__7745;
    wire N__7740;
    wire N__7737;
    wire N__7734;
    wire N__7733;
    wire N__7730;
    wire N__7727;
    wire N__7722;
    wire N__7719;
    wire N__7718;
    wire N__7715;
    wire N__7712;
    wire N__7707;
    wire N__7704;
    wire N__7701;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7686;
    wire N__7683;
    wire N__7682;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7668;
    wire N__7665;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7653;
    wire N__7650;
    wire N__7647;
    wire N__7644;
    wire N__7641;
    wire N__7638;
    wire N__7635;
    wire N__7632;
    wire N__7629;
    wire N__7626;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7602;
    wire N__7599;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7581;
    wire N__7578;
    wire N__7575;
    wire N__7572;
    wire N__7569;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7551;
    wire N__7548;
    wire N__7545;
    wire N__7542;
    wire N__7539;
    wire N__7536;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7485;
    wire N__7482;
    wire N__7479;
    wire N__7476;
    wire N__7473;
    wire N__7470;
    wire N__7467;
    wire N__7464;
    wire N__7461;
    wire N__7458;
    wire N__7455;
    wire N__7452;
    wire N__7449;
    wire N__7446;
    wire N__7443;
    wire N__7440;
    wire N__7437;
    wire N__7434;
    wire N__7431;
    wire N__7428;
    wire N__7425;
    wire N__7422;
    wire N__7419;
    wire N__7416;
    wire N__7413;
    wire N__7410;
    wire N__7407;
    wire N__7404;
    wire N__7401;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7389;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7374;
    wire N__7371;
    wire N__7368;
    wire N__7365;
    wire N__7362;
    wire N__7359;
    wire N__7356;
    wire N__7353;
    wire N__7350;
    wire N__7347;
    wire N__7344;
    wire N__7341;
    wire N__7338;
    wire N__7335;
    wire N__7332;
    wire N__7329;
    wire N__7326;
    wire N__7323;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7311;
    wire N__7308;
    wire N__7305;
    wire N__7302;
    wire N__7299;
    wire N__7296;
    wire N__7293;
    wire N__7290;
    wire N__7287;
    wire N__7286;
    wire N__7285;
    wire N__7284;
    wire N__7281;
    wire N__7276;
    wire N__7275;
    wire N__7272;
    wire N__7269;
    wire N__7266;
    wire N__7263;
    wire N__7254;
    wire N__7253;
    wire N__7252;
    wire N__7251;
    wire N__7250;
    wire N__7247;
    wire N__7246;
    wire N__7245;
    wire N__7244;
    wire N__7243;
    wire N__7240;
    wire N__7239;
    wire N__7238;
    wire N__7237;
    wire N__7234;
    wire N__7231;
    wire N__7230;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7218;
    wire N__7217;
    wire N__7216;
    wire N__7209;
    wire N__7204;
    wire N__7197;
    wire N__7194;
    wire N__7191;
    wire N__7184;
    wire N__7181;
    wire N__7180;
    wire N__7179;
    wire N__7178;
    wire N__7177;
    wire N__7174;
    wire N__7169;
    wire N__7164;
    wire N__7157;
    wire N__7154;
    wire N__7149;
    wire N__7146;
    wire N__7131;
    wire N__7130;
    wire N__7129;
    wire N__7128;
    wire N__7125;
    wire N__7122;
    wire N__7119;
    wire N__7116;
    wire N__7115;
    wire N__7114;
    wire N__7113;
    wire N__7112;
    wire N__7109;
    wire N__7104;
    wire N__7101;
    wire N__7098;
    wire N__7097;
    wire N__7092;
    wire N__7089;
    wire N__7086;
    wire N__7083;
    wire N__7078;
    wire N__7075;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7049;
    wire N__7048;
    wire N__7045;
    wire N__7044;
    wire N__7043;
    wire N__7042;
    wire N__7041;
    wire N__7040;
    wire N__7039;
    wire N__7038;
    wire N__7035;
    wire N__7032;
    wire N__7031;
    wire N__7030;
    wire N__7029;
    wire N__7026;
    wire N__7025;
    wire N__7022;
    wire N__7021;
    wire N__7010;
    wire N__7009;
    wire N__7008;
    wire N__7005;
    wire N__7000;
    wire N__6997;
    wire N__6992;
    wire N__6991;
    wire N__6990;
    wire N__6987;
    wire N__6984;
    wire N__6981;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6960;
    wire N__6955;
    wire N__6950;
    wire N__6933;
    wire N__6932;
    wire N__6931;
    wire N__6930;
    wire N__6929;
    wire N__6926;
    wire N__6925;
    wire N__6924;
    wire N__6921;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6913;
    wire N__6912;
    wire N__6911;
    wire N__6910;
    wire N__6907;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6885;
    wire N__6884;
    wire N__6881;
    wire N__6880;
    wire N__6877;
    wire N__6874;
    wire N__6869;
    wire N__6858;
    wire N__6853;
    wire N__6848;
    wire N__6837;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6819;
    wire N__6816;
    wire N__6813;
    wire N__6810;
    wire N__6807;
    wire N__6804;
    wire N__6801;
    wire N__6798;
    wire N__6795;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6783;
    wire N__6782;
    wire N__6781;
    wire N__6780;
    wire N__6777;
    wire N__6770;
    wire N__6765;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6757;
    wire N__6756;
    wire N__6755;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6745;
    wire N__6742;
    wire N__6739;
    wire N__6736;
    wire N__6727;
    wire N__6724;
    wire N__6723;
    wire N__6720;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6702;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6688;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6676;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6660;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6650;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6639;
    wire N__6632;
    wire N__6629;
    wire N__6626;
    wire N__6623;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6606;
    wire N__6603;
    wire N__6600;
    wire N__6597;
    wire N__6594;
    wire N__6591;
    wire N__6588;
    wire N__6585;
    wire N__6582;
    wire N__6579;
    wire N__6576;
    wire N__6573;
    wire N__6570;
    wire N__6567;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6555;
    wire N__6552;
    wire N__6549;
    wire N__6546;
    wire N__6543;
    wire N__6540;
    wire N__6537;
    wire N__6534;
    wire N__6531;
    wire N__6528;
    wire N__6525;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6501;
    wire N__6498;
    wire N__6495;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6483;
    wire N__6480;
    wire N__6477;
    wire N__6474;
    wire N__6471;
    wire N__6468;
    wire N__6465;
    wire N__6462;
    wire N__6461;
    wire N__6458;
    wire N__6455;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6441;
    wire N__6440;
    wire N__6437;
    wire N__6434;
    wire N__6429;
    wire N__6426;
    wire N__6425;
    wire N__6422;
    wire N__6419;
    wire N__6418;
    wire N__6413;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6399;
    wire N__6396;
    wire N__6395;
    wire N__6392;
    wire N__6391;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6379;
    wire N__6372;
    wire N__6369;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6359;
    wire N__6354;
    wire N__6351;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6336;
    wire N__6335;
    wire N__6330;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6315;
    wire N__6312;
    wire N__6309;
    wire N__6306;
    wire N__6303;
    wire N__6300;
    wire N__6297;
    wire N__6294;
    wire N__6291;
    wire N__6288;
    wire N__6285;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6255;
    wire N__6254;
    wire N__6253;
    wire N__6252;
    wire N__6249;
    wire N__6246;
    wire N__6245;
    wire N__6242;
    wire N__6241;
    wire N__6240;
    wire N__6239;
    wire N__6238;
    wire N__6235;
    wire N__6226;
    wire N__6221;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6202;
    wire N__6201;
    wire N__6200;
    wire N__6197;
    wire N__6188;
    wire N__6181;
    wire N__6174;
    wire N__6171;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6163;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6147;
    wire N__6144;
    wire N__6141;
    wire N__6140;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6129;
    wire N__6128;
    wire N__6127;
    wire N__6126;
    wire N__6125;
    wire N__6122;
    wire N__6121;
    wire N__6120;
    wire N__6119;
    wire N__6118;
    wire N__6117;
    wire N__6116;
    wire N__6111;
    wire N__6108;
    wire N__6107;
    wire N__6104;
    wire N__6099;
    wire N__6096;
    wire N__6093;
    wire N__6090;
    wire N__6083;
    wire N__6082;
    wire N__6081;
    wire N__6078;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6065;
    wire N__6060;
    wire N__6055;
    wire N__6050;
    wire N__6047;
    wire N__6044;
    wire N__6039;
    wire N__6018;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5985;
    wire N__5982;
    wire N__5979;
    wire N__5978;
    wire N__5977;
    wire N__5972;
    wire N__5969;
    wire N__5964;
    wire N__5963;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5946;
    wire N__5943;
    wire N__5942;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5925;
    wire N__5922;
    wire N__5921;
    wire N__5918;
    wire N__5915;
    wire N__5910;
    wire N__5907;
    wire N__5904;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5894;
    wire N__5891;
    wire N__5888;
    wire N__5883;
    wire N__5880;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5862;
    wire N__5859;
    wire N__5856;
    wire N__5853;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5829;
    wire N__5828;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5811;
    wire N__5810;
    wire N__5809;
    wire N__5806;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5793;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5766;
    wire N__5763;
    wire N__5762;
    wire N__5761;
    wire N__5760;
    wire N__5759;
    wire N__5758;
    wire N__5757;
    wire N__5756;
    wire N__5751;
    wire N__5746;
    wire N__5745;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5737;
    wire N__5734;
    wire N__5733;
    wire N__5730;
    wire N__5725;
    wire N__5720;
    wire N__5715;
    wire N__5712;
    wire N__5709;
    wire N__5706;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5682;
    wire N__5681;
    wire N__5678;
    wire N__5677;
    wire N__5676;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5662;
    wire N__5659;
    wire N__5652;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5633;
    wire N__5630;
    wire N__5625;
    wire N__5622;
    wire N__5619;
    wire N__5616;
    wire N__5613;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5598;
    wire N__5595;
    wire N__5592;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5577;
    wire N__5576;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5565;
    wire N__5560;
    wire N__5559;
    wire N__5554;
    wire N__5551;
    wire N__5548;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5532;
    wire N__5531;
    wire N__5530;
    wire N__5529;
    wire N__5528;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5511;
    wire N__5502;
    wire N__5499;
    wire N__5496;
    wire N__5493;
    wire N__5490;
    wire N__5487;
    wire N__5484;
    wire N__5481;
    wire N__5478;
    wire N__5475;
    wire N__5472;
    wire N__5469;
    wire N__5466;
    wire N__5465;
    wire N__5462;
    wire N__5459;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5448;
    wire N__5445;
    wire N__5440;
    wire N__5437;
    wire N__5436;
    wire N__5433;
    wire N__5428;
    wire N__5425;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5409;
    wire N__5408;
    wire N__5407;
    wire N__5404;
    wire N__5401;
    wire N__5398;
    wire N__5391;
    wire N__5388;
    wire N__5385;
    wire N__5382;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5345;
    wire N__5342;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5325;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5307;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5285;
    wire N__5282;
    wire N__5277;
    wire N__5274;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5262;
    wire N__5259;
    wire N__5256;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5205;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5187;
    wire N__5184;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5166;
    wire N__5165;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5148;
    wire N__5145;
    wire N__5142;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5130;
    wire N__5127;
    wire N__5124;
    wire N__5121;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5091;
    wire N__5088;
    wire N__5087;
    wire N__5086;
    wire N__5085;
    wire N__5084;
    wire N__5081;
    wire N__5080;
    wire N__5079;
    wire N__5070;
    wire N__5067;
    wire N__5062;
    wire N__5059;
    wire N__5052;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire N__5040;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5004;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4977;
    wire N__4976;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4963;
    wire N__4960;
    wire N__4957;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4872;
    wire N__4869;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4857;
    wire N__4854;
    wire N__4851;
    wire N__4848;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4836;
    wire N__4835;
    wire N__4834;
    wire N__4831;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4809;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4781;
    wire N__4780;
    wire N__4777;
    wire N__4774;
    wire N__4771;
    wire N__4764;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4743;
    wire N__4742;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4725;
    wire N__4722;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4704;
    wire N__4701;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4691;
    wire N__4686;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4674;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4662;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4647;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4593;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4575;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4545;
    wire N__4542;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4530;
    wire N__4527;
    wire N__4524;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4512;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4500;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4488;
    wire N__4485;
    wire N__4482;
    wire N__4479;
    wire N__4478;
    wire N__4477;
    wire N__4474;
    wire N__4469;
    wire N__4468;
    wire N__4467;
    wire N__4466;
    wire N__4465;
    wire N__4460;
    wire N__4451;
    wire N__4446;
    wire N__4445;
    wire N__4444;
    wire N__4443;
    wire N__4438;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4415;
    wire N__4414;
    wire N__4413;
    wire N__4410;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4383;
    wire N__4382;
    wire N__4381;
    wire N__4380;
    wire N__4377;
    wire N__4376;
    wire N__4375;
    wire N__4374;
    wire N__4371;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4356;
    wire N__4349;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4313;
    wire N__4312;
    wire N__4311;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4293;
    wire N__4284;
    wire N__4283;
    wire N__4280;
    wire N__4279;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4267;
    wire N__4260;
    wire N__4257;
    wire N__4256;
    wire N__4255;
    wire N__4254;
    wire N__4253;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4212;
    wire N__4209;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4197;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4178;
    wire N__4177;
    wire N__4176;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4136;
    wire N__4133;
    wire N__4130;
    wire N__4125;
    wire N__4124;
    wire N__4123;
    wire N__4122;
    wire N__4121;
    wire N__4120;
    wire N__4115;
    wire N__4110;
    wire N__4105;
    wire N__4098;
    wire N__4095;
    wire N__4092;
    wire N__4091;
    wire N__4088;
    wire N__4087;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4075;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4059;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4038;
    wire N__4037;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4023;
    wire N__4020;
    wire N__4017;
    wire N__4014;
    wire N__4011;
    wire N__4008;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3957;
    wire N__3954;
    wire N__3953;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3941;
    wire N__3938;
    wire N__3935;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3900;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3885;
    wire N__3882;
    wire N__3879;
    wire N__3876;
    wire N__3873;
    wire N__3870;
    wire N__3867;
    wire N__3864;
    wire N__3861;
    wire N__3858;
    wire N__3855;
    wire N__3852;
    wire N__3849;
    wire N__3846;
    wire N__3843;
    wire N__3840;
    wire N__3837;
    wire N__3834;
    wire N__3831;
    wire N__3828;
    wire N__3827;
    wire N__3824;
    wire N__3821;
    wire N__3816;
    wire N__3813;
    wire N__3812;
    wire N__3809;
    wire N__3806;
    wire N__3801;
    wire N__3800;
    wire N__3797;
    wire N__3794;
    wire N__3789;
    wire N__3788;
    wire N__3785;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3759;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire N_991_i;
    wire CLK80_PLL_i_i;
    wire ASn_c;
    wire \U712_REG_SM.N_238_cascade_ ;
    wire \U712_REG_SM.N_238 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire \U712_REG_SM.ASn_0_sqmuxa_1 ;
    wire \U712_REG_SM.N_219_cascade_ ;
    wire \U712_REG_SM.N_304 ;
    wire \U712_REG_SM.N_304_cascade_ ;
    wire \U712_REG_SM.STATE_COUNT_srsts_i_0_i_0_1 ;
    wire C3_c;
    wire C1_c;
    wire REGSPACEn_c;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire REGENn_c;
    wire \U712_REG_SM.N_307 ;
    wire \U712_REG_SM.N_219 ;
    wire \U712_REG_SM.REG_TACK_RNOZ0Z_0 ;
    wire \U712_REG_SM.N_235 ;
    wire \U712_CHIP_RAM.un5_DMA_CYCLE_START_0_cascade_ ;
    wire \U712_REG_SM.N_225 ;
    wire \U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_1_1_3_cascade_ ;
    wire \U712_REG_SM.N_259 ;
    wire \U712_REG_SM.N_259_cascade_ ;
    wire \U712_REG_SM.N_236 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.STATE_COUNT_srsts_i_i_0_0_3 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire N_40_i;
    wire \U712_REG_SM.N_261 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire N_41_i;
    wire \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_0 ;
    wire \U712_REG_SM.DS_EN_RNOZ0Z_0 ;
    wire \U712_REG_SM.N_314 ;
    wire REG_TACK;
    wire \U712_CYCLE_TERM.TACK_EN6_0_cascade_ ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_2 ;
    wire TACK_OUTn;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire bfn_7_9_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.N_282_cascade_ ;
    wire \U712_CHIP_RAM.N_265_cascade_ ;
    wire \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_i_2_cascade_ ;
    wire CPU_TACKm;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.N_218 ;
    wire \U712_CHIP_RAM.N_208_cascade_ ;
    wire \U712_CHIP_RAM.N_245_cascade_ ;
    wire \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a3_0_2 ;
    wire A_c_4;
    wire A_c_11;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ;
    wire \U712_BYTE_ENABLE.N_327 ;
    wire CASUn_c;
    wire \U712_BYTE_ENABLE.N_319_cascade_ ;
    wire N_43_i;
    wire SIZ_c_1;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0 ;
    wire \U712_BYTE_ENABLE.N_321 ;
    wire A_c_1;
    wire \U712_BYTE_ENABLE.un1_CLMBEn_i_0Z0Z_0 ;
    wire TACK_EN_i_ess;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.N_233_i_0_en_cascade_ ;
    wire \U712_CYCLE_TERM.N_233_i_0_en_0 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ;
    wire VBENn_c;
    wire \U712_CHIP_RAM.N_209_cascade_ ;
    wire \U712_CHIP_RAM.N_359_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0_cascade_ ;
    wire \U712_CHIP_RAM.N_290_cascade_ ;
    wire \U712_CHIP_RAM.N_181_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_a4_0_a3_0 ;
    wire \U712_CHIP_RAM.N_216_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.N_181 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.N_204_cascade_ ;
    wire \U712_CHIP_RAM.N_279_1 ;
    wire \U712_CHIP_RAM.N_279_1_cascade_ ;
    wire \U712_CHIP_RAM.N_398 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_393 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0 ;
    wire \U712_CHIP_RAM.REFRESH_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.N_227_cascade_ ;
    wire \U712_CHIP_RAM.N_226 ;
    wire \U712_CHIP_RAM.N_245 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ;
    wire DBENn_c;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0 ;
    wire \U712_BYTE_ENABLE.N_319 ;
    wire \U712_BYTE_ENABLE.N_322 ;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_cascade_ ;
    wire CASLn_c;
    wire N_42_i;
    wire REG_CYCLEm;
    wire DRDENn_c;
    wire A_c_8;
    wire A_c_15;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0 ;
    wire A_c_6;
    wire A_c_13;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ;
    wire \U712_CHIP_RAM.N_257 ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_205 ;
    wire \U712_CHIP_RAM.N_205_cascade_ ;
    wire \U712_CHIP_RAM.N_216 ;
    wire \U712_CHIP_RAM.N_291 ;
    wire \U712_CHIP_RAM.N_291_cascade_ ;
    wire \U712_CHIP_RAM.N_204 ;
    wire \U712_CHIP_RAM.N_342_cascade_ ;
    wire A_c_20;
    wire \U712_CHIP_RAM.N_352_cascade_ ;
    wire \U712_CHIP_RAM.N_395 ;
    wire \U712_CHIP_RAM.N_352 ;
    wire \U712_CHIP_RAM.N_293_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_99_cascade_ ;
    wire \U712_CHIP_RAM.N_290 ;
    wire BANK0_c;
    wire TSn_c;
    wire RAMSPACEn_c;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_359 ;
    wire DBDIR_c;
    wire DBR_SYNCZ0Z_0;
    wire DBR_SYNCZ0Z_1;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire RAS1n_c;
    wire \U712_CHIP_RAM.REFRESH_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0 ;
    wire \U712_CHIP_RAM.N_301 ;
    wire \U712_CHIP_RAM.N_243 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_209 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.N_227 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_2 ;
    wire \U712_CHIP_RAM.N_303 ;
    wire \U712_CHIP_RAM.N_241 ;
    wire DMA_CYCLEm;
    wire AWEn_c;
    wire RnW_c;
    wire N_256;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire CONSTANT_ONE_NET;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire CMA_c_4;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire A_c_7;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ;
    wire \U712_CHIP_RAM.N_289 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.N_342 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.N_208 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_a3_0 ;
    wire A_c_16;
    wire A_c_18;
    wire A_c_10;
    wire A_c_3;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ;
    wire A_c_12;
    wire A_c_5;
    wire A_c_2;
    wire A_c_9;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire A_c_17;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.un1_CMA28_0_i ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CMA_c_2;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire A_c_14;
    wire CPU_CYCLEm;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_11_11_0_;
    wire \U712_CHIP_RAM.REFRESH5lto1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH5lto2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire un1_LDSn_i_0_0;
    wire DS_ENm;
    wire A_c_0;
    wire SIZ_c_0;
    wire un1_UDSn_i_0_0;
    wire RASn_c;
    wire CRCSn_c;
    wire WEn_c;
    wire CASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire CMA_c_10;
    wire RAS0n_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire CLK80_PLL;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire \U712_CHIP_RAM.DMA_AZ0Z20 ;
    wire \INVU712_CHIP_RAM.DMA_A20C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10_cascade_ ;
    wire DBRn_c;
    wire C1_c_g;
    wire CLK40_PLL_i;
    wire CLK40_PLL_i_i;
    wire RESETn_c;
    wire RESETn_c_i;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire DRA_c_9;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire DRA_c_2;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire DRA_c_6;
    wire AGNUS_REV_c;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire _gnd_net_;
    wire C3_c_g;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ;
    wire RESETn_c_i_g;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__3777),
            .RESETB(N__6582),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__11197),
            .DIN(N__11196),
            .DOUT(N__11195),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__11197),
            .PADOUT(N__11196),
            .PADIN(N__11195),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5469),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11188),
            .DIN(N__11187),
            .DOUT(N__11186),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11188),
            .PADOUT(N__11187),
            .PADIN(N__11186),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__11179),
            .DIN(N__11178),
            .DOUT(N__11177),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__11179),
            .PADOUT(N__11178),
            .PADIN(N__11177),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8322),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__11170),
            .DIN(N__11169),
            .DOUT(N__11168),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__11170),
            .PADOUT(N__11169),
            .PADIN(N__11168),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6609),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__11161),
            .DIN(N__11160),
            .DOUT(N__11159),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__11161),
            .PADOUT(N__11160),
            .PADIN(N__11159),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__11152),
            .DIN(N__11151),
            .DOUT(N__11150),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__11152),
            .PADOUT(N__11151),
            .PADIN(N__11150),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__11143),
            .DIN(N__11142),
            .DOUT(N__11141),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__11143),
            .PADOUT(N__11142),
            .PADIN(N__11141),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__11134),
            .DIN(N__11133),
            .DOUT(N__11132),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__11134),
            .PADOUT(N__11133),
            .PADIN(N__11132),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__11125),
            .DIN(N__11124),
            .DOUT(N__11123),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__11125),
            .PADOUT(N__11124),
            .PADIN(N__11123),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__11116),
            .DIN(N__11115),
            .DOUT(N__11114),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__11116),
            .PADOUT(N__11115),
            .PADIN(N__11114),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11107),
            .DIN(N__11106),
            .DOUT(N__11105),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11107),
            .PADOUT(N__11106),
            .PADIN(N__11105),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__11098),
            .DIN(N__11097),
            .DOUT(N__11096),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__11098),
            .PADOUT(N__11097),
            .PADIN(N__11096),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7620),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__11089),
            .DIN(N__11088),
            .DOUT(N__11087),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__11089),
            .PADOUT(N__11088),
            .PADIN(N__11087),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__11080),
            .DIN(N__11079),
            .DOUT(N__11078),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__11080),
            .PADOUT(N__11079),
            .PADIN(N__11078),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__11071),
            .DIN(N__11070),
            .DOUT(N__11069),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__11071),
            .PADOUT(N__11070),
            .PADIN(N__11069),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__11062),
            .DIN(N__11061),
            .DOUT(N__11060),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__11062),
            .PADOUT(N__11061),
            .PADIN(N__11060),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5001),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__11053),
            .DIN(N__11052),
            .DOUT(N__11051),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__11053),
            .PADOUT(N__11052),
            .PADIN(N__11051),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11044),
            .DIN(N__11043),
            .DOUT(N__11042),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11044),
            .PADOUT(N__11043),
            .PADIN(N__11042),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__11035),
            .DIN(N__11034),
            .DOUT(N__11033),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__11035),
            .PADOUT(N__11034),
            .PADIN(N__11033),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7353),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__11026),
            .DIN(N__11025),
            .DOUT(N__11024),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__11026),
            .PADOUT(N__11025),
            .PADIN(N__11024),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__11017),
            .DIN(N__11016),
            .DOUT(N__11015),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__11017),
            .PADOUT(N__11016),
            .PADIN(N__11015),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8355),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11008),
            .DIN(N__11007),
            .DOUT(N__11006),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11008),
            .PADOUT(N__11007),
            .PADIN(N__11006),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__10999),
            .DIN(N__10998),
            .DOUT(N__10997),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__10999),
            .PADOUT(N__10998),
            .PADIN(N__10997),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__10990),
            .DIN(N__10989),
            .DOUT(N__10988),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__10990),
            .PADOUT(N__10989),
            .PADIN(N__10988),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__10981),
            .DIN(N__10980),
            .DOUT(N__10979),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__10981),
            .PADOUT(N__10980),
            .PADIN(N__10979),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__10972),
            .DIN(N__10971),
            .DOUT(N__10970),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__10972),
            .PADOUT(N__10971),
            .PADIN(N__10970),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__10963),
            .DIN(N__10962),
            .DOUT(N__10961),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__10963),
            .PADOUT(N__10962),
            .PADIN(N__10961),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__10954),
            .DIN(N__10953),
            .DOUT(N__10952),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__10954),
            .PADOUT(N__10953),
            .PADIN(N__10952),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__10945),
            .DIN(N__10944),
            .DOUT(N__10943),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__10945),
            .PADOUT(N__10944),
            .PADIN(N__10943),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__10936),
            .DIN(N__10935),
            .DOUT(N__10934),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__10936),
            .PADOUT(N__10935),
            .PADIN(N__10934),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7368),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__10927),
            .DIN(N__10926),
            .DOUT(N__10925),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__10927),
            .PADOUT(N__10926),
            .PADIN(N__10925),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__10918),
            .DIN(N__10917),
            .DOUT(N__10916),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__10918),
            .PADOUT(N__10917),
            .PADIN(N__10916),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__10909),
            .DIN(N__10908),
            .DOUT(N__10907),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__10909),
            .PADOUT(N__10908),
            .PADIN(N__10907),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__10900),
            .DIN(N__10899),
            .DOUT(N__10898),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__10900),
            .PADOUT(N__10899),
            .PADIN(N__10898),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__10891),
            .DIN(N__10890),
            .DOUT(N__10889),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__10891),
            .PADOUT(N__10890),
            .PADIN(N__10889),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__10882),
            .DIN(N__10881),
            .DOUT(N__10880),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__10882),
            .PADOUT(N__10881),
            .PADIN(N__10880),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8508),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__10873),
            .DIN(N__10872),
            .DOUT(N__10871),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__10873),
            .PADOUT(N__10872),
            .PADIN(N__10871),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8766),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__10864),
            .DIN(N__10863),
            .DOUT(N__10862),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__10864),
            .PADOUT(N__10863),
            .PADIN(N__10862),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__10855),
            .DIN(N__10854),
            .DOUT(N__10853),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__10855),
            .PADOUT(N__10854),
            .PADIN(N__10853),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8376),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__10846),
            .DIN(N__10845),
            .DOUT(N__10844),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__10846),
            .PADOUT(N__10845),
            .PADIN(N__10844),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__10837),
            .DIN(N__10836),
            .DOUT(N__10835),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__10837),
            .PADOUT(N__10836),
            .PADIN(N__10835),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5910),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__10828),
            .DIN(N__10827),
            .DOUT(N__10826),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__10828),
            .PADOUT(N__10827),
            .PADIN(N__10826),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8762),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__10819),
            .DIN(N__10818),
            .DOUT(N__10817),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__10819),
            .PADOUT(N__10818),
            .PADIN(N__10817),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3867),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__10810),
            .DIN(N__10809),
            .DOUT(N__10808),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__10810),
            .PADOUT(N__10809),
            .PADIN(N__10808),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__10801),
            .DIN(N__10800),
            .DOUT(N__10799),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__10801),
            .PADOUT(N__10800),
            .PADIN(N__10799),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3849),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__10792),
            .DIN(N__10791),
            .DOUT(N__10790),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__10792),
            .PADOUT(N__10791),
            .PADIN(N__10790),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9120),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__10783),
            .DIN(N__10782),
            .DOUT(N__10781),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__10783),
            .PADOUT(N__10782),
            .PADIN(N__10781),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__10774),
            .DIN(N__10773),
            .DOUT(N__10772),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__10774),
            .PADOUT(N__10773),
            .PADIN(N__10772),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__10765),
            .DIN(N__10764),
            .DOUT(N__10763),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__10765),
            .PADOUT(N__10764),
            .PADIN(N__10763),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_0_iopad (
            .OE(N__10756),
            .DIN(N__10755),
            .DOUT(N__10754),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__10756),
            .PADOUT(N__10755),
            .PADIN(N__10754),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__10747),
            .DIN(N__10746),
            .DOUT(N__10745),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__10747),
            .PADOUT(N__10746),
            .PADIN(N__10745),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8001),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__10738),
            .DIN(N__10737),
            .DOUT(N__10736),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__10738),
            .PADOUT(N__10737),
            .PADIN(N__10736),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__10729),
            .DIN(N__10728),
            .DOUT(N__10727),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__10729),
            .PADOUT(N__10728),
            .PADIN(N__10727),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8761),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__10720),
            .DIN(N__10719),
            .DOUT(N__10718),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__10720),
            .PADOUT(N__10719),
            .PADIN(N__10718),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6507),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__10711),
            .DIN(N__10710),
            .DOUT(N__10709),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__10711),
            .PADOUT(N__10710),
            .PADIN(N__10709),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5277),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__10702),
            .DIN(N__10701),
            .DOUT(N__10700),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__10702),
            .PADOUT(N__10701),
            .PADIN(N__10700),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4338),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__10693),
            .DIN(N__10692),
            .DOUT(N__10691),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__10693),
            .PADOUT(N__10692),
            .PADIN(N__10691),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6537),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__10684),
            .DIN(N__10683),
            .DOUT(N__10682),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__10684),
            .PADOUT(N__10683),
            .PADIN(N__10682),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4098),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__10675),
            .DIN(N__10674),
            .DOUT(N__10673),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__10675),
            .PADOUT(N__10674),
            .PADIN(N__10673),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__10666),
            .DIN(N__10665),
            .DOUT(N__10664),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__10666),
            .PADOUT(N__10665),
            .PADIN(N__10664),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__10657),
            .DIN(N__10656),
            .DOUT(N__10655),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__10657),
            .PADOUT(N__10656),
            .PADIN(N__10655),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4221),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__10648),
            .DIN(N__10647),
            .DOUT(N__10646),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__10648),
            .PADOUT(N__10647),
            .PADIN(N__10646),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8337),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__10639),
            .DIN(N__10638),
            .DOUT(N__10637),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__10639),
            .PADOUT(N__10638),
            .PADIN(N__10637),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5652),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__10630),
            .DIN(N__10629),
            .DOUT(N__10628),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__10630),
            .PADOUT(N__10629),
            .PADIN(N__10628),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5337),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_obuf_iopad (
            .OE(N__10621),
            .DIN(N__10620),
            .DOUT(N__10619),
            .PACKAGEPIN(DMA_LATCH));
    defparam DMA_LATCH_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_obuf_preio (
            .PADOEN(N__10621),
            .PADOUT(N__10620),
            .PADIN(N__10619),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__10612),
            .DIN(N__10611),
            .DOUT(N__10610),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__10612),
            .PADOUT(N__10611),
            .PADIN(N__10610),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__10603),
            .DIN(N__10602),
            .DOUT(N__10601),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__10603),
            .PADOUT(N__10602),
            .PADIN(N__10601),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__10594),
            .DIN(N__10593),
            .DOUT(N__10592),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__10594),
            .PADOUT(N__10593),
            .PADIN(N__10592),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__10585),
            .DIN(N__10584),
            .DOUT(N__10583),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__10585),
            .PADOUT(N__10584),
            .PADIN(N__10583),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__10576),
            .DIN(N__10575),
            .DOUT(N__10574),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__10576),
            .PADOUT(N__10575),
            .PADIN(N__10574),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6492),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__10567),
            .DIN(N__10566),
            .DOUT(N__10565),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__10567),
            .PADOUT(N__10566),
            .PADIN(N__10565),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__10558),
            .DIN(N__10557),
            .DOUT(N__10556),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__10558),
            .PADOUT(N__10557),
            .PADIN(N__10556),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4929),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__10549),
            .DIN(N__10548),
            .DOUT(N__10547),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__10549),
            .PADOUT(N__10548),
            .PADIN(N__10547),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3885),
            .DIN0(),
            .DOUT0(N__4536),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__10540),
            .DIN(N__10539),
            .DOUT(N__10538),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__10540),
            .PADOUT(N__10539),
            .PADIN(N__10538),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7632),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__10531),
            .DIN(N__10530),
            .DOUT(N__10529),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__10531),
            .PADOUT(N__10530),
            .PADIN(N__10529),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__10522),
            .DIN(N__10521),
            .DOUT(N__10520),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__10522),
            .PADOUT(N__10521),
            .PADIN(N__10520),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__10513),
            .DIN(N__10512),
            .DOUT(N__10511),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__10513),
            .PADOUT(N__10512),
            .PADIN(N__10511),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7398),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__10504),
            .DIN(N__10503),
            .DOUT(N__10502),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__10504),
            .PADOUT(N__10503),
            .PADIN(N__10502),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__10495),
            .DIN(N__10494),
            .DOUT(N__10493),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__10495),
            .PADOUT(N__10494),
            .PADIN(N__10493),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__10486),
            .DIN(N__10485),
            .DOUT(N__10484),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__10486),
            .PADOUT(N__10485),
            .PADIN(N__10484),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__10477),
            .DIN(N__10476),
            .DOUT(N__10475),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__10477),
            .PADOUT(N__10476),
            .PADIN(N__10475),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__10468),
            .DIN(N__10467),
            .DOUT(N__10466),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__10468),
            .PADOUT(N__10467),
            .PADIN(N__10466),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7593),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__10459),
            .DIN(N__10458),
            .DOUT(N__10457),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__10459),
            .PADOUT(N__10458),
            .PADIN(N__10457),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8391),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__10450),
            .DIN(N__10449),
            .DOUT(N__10448),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__10450),
            .PADOUT(N__10449),
            .PADIN(N__10448),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5217),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__10441),
            .DIN(N__10440),
            .DOUT(N__10439),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__10441),
            .PADOUT(N__10440),
            .PADIN(N__10439),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__10432),
            .DIN(N__10431),
            .DOUT(N__10430),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__10432),
            .PADOUT(N__10431),
            .PADIN(N__10430),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2541 (
            .O(N__10413),
            .I(N__10408));
    InMux I__2540 (
            .O(N__10412),
            .I(N__10405));
    InMux I__2539 (
            .O(N__10411),
            .I(N__10401));
    LocalMux I__2538 (
            .O(N__10408),
            .I(N__10398));
    LocalMux I__2537 (
            .O(N__10405),
            .I(N__10395));
    InMux I__2536 (
            .O(N__10404),
            .I(N__10392));
    LocalMux I__2535 (
            .O(N__10401),
            .I(N__10389));
    Span4Mux_v I__2534 (
            .O(N__10398),
            .I(N__10382));
    Span4Mux_h I__2533 (
            .O(N__10395),
            .I(N__10382));
    LocalMux I__2532 (
            .O(N__10392),
            .I(N__10382));
    Sp12to4 I__2531 (
            .O(N__10389),
            .I(N__10379));
    Span4Mux_h I__2530 (
            .O(N__10382),
            .I(N__10376));
    Span12Mux_v I__2529 (
            .O(N__10379),
            .I(N__10373));
    Span4Mux_v I__2528 (
            .O(N__10376),
            .I(N__10370));
    Span12Mux_h I__2527 (
            .O(N__10373),
            .I(N__10367));
    Sp12to4 I__2526 (
            .O(N__10370),
            .I(N__10364));
    Odrv12 I__2525 (
            .O(N__10367),
            .I(DRA_c_6));
    Odrv12 I__2524 (
            .O(N__10364),
            .I(DRA_c_6));
    InMux I__2523 (
            .O(N__10359),
            .I(N__10354));
    InMux I__2522 (
            .O(N__10358),
            .I(N__10348));
    CascadeMux I__2521 (
            .O(N__10357),
            .I(N__10343));
    LocalMux I__2520 (
            .O(N__10354),
            .I(N__10335));
    InMux I__2519 (
            .O(N__10353),
            .I(N__10332));
    InMux I__2518 (
            .O(N__10352),
            .I(N__10329));
    InMux I__2517 (
            .O(N__10351),
            .I(N__10326));
    LocalMux I__2516 (
            .O(N__10348),
            .I(N__10323));
    InMux I__2515 (
            .O(N__10347),
            .I(N__10320));
    InMux I__2514 (
            .O(N__10346),
            .I(N__10317));
    InMux I__2513 (
            .O(N__10343),
            .I(N__10308));
    InMux I__2512 (
            .O(N__10342),
            .I(N__10308));
    InMux I__2511 (
            .O(N__10341),
            .I(N__10308));
    InMux I__2510 (
            .O(N__10340),
            .I(N__10308));
    InMux I__2509 (
            .O(N__10339),
            .I(N__10305));
    InMux I__2508 (
            .O(N__10338),
            .I(N__10300));
    Span4Mux_h I__2507 (
            .O(N__10335),
            .I(N__10285));
    LocalMux I__2506 (
            .O(N__10332),
            .I(N__10285));
    LocalMux I__2505 (
            .O(N__10329),
            .I(N__10285));
    LocalMux I__2504 (
            .O(N__10326),
            .I(N__10285));
    Span4Mux_v I__2503 (
            .O(N__10323),
            .I(N__10282));
    LocalMux I__2502 (
            .O(N__10320),
            .I(N__10273));
    LocalMux I__2501 (
            .O(N__10317),
            .I(N__10273));
    LocalMux I__2500 (
            .O(N__10308),
            .I(N__10273));
    LocalMux I__2499 (
            .O(N__10305),
            .I(N__10273));
    InMux I__2498 (
            .O(N__10304),
            .I(N__10268));
    InMux I__2497 (
            .O(N__10303),
            .I(N__10268));
    LocalMux I__2496 (
            .O(N__10300),
            .I(N__10265));
    InMux I__2495 (
            .O(N__10299),
            .I(N__10260));
    InMux I__2494 (
            .O(N__10298),
            .I(N__10260));
    InMux I__2493 (
            .O(N__10297),
            .I(N__10257));
    InMux I__2492 (
            .O(N__10296),
            .I(N__10252));
    InMux I__2491 (
            .O(N__10295),
            .I(N__10252));
    InMux I__2490 (
            .O(N__10294),
            .I(N__10249));
    Span4Mux_v I__2489 (
            .O(N__10285),
            .I(N__10246));
    Span4Mux_h I__2488 (
            .O(N__10282),
            .I(N__10239));
    Span4Mux_v I__2487 (
            .O(N__10273),
            .I(N__10239));
    LocalMux I__2486 (
            .O(N__10268),
            .I(N__10239));
    Sp12to4 I__2485 (
            .O(N__10265),
            .I(N__10232));
    LocalMux I__2484 (
            .O(N__10260),
            .I(N__10232));
    LocalMux I__2483 (
            .O(N__10257),
            .I(N__10232));
    LocalMux I__2482 (
            .O(N__10252),
            .I(N__10227));
    LocalMux I__2481 (
            .O(N__10249),
            .I(N__10227));
    Sp12to4 I__2480 (
            .O(N__10246),
            .I(N__10222));
    Sp12to4 I__2479 (
            .O(N__10239),
            .I(N__10222));
    Span12Mux_h I__2478 (
            .O(N__10232),
            .I(N__10219));
    Span12Mux_v I__2477 (
            .O(N__10227),
            .I(N__10216));
    Span12Mux_h I__2476 (
            .O(N__10222),
            .I(N__10213));
    Span12Mux_v I__2475 (
            .O(N__10219),
            .I(N__10208));
    Span12Mux_h I__2474 (
            .O(N__10216),
            .I(N__10208));
    Span12Mux_v I__2473 (
            .O(N__10213),
            .I(N__10205));
    Odrv12 I__2472 (
            .O(N__10208),
            .I(AGNUS_REV_c));
    Odrv12 I__2471 (
            .O(N__10205),
            .I(AGNUS_REV_c));
    InMux I__2470 (
            .O(N__10200),
            .I(N__10195));
    InMux I__2469 (
            .O(N__10199),
            .I(N__10192));
    InMux I__2468 (
            .O(N__10198),
            .I(N__10189));
    LocalMux I__2467 (
            .O(N__10195),
            .I(N__10183));
    LocalMux I__2466 (
            .O(N__10192),
            .I(N__10183));
    LocalMux I__2465 (
            .O(N__10189),
            .I(N__10180));
    InMux I__2464 (
            .O(N__10188),
            .I(N__10177));
    Span4Mux_v I__2463 (
            .O(N__10183),
            .I(N__10174));
    Span4Mux_v I__2462 (
            .O(N__10180),
            .I(N__10169));
    LocalMux I__2461 (
            .O(N__10177),
            .I(N__10169));
    Span4Mux_v I__2460 (
            .O(N__10174),
            .I(N__10166));
    Span4Mux_v I__2459 (
            .O(N__10169),
            .I(N__10163));
    Sp12to4 I__2458 (
            .O(N__10166),
            .I(N__10158));
    Sp12to4 I__2457 (
            .O(N__10163),
            .I(N__10158));
    Span12Mux_h I__2456 (
            .O(N__10158),
            .I(N__10155));
    Odrv12 I__2455 (
            .O(N__10155),
            .I(DRA_c_5));
    InMux I__2454 (
            .O(N__10152),
            .I(N__10146));
    InMux I__2453 (
            .O(N__10151),
            .I(N__10146));
    LocalMux I__2452 (
            .O(N__10146),
            .I(N__10143));
    Odrv12 I__2451 (
            .O(N__10143),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__2450 (
            .O(N__10140),
            .I(N__10137));
    LocalMux I__2449 (
            .O(N__10137),
            .I(N__10125));
    ClkMux I__2448 (
            .O(N__10136),
            .I(N__10104));
    ClkMux I__2447 (
            .O(N__10135),
            .I(N__10104));
    ClkMux I__2446 (
            .O(N__10134),
            .I(N__10104));
    ClkMux I__2445 (
            .O(N__10133),
            .I(N__10104));
    ClkMux I__2444 (
            .O(N__10132),
            .I(N__10104));
    ClkMux I__2443 (
            .O(N__10131),
            .I(N__10104));
    ClkMux I__2442 (
            .O(N__10130),
            .I(N__10104));
    ClkMux I__2441 (
            .O(N__10129),
            .I(N__10104));
    ClkMux I__2440 (
            .O(N__10128),
            .I(N__10104));
    Glb2LocalMux I__2439 (
            .O(N__10125),
            .I(N__10104));
    GlobalMux I__2438 (
            .O(N__10104),
            .I(N__10101));
    gio2CtrlBuf I__2437 (
            .O(N__10101),
            .I(C3_c_g));
    CEMux I__2436 (
            .O(N__10098),
            .I(N__10094));
    CEMux I__2435 (
            .O(N__10097),
            .I(N__10087));
    LocalMux I__2434 (
            .O(N__10094),
            .I(N__10083));
    CEMux I__2433 (
            .O(N__10093),
            .I(N__10080));
    CEMux I__2432 (
            .O(N__10092),
            .I(N__10077));
    CEMux I__2431 (
            .O(N__10091),
            .I(N__10074));
    CEMux I__2430 (
            .O(N__10090),
            .I(N__10071));
    LocalMux I__2429 (
            .O(N__10087),
            .I(N__10068));
    CEMux I__2428 (
            .O(N__10086),
            .I(N__10065));
    Span4Mux_v I__2427 (
            .O(N__10083),
            .I(N__10059));
    LocalMux I__2426 (
            .O(N__10080),
            .I(N__10059));
    LocalMux I__2425 (
            .O(N__10077),
            .I(N__10056));
    LocalMux I__2424 (
            .O(N__10074),
            .I(N__10053));
    LocalMux I__2423 (
            .O(N__10071),
            .I(N__10046));
    Span4Mux_v I__2422 (
            .O(N__10068),
            .I(N__10046));
    LocalMux I__2421 (
            .O(N__10065),
            .I(N__10046));
    CEMux I__2420 (
            .O(N__10064),
            .I(N__10043));
    Span4Mux_h I__2419 (
            .O(N__10059),
            .I(N__10038));
    Span4Mux_h I__2418 (
            .O(N__10056),
            .I(N__10038));
    Span4Mux_h I__2417 (
            .O(N__10053),
            .I(N__10035));
    Span4Mux_h I__2416 (
            .O(N__10046),
            .I(N__10032));
    LocalMux I__2415 (
            .O(N__10043),
            .I(N__10029));
    Odrv4 I__2414 (
            .O(N__10038),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ));
    Odrv4 I__2413 (
            .O(N__10035),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ));
    Odrv4 I__2412 (
            .O(N__10032),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ));
    Odrv12 I__2411 (
            .O(N__10029),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ));
    InMux I__2410 (
            .O(N__10020),
            .I(N__10012));
    InMux I__2409 (
            .O(N__10019),
            .I(N__10009));
    InMux I__2408 (
            .O(N__10018),
            .I(N__10006));
    InMux I__2407 (
            .O(N__10017),
            .I(N__10003));
    InMux I__2406 (
            .O(N__10016),
            .I(N__9998));
    InMux I__2405 (
            .O(N__10015),
            .I(N__9998));
    LocalMux I__2404 (
            .O(N__10012),
            .I(N__9991));
    LocalMux I__2403 (
            .O(N__10009),
            .I(N__9983));
    LocalMux I__2402 (
            .O(N__10006),
            .I(N__9975));
    LocalMux I__2401 (
            .O(N__10003),
            .I(N__9965));
    LocalMux I__2400 (
            .O(N__9998),
            .I(N__9943));
    SRMux I__2399 (
            .O(N__9997),
            .I(N__9852));
    SRMux I__2398 (
            .O(N__9996),
            .I(N__9852));
    SRMux I__2397 (
            .O(N__9995),
            .I(N__9852));
    SRMux I__2396 (
            .O(N__9994),
            .I(N__9852));
    Glb2LocalMux I__2395 (
            .O(N__9991),
            .I(N__9852));
    SRMux I__2394 (
            .O(N__9990),
            .I(N__9852));
    SRMux I__2393 (
            .O(N__9989),
            .I(N__9852));
    SRMux I__2392 (
            .O(N__9988),
            .I(N__9852));
    SRMux I__2391 (
            .O(N__9987),
            .I(N__9852));
    SRMux I__2390 (
            .O(N__9986),
            .I(N__9852));
    Glb2LocalMux I__2389 (
            .O(N__9983),
            .I(N__9852));
    SRMux I__2388 (
            .O(N__9982),
            .I(N__9852));
    SRMux I__2387 (
            .O(N__9981),
            .I(N__9852));
    SRMux I__2386 (
            .O(N__9980),
            .I(N__9852));
    SRMux I__2385 (
            .O(N__9979),
            .I(N__9852));
    SRMux I__2384 (
            .O(N__9978),
            .I(N__9852));
    Glb2LocalMux I__2383 (
            .O(N__9975),
            .I(N__9852));
    SRMux I__2382 (
            .O(N__9974),
            .I(N__9852));
    SRMux I__2381 (
            .O(N__9973),
            .I(N__9852));
    SRMux I__2380 (
            .O(N__9972),
            .I(N__9852));
    SRMux I__2379 (
            .O(N__9971),
            .I(N__9852));
    SRMux I__2378 (
            .O(N__9970),
            .I(N__9852));
    SRMux I__2377 (
            .O(N__9969),
            .I(N__9852));
    SRMux I__2376 (
            .O(N__9968),
            .I(N__9852));
    Glb2LocalMux I__2375 (
            .O(N__9965),
            .I(N__9852));
    SRMux I__2374 (
            .O(N__9964),
            .I(N__9852));
    SRMux I__2373 (
            .O(N__9963),
            .I(N__9852));
    SRMux I__2372 (
            .O(N__9962),
            .I(N__9852));
    SRMux I__2371 (
            .O(N__9961),
            .I(N__9852));
    SRMux I__2370 (
            .O(N__9960),
            .I(N__9852));
    SRMux I__2369 (
            .O(N__9959),
            .I(N__9852));
    SRMux I__2368 (
            .O(N__9958),
            .I(N__9852));
    SRMux I__2367 (
            .O(N__9957),
            .I(N__9852));
    SRMux I__2366 (
            .O(N__9956),
            .I(N__9852));
    SRMux I__2365 (
            .O(N__9955),
            .I(N__9852));
    SRMux I__2364 (
            .O(N__9954),
            .I(N__9852));
    SRMux I__2363 (
            .O(N__9953),
            .I(N__9852));
    SRMux I__2362 (
            .O(N__9952),
            .I(N__9852));
    SRMux I__2361 (
            .O(N__9951),
            .I(N__9852));
    SRMux I__2360 (
            .O(N__9950),
            .I(N__9852));
    SRMux I__2359 (
            .O(N__9949),
            .I(N__9852));
    SRMux I__2358 (
            .O(N__9948),
            .I(N__9852));
    SRMux I__2357 (
            .O(N__9947),
            .I(N__9852));
    SRMux I__2356 (
            .O(N__9946),
            .I(N__9852));
    Glb2LocalMux I__2355 (
            .O(N__9943),
            .I(N__9852));
    GlobalMux I__2354 (
            .O(N__9852),
            .I(N__9849));
    gio2CtrlBuf I__2353 (
            .O(N__9849),
            .I(RESETn_c_i_g));
    CascadeMux I__2352 (
            .O(N__9846),
            .I(N__9843));
    InMux I__2351 (
            .O(N__9843),
            .I(N__9840));
    LocalMux I__2350 (
            .O(N__9840),
            .I(N__9837));
    Span4Mux_h I__2349 (
            .O(N__9837),
            .I(N__9834));
    Odrv4 I__2348 (
            .O(N__9834),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2347 (
            .O(N__9831),
            .I(N__9823));
    InMux I__2346 (
            .O(N__9830),
            .I(N__9823));
    InMux I__2345 (
            .O(N__9829),
            .I(N__9820));
    InMux I__2344 (
            .O(N__9828),
            .I(N__9817));
    LocalMux I__2343 (
            .O(N__9823),
            .I(N__9814));
    LocalMux I__2342 (
            .O(N__9820),
            .I(N__9809));
    LocalMux I__2341 (
            .O(N__9817),
            .I(N__9809));
    Span4Mux_v I__2340 (
            .O(N__9814),
            .I(N__9806));
    Span4Mux_v I__2339 (
            .O(N__9809),
            .I(N__9803));
    Span4Mux_h I__2338 (
            .O(N__9806),
            .I(N__9800));
    Sp12to4 I__2337 (
            .O(N__9803),
            .I(N__9797));
    Sp12to4 I__2336 (
            .O(N__9800),
            .I(N__9792));
    Span12Mux_h I__2335 (
            .O(N__9797),
            .I(N__9792));
    Odrv12 I__2334 (
            .O(N__9792),
            .I(DRA_c_7));
    InMux I__2333 (
            .O(N__9789),
            .I(N__9786));
    LocalMux I__2332 (
            .O(N__9786),
            .I(N__9783));
    Span4Mux_h I__2331 (
            .O(N__9783),
            .I(N__9780));
    Odrv4 I__2330 (
            .O(N__9780),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2329 (
            .O(N__9777),
            .I(N__9774));
    LocalMux I__2328 (
            .O(N__9774),
            .I(N__9771));
    Odrv4 I__2327 (
            .O(N__9771),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2326 (
            .O(N__9768),
            .I(N__9765));
    LocalMux I__2325 (
            .O(N__9765),
            .I(N__9759));
    InMux I__2324 (
            .O(N__9764),
            .I(N__9756));
    InMux I__2323 (
            .O(N__9763),
            .I(N__9751));
    InMux I__2322 (
            .O(N__9762),
            .I(N__9751));
    Span4Mux_h I__2321 (
            .O(N__9759),
            .I(N__9746));
    LocalMux I__2320 (
            .O(N__9756),
            .I(N__9746));
    LocalMux I__2319 (
            .O(N__9751),
            .I(N__9741));
    Sp12to4 I__2318 (
            .O(N__9746),
            .I(N__9741));
    Span12Mux_v I__2317 (
            .O(N__9741),
            .I(N__9738));
    Span12Mux_h I__2316 (
            .O(N__9738),
            .I(N__9735));
    Odrv12 I__2315 (
            .O(N__9735),
            .I(DRA_c_3));
    InMux I__2314 (
            .O(N__9732),
            .I(N__9729));
    LocalMux I__2313 (
            .O(N__9729),
            .I(N__9726));
    Odrv4 I__2312 (
            .O(N__9726),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__2311 (
            .O(N__9723),
            .I(N__9717));
    InMux I__2310 (
            .O(N__9722),
            .I(N__9714));
    InMux I__2309 (
            .O(N__9721),
            .I(N__9709));
    InMux I__2308 (
            .O(N__9720),
            .I(N__9709));
    LocalMux I__2307 (
            .O(N__9717),
            .I(N__9704));
    LocalMux I__2306 (
            .O(N__9714),
            .I(N__9704));
    LocalMux I__2305 (
            .O(N__9709),
            .I(N__9701));
    Span4Mux_v I__2304 (
            .O(N__9704),
            .I(N__9698));
    Span4Mux_h I__2303 (
            .O(N__9701),
            .I(N__9695));
    Span4Mux_v I__2302 (
            .O(N__9698),
            .I(N__9692));
    Span4Mux_v I__2301 (
            .O(N__9695),
            .I(N__9689));
    Sp12to4 I__2300 (
            .O(N__9692),
            .I(N__9684));
    Sp12to4 I__2299 (
            .O(N__9689),
            .I(N__9684));
    Span12Mux_h I__2298 (
            .O(N__9684),
            .I(N__9681));
    Odrv12 I__2297 (
            .O(N__9681),
            .I(DRA_c_4));
    InMux I__2296 (
            .O(N__9678),
            .I(N__9675));
    LocalMux I__2295 (
            .O(N__9675),
            .I(N__9672));
    Span4Mux_h I__2294 (
            .O(N__9672),
            .I(N__9669));
    Odrv4 I__2293 (
            .O(N__9669),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    CascadeMux I__2292 (
            .O(N__9666),
            .I(N__9663));
    InMux I__2291 (
            .O(N__9663),
            .I(N__9659));
    InMux I__2290 (
            .O(N__9662),
            .I(N__9656));
    LocalMux I__2289 (
            .O(N__9659),
            .I(N__9651));
    LocalMux I__2288 (
            .O(N__9656),
            .I(N__9651));
    Span12Mux_h I__2287 (
            .O(N__9651),
            .I(N__9648));
    Span12Mux_v I__2286 (
            .O(N__9648),
            .I(N__9645));
    Odrv12 I__2285 (
            .O(N__9645),
            .I(DRA_c_0));
    InMux I__2284 (
            .O(N__9642),
            .I(N__9639));
    LocalMux I__2283 (
            .O(N__9639),
            .I(N__9636));
    Span4Mux_h I__2282 (
            .O(N__9636),
            .I(N__9633));
    Odrv4 I__2281 (
            .O(N__9633),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__2280 (
            .O(N__9630),
            .I(N__9625));
    InMux I__2279 (
            .O(N__9629),
            .I(N__9622));
    CascadeMux I__2278 (
            .O(N__9628),
            .I(N__9619));
    LocalMux I__2277 (
            .O(N__9625),
            .I(N__9615));
    LocalMux I__2276 (
            .O(N__9622),
            .I(N__9612));
    InMux I__2275 (
            .O(N__9619),
            .I(N__9609));
    InMux I__2274 (
            .O(N__9618),
            .I(N__9606));
    Span4Mux_v I__2273 (
            .O(N__9615),
            .I(N__9603));
    Span4Mux_v I__2272 (
            .O(N__9612),
            .I(N__9596));
    LocalMux I__2271 (
            .O(N__9609),
            .I(N__9596));
    LocalMux I__2270 (
            .O(N__9606),
            .I(N__9596));
    Span4Mux_v I__2269 (
            .O(N__9603),
            .I(N__9593));
    Span4Mux_v I__2268 (
            .O(N__9596),
            .I(N__9590));
    Sp12to4 I__2267 (
            .O(N__9593),
            .I(N__9585));
    Sp12to4 I__2266 (
            .O(N__9590),
            .I(N__9585));
    Span12Mux_h I__2265 (
            .O(N__9585),
            .I(N__9582));
    Span12Mux_v I__2264 (
            .O(N__9582),
            .I(N__9579));
    Odrv12 I__2263 (
            .O(N__9579),
            .I(DRA_c_9));
    InMux I__2262 (
            .O(N__9576),
            .I(N__9571));
    InMux I__2261 (
            .O(N__9575),
            .I(N__9568));
    InMux I__2260 (
            .O(N__9574),
            .I(N__9565));
    LocalMux I__2259 (
            .O(N__9571),
            .I(N__9562));
    LocalMux I__2258 (
            .O(N__9568),
            .I(N__9557));
    LocalMux I__2257 (
            .O(N__9565),
            .I(N__9557));
    Span4Mux_v I__2256 (
            .O(N__9562),
            .I(N__9553));
    Span4Mux_v I__2255 (
            .O(N__9557),
            .I(N__9550));
    InMux I__2254 (
            .O(N__9556),
            .I(N__9547));
    Span4Mux_h I__2253 (
            .O(N__9553),
            .I(N__9544));
    Span4Mux_h I__2252 (
            .O(N__9550),
            .I(N__9541));
    LocalMux I__2251 (
            .O(N__9547),
            .I(N__9538));
    Sp12to4 I__2250 (
            .O(N__9544),
            .I(N__9531));
    Sp12to4 I__2249 (
            .O(N__9541),
            .I(N__9531));
    Span12Mux_h I__2248 (
            .O(N__9538),
            .I(N__9531));
    Odrv12 I__2247 (
            .O(N__9531),
            .I(DRA_c_8));
    InMux I__2246 (
            .O(N__9528),
            .I(N__9525));
    LocalMux I__2245 (
            .O(N__9525),
            .I(N__9522));
    Span12Mux_v I__2244 (
            .O(N__9522),
            .I(N__9519));
    Odrv12 I__2243 (
            .O(N__9519),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2242 (
            .O(N__9516),
            .I(N__9509));
    InMux I__2241 (
            .O(N__9515),
            .I(N__9509));
    InMux I__2240 (
            .O(N__9514),
            .I(N__9505));
    LocalMux I__2239 (
            .O(N__9509),
            .I(N__9502));
    InMux I__2238 (
            .O(N__9508),
            .I(N__9499));
    LocalMux I__2237 (
            .O(N__9505),
            .I(N__9492));
    Span4Mux_h I__2236 (
            .O(N__9502),
            .I(N__9492));
    LocalMux I__2235 (
            .O(N__9499),
            .I(N__9492));
    Span4Mux_v I__2234 (
            .O(N__9492),
            .I(N__9489));
    Sp12to4 I__2233 (
            .O(N__9489),
            .I(N__9486));
    Span12Mux_h I__2232 (
            .O(N__9486),
            .I(N__9483));
    Span12Mux_v I__2231 (
            .O(N__9483),
            .I(N__9480));
    Odrv12 I__2230 (
            .O(N__9480),
            .I(DRA_c_2));
    InMux I__2229 (
            .O(N__9477),
            .I(N__9474));
    LocalMux I__2228 (
            .O(N__9474),
            .I(N__9469));
    InMux I__2227 (
            .O(N__9473),
            .I(N__9466));
    InMux I__2226 (
            .O(N__9472),
            .I(N__9462));
    Span4Mux_v I__2225 (
            .O(N__9469),
            .I(N__9459));
    LocalMux I__2224 (
            .O(N__9466),
            .I(N__9456));
    InMux I__2223 (
            .O(N__9465),
            .I(N__9453));
    LocalMux I__2222 (
            .O(N__9462),
            .I(N__9450));
    Sp12to4 I__2221 (
            .O(N__9459),
            .I(N__9447));
    Sp12to4 I__2220 (
            .O(N__9456),
            .I(N__9442));
    LocalMux I__2219 (
            .O(N__9453),
            .I(N__9442));
    Span12Mux_h I__2218 (
            .O(N__9450),
            .I(N__9439));
    Span12Mux_h I__2217 (
            .O(N__9447),
            .I(N__9436));
    Span12Mux_v I__2216 (
            .O(N__9442),
            .I(N__9433));
    Span12Mux_v I__2215 (
            .O(N__9439),
            .I(N__9430));
    Span12Mux_v I__2214 (
            .O(N__9436),
            .I(N__9425));
    Span12Mux_h I__2213 (
            .O(N__9433),
            .I(N__9425));
    Odrv12 I__2212 (
            .O(N__9430),
            .I(DRA_c_1));
    Odrv12 I__2211 (
            .O(N__9425),
            .I(DRA_c_1));
    InMux I__2210 (
            .O(N__9420),
            .I(N__9414));
    InMux I__2209 (
            .O(N__9419),
            .I(N__9414));
    LocalMux I__2208 (
            .O(N__9414),
            .I(N__9411));
    Odrv12 I__2207 (
            .O(N__9411),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__2206 (
            .O(N__9408),
            .I(N__9405));
    LocalMux I__2205 (
            .O(N__9405),
            .I(N__9402));
    Span4Mux_h I__2204 (
            .O(N__9402),
            .I(N__9399));
    Odrv4 I__2203 (
            .O(N__9399),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2202 (
            .O(N__9396),
            .I(N__9393));
    LocalMux I__2201 (
            .O(N__9393),
            .I(N__9390));
    Odrv4 I__2200 (
            .O(N__9390),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2199 (
            .O(N__9387),
            .I(N__9384));
    LocalMux I__2198 (
            .O(N__9384),
            .I(N__9381));
    Span4Mux_h I__2197 (
            .O(N__9381),
            .I(N__9378));
    Odrv4 I__2196 (
            .O(N__9378),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2195 (
            .O(N__9375),
            .I(N__9372));
    LocalMux I__2194 (
            .O(N__9372),
            .I(N__9369));
    Odrv4 I__2193 (
            .O(N__9369),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__2192 (
            .O(N__9366),
            .I(N__9363));
    LocalMux I__2191 (
            .O(N__9363),
            .I(N__9360));
    Odrv4 I__2190 (
            .O(N__9360),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__2189 (
            .O(N__9357),
            .I(N__9354));
    LocalMux I__2188 (
            .O(N__9354),
            .I(N__9351));
    Span4Mux_h I__2187 (
            .O(N__9351),
            .I(N__9348));
    Odrv4 I__2186 (
            .O(N__9348),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__2185 (
            .O(N__9345),
            .I(N__9342));
    LocalMux I__2184 (
            .O(N__9342),
            .I(N__9339));
    Span4Mux_h I__2183 (
            .O(N__9339),
            .I(N__9336));
    Span4Mux_h I__2182 (
            .O(N__9336),
            .I(N__9333));
    Odrv4 I__2181 (
            .O(N__9333),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__2180 (
            .O(N__9330),
            .I(N__9327));
    LocalMux I__2179 (
            .O(N__9327),
            .I(N__9324));
    Span4Mux_h I__2178 (
            .O(N__9324),
            .I(N__9321));
    Odrv4 I__2177 (
            .O(N__9321),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2176 (
            .O(N__9318),
            .I(N__9315));
    LocalMux I__2175 (
            .O(N__9315),
            .I(N__9312));
    Span4Mux_h I__2174 (
            .O(N__9312),
            .I(N__9309));
    Odrv4 I__2173 (
            .O(N__9309),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    CEMux I__2172 (
            .O(N__9306),
            .I(N__9302));
    CEMux I__2171 (
            .O(N__9305),
            .I(N__9299));
    LocalMux I__2170 (
            .O(N__9302),
            .I(N__9296));
    LocalMux I__2169 (
            .O(N__9299),
            .I(N__9293));
    Span4Mux_v I__2168 (
            .O(N__9296),
            .I(N__9287));
    Span12Mux_h I__2167 (
            .O(N__9293),
            .I(N__9284));
    CEMux I__2166 (
            .O(N__9292),
            .I(N__9281));
    CEMux I__2165 (
            .O(N__9291),
            .I(N__9278));
    CEMux I__2164 (
            .O(N__9290),
            .I(N__9275));
    Odrv4 I__2163 (
            .O(N__9287),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ));
    Odrv12 I__2162 (
            .O(N__9284),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ));
    LocalMux I__2161 (
            .O(N__9281),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ));
    LocalMux I__2160 (
            .O(N__9278),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ));
    LocalMux I__2159 (
            .O(N__9275),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ));
    InMux I__2158 (
            .O(N__9264),
            .I(N__9261));
    LocalMux I__2157 (
            .O(N__9261),
            .I(N__9257));
    InMux I__2156 (
            .O(N__9260),
            .I(N__9254));
    Span4Mux_v I__2155 (
            .O(N__9257),
            .I(N__9251));
    LocalMux I__2154 (
            .O(N__9254),
            .I(N__9248));
    Span4Mux_h I__2153 (
            .O(N__9251),
            .I(N__9243));
    Span4Mux_v I__2152 (
            .O(N__9248),
            .I(N__9243));
    Sp12to4 I__2151 (
            .O(N__9243),
            .I(N__9240));
    Span12Mux_h I__2150 (
            .O(N__9240),
            .I(N__9237));
    Odrv12 I__2149 (
            .O(N__9237),
            .I(RAS0n_c));
    InMux I__2148 (
            .O(N__9234),
            .I(N__9231));
    LocalMux I__2147 (
            .O(N__9231),
            .I(N__9228));
    Span4Mux_h I__2146 (
            .O(N__9228),
            .I(N__9225));
    Odrv4 I__2145 (
            .O(N__9225),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    InMux I__2144 (
            .O(N__9222),
            .I(N__9214));
    InMux I__2143 (
            .O(N__9221),
            .I(N__9211));
    InMux I__2142 (
            .O(N__9220),
            .I(N__9206));
    InMux I__2141 (
            .O(N__9219),
            .I(N__9206));
    InMux I__2140 (
            .O(N__9218),
            .I(N__9201));
    InMux I__2139 (
            .O(N__9217),
            .I(N__9201));
    LocalMux I__2138 (
            .O(N__9214),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    LocalMux I__2137 (
            .O(N__9211),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    LocalMux I__2136 (
            .O(N__9206),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    LocalMux I__2135 (
            .O(N__9201),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    CascadeMux I__2134 (
            .O(N__9192),
            .I(N__9185));
    CascadeMux I__2133 (
            .O(N__9191),
            .I(N__9182));
    CascadeMux I__2132 (
            .O(N__9190),
            .I(N__9179));
    CascadeMux I__2131 (
            .O(N__9189),
            .I(N__9174));
    CascadeMux I__2130 (
            .O(N__9188),
            .I(N__9171));
    InMux I__2129 (
            .O(N__9185),
            .I(N__9166));
    InMux I__2128 (
            .O(N__9182),
            .I(N__9166));
    InMux I__2127 (
            .O(N__9179),
            .I(N__9163));
    CascadeMux I__2126 (
            .O(N__9178),
            .I(N__9159));
    InMux I__2125 (
            .O(N__9177),
            .I(N__9156));
    InMux I__2124 (
            .O(N__9174),
            .I(N__9153));
    InMux I__2123 (
            .O(N__9171),
            .I(N__9150));
    LocalMux I__2122 (
            .O(N__9166),
            .I(N__9147));
    LocalMux I__2121 (
            .O(N__9163),
            .I(N__9144));
    InMux I__2120 (
            .O(N__9162),
            .I(N__9139));
    InMux I__2119 (
            .O(N__9159),
            .I(N__9139));
    LocalMux I__2118 (
            .O(N__9156),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__2117 (
            .O(N__9153),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__2116 (
            .O(N__9150),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__2115 (
            .O(N__9147),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__2114 (
            .O(N__9144),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__2113 (
            .O(N__9139),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    InMux I__2112 (
            .O(N__9126),
            .I(N__9123));
    LocalMux I__2111 (
            .O(N__9123),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__2110 (
            .O(N__9120),
            .I(N__9117));
    LocalMux I__2109 (
            .O(N__9117),
            .I(N__9114));
    Span12Mux_s7_h I__2108 (
            .O(N__9114),
            .I(N__9111));
    Span12Mux_v I__2107 (
            .O(N__9111),
            .I(N__9108));
    Odrv12 I__2106 (
            .O(N__9108),
            .I(CMA_c_3));
    InMux I__2105 (
            .O(N__9105),
            .I(N__9102));
    LocalMux I__2104 (
            .O(N__9102),
            .I(N__9072));
    ClkMux I__2103 (
            .O(N__9101),
            .I(N__8997));
    ClkMux I__2102 (
            .O(N__9100),
            .I(N__8997));
    ClkMux I__2101 (
            .O(N__9099),
            .I(N__8997));
    ClkMux I__2100 (
            .O(N__9098),
            .I(N__8997));
    ClkMux I__2099 (
            .O(N__9097),
            .I(N__8997));
    ClkMux I__2098 (
            .O(N__9096),
            .I(N__8997));
    ClkMux I__2097 (
            .O(N__9095),
            .I(N__8997));
    ClkMux I__2096 (
            .O(N__9094),
            .I(N__8997));
    ClkMux I__2095 (
            .O(N__9093),
            .I(N__8997));
    ClkMux I__2094 (
            .O(N__9092),
            .I(N__8997));
    ClkMux I__2093 (
            .O(N__9091),
            .I(N__8997));
    ClkMux I__2092 (
            .O(N__9090),
            .I(N__8997));
    ClkMux I__2091 (
            .O(N__9089),
            .I(N__8997));
    ClkMux I__2090 (
            .O(N__9088),
            .I(N__8997));
    ClkMux I__2089 (
            .O(N__9087),
            .I(N__8997));
    ClkMux I__2088 (
            .O(N__9086),
            .I(N__8997));
    ClkMux I__2087 (
            .O(N__9085),
            .I(N__8997));
    ClkMux I__2086 (
            .O(N__9084),
            .I(N__8997));
    ClkMux I__2085 (
            .O(N__9083),
            .I(N__8997));
    ClkMux I__2084 (
            .O(N__9082),
            .I(N__8997));
    ClkMux I__2083 (
            .O(N__9081),
            .I(N__8997));
    ClkMux I__2082 (
            .O(N__9080),
            .I(N__8997));
    ClkMux I__2081 (
            .O(N__9079),
            .I(N__8997));
    ClkMux I__2080 (
            .O(N__9078),
            .I(N__8997));
    ClkMux I__2079 (
            .O(N__9077),
            .I(N__8997));
    ClkMux I__2078 (
            .O(N__9076),
            .I(N__8997));
    ClkMux I__2077 (
            .O(N__9075),
            .I(N__8997));
    Glb2LocalMux I__2076 (
            .O(N__9072),
            .I(N__8997));
    ClkMux I__2075 (
            .O(N__9071),
            .I(N__8997));
    ClkMux I__2074 (
            .O(N__9070),
            .I(N__8997));
    ClkMux I__2073 (
            .O(N__9069),
            .I(N__8997));
    ClkMux I__2072 (
            .O(N__9068),
            .I(N__8997));
    ClkMux I__2071 (
            .O(N__9067),
            .I(N__8997));
    ClkMux I__2070 (
            .O(N__9066),
            .I(N__8997));
    GlobalMux I__2069 (
            .O(N__8997),
            .I(CLK80_PLL));
    CEMux I__2068 (
            .O(N__8994),
            .I(N__8990));
    CEMux I__2067 (
            .O(N__8993),
            .I(N__8985));
    LocalMux I__2066 (
            .O(N__8990),
            .I(N__8980));
    CEMux I__2065 (
            .O(N__8989),
            .I(N__8977));
    CEMux I__2064 (
            .O(N__8988),
            .I(N__8974));
    LocalMux I__2063 (
            .O(N__8985),
            .I(N__8971));
    CEMux I__2062 (
            .O(N__8984),
            .I(N__8968));
    CEMux I__2061 (
            .O(N__8983),
            .I(N__8965));
    Odrv4 I__2060 (
            .O(N__8980),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__2059 (
            .O(N__8977),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__2058 (
            .O(N__8974),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__2057 (
            .O(N__8971),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__2056 (
            .O(N__8968),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__2055 (
            .O(N__8965),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    InMux I__2054 (
            .O(N__8952),
            .I(N__8948));
    InMux I__2053 (
            .O(N__8951),
            .I(N__8945));
    LocalMux I__2052 (
            .O(N__8948),
            .I(N__8942));
    LocalMux I__2051 (
            .O(N__8945),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    Odrv4 I__2050 (
            .O(N__8942),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    InMux I__2049 (
            .O(N__8937),
            .I(N__8934));
    LocalMux I__2048 (
            .O(N__8934),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10 ));
    CascadeMux I__2047 (
            .O(N__8931),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10_cascade_ ));
    CascadeMux I__2046 (
            .O(N__8928),
            .I(N__8925));
    InMux I__2045 (
            .O(N__8925),
            .I(N__8918));
    InMux I__2044 (
            .O(N__8924),
            .I(N__8918));
    InMux I__2043 (
            .O(N__8923),
            .I(N__8915));
    LocalMux I__2042 (
            .O(N__8918),
            .I(N__8912));
    LocalMux I__2041 (
            .O(N__8915),
            .I(N__8908));
    Span4Mux_v I__2040 (
            .O(N__8912),
            .I(N__8905));
    InMux I__2039 (
            .O(N__8911),
            .I(N__8902));
    Span4Mux_h I__2038 (
            .O(N__8908),
            .I(N__8899));
    Sp12to4 I__2037 (
            .O(N__8905),
            .I(N__8894));
    LocalMux I__2036 (
            .O(N__8902),
            .I(N__8894));
    Sp12to4 I__2035 (
            .O(N__8899),
            .I(N__8889));
    Span12Mux_h I__2034 (
            .O(N__8894),
            .I(N__8889));
    Span12Mux_v I__2033 (
            .O(N__8889),
            .I(N__8886));
    Odrv12 I__2032 (
            .O(N__8886),
            .I(DBRn_c));
    InMux I__2031 (
            .O(N__8883),
            .I(N__8877));
    InMux I__2030 (
            .O(N__8882),
            .I(N__8874));
    InMux I__2029 (
            .O(N__8881),
            .I(N__8869));
    InMux I__2028 (
            .O(N__8880),
            .I(N__8869));
    LocalMux I__2027 (
            .O(N__8877),
            .I(N__8859));
    LocalMux I__2026 (
            .O(N__8874),
            .I(N__8856));
    LocalMux I__2025 (
            .O(N__8869),
            .I(N__8853));
    ClkMux I__2024 (
            .O(N__8868),
            .I(N__8832));
    ClkMux I__2023 (
            .O(N__8867),
            .I(N__8832));
    ClkMux I__2022 (
            .O(N__8866),
            .I(N__8832));
    ClkMux I__2021 (
            .O(N__8865),
            .I(N__8832));
    ClkMux I__2020 (
            .O(N__8864),
            .I(N__8832));
    ClkMux I__2019 (
            .O(N__8863),
            .I(N__8832));
    ClkMux I__2018 (
            .O(N__8862),
            .I(N__8832));
    Glb2LocalMux I__2017 (
            .O(N__8859),
            .I(N__8832));
    Glb2LocalMux I__2016 (
            .O(N__8856),
            .I(N__8832));
    Glb2LocalMux I__2015 (
            .O(N__8853),
            .I(N__8832));
    GlobalMux I__2014 (
            .O(N__8832),
            .I(N__8829));
    gio2CtrlBuf I__2013 (
            .O(N__8829),
            .I(C1_c_g));
    CascadeMux I__2012 (
            .O(N__8826),
            .I(N__8822));
    InMux I__2011 (
            .O(N__8825),
            .I(N__8818));
    InMux I__2010 (
            .O(N__8822),
            .I(N__8814));
    InMux I__2009 (
            .O(N__8821),
            .I(N__8811));
    LocalMux I__2008 (
            .O(N__8818),
            .I(N__8808));
    InMux I__2007 (
            .O(N__8817),
            .I(N__8805));
    LocalMux I__2006 (
            .O(N__8814),
            .I(N__8802));
    LocalMux I__2005 (
            .O(N__8811),
            .I(N__8799));
    Span4Mux_v I__2004 (
            .O(N__8808),
            .I(N__8796));
    LocalMux I__2003 (
            .O(N__8805),
            .I(N__8793));
    Span4Mux_v I__2002 (
            .O(N__8802),
            .I(N__8790));
    Span4Mux_v I__2001 (
            .O(N__8799),
            .I(N__8785));
    Span4Mux_h I__2000 (
            .O(N__8796),
            .I(N__8785));
    Span4Mux_v I__1999 (
            .O(N__8793),
            .I(N__8780));
    Span4Mux_v I__1998 (
            .O(N__8790),
            .I(N__8780));
    Span4Mux_v I__1997 (
            .O(N__8785),
            .I(N__8777));
    Sp12to4 I__1996 (
            .O(N__8780),
            .I(N__8774));
    Sp12to4 I__1995 (
            .O(N__8777),
            .I(N__8769));
    Span12Mux_h I__1994 (
            .O(N__8774),
            .I(N__8769));
    Odrv12 I__1993 (
            .O(N__8769),
            .I(CLK40_PLL_i));
    IoInMux I__1992 (
            .O(N__8766),
            .I(N__8763));
    LocalMux I__1991 (
            .O(N__8763),
            .I(N__8758));
    IoInMux I__1990 (
            .O(N__8762),
            .I(N__8755));
    IoInMux I__1989 (
            .O(N__8761),
            .I(N__8752));
    Span4Mux_s3_v I__1988 (
            .O(N__8758),
            .I(N__8749));
    LocalMux I__1987 (
            .O(N__8755),
            .I(N__8746));
    LocalMux I__1986 (
            .O(N__8752),
            .I(N__8743));
    Span4Mux_h I__1985 (
            .O(N__8749),
            .I(N__8740));
    Span4Mux_s3_v I__1984 (
            .O(N__8746),
            .I(N__8737));
    Span4Mux_s3_h I__1983 (
            .O(N__8743),
            .I(N__8734));
    Sp12to4 I__1982 (
            .O(N__8740),
            .I(N__8729));
    Sp12to4 I__1981 (
            .O(N__8737),
            .I(N__8729));
    Span4Mux_h I__1980 (
            .O(N__8734),
            .I(N__8726));
    Span12Mux_h I__1979 (
            .O(N__8729),
            .I(N__8723));
    Span4Mux_h I__1978 (
            .O(N__8726),
            .I(N__8720));
    Span12Mux_v I__1977 (
            .O(N__8723),
            .I(N__8717));
    Span4Mux_h I__1976 (
            .O(N__8720),
            .I(N__8714));
    Odrv12 I__1975 (
            .O(N__8717),
            .I(CLK40_PLL_i_i));
    Odrv4 I__1974 (
            .O(N__8714),
            .I(CLK40_PLL_i_i));
    InMux I__1973 (
            .O(N__8709),
            .I(N__8696));
    InMux I__1972 (
            .O(N__8708),
            .I(N__8693));
    InMux I__1971 (
            .O(N__8707),
            .I(N__8688));
    InMux I__1970 (
            .O(N__8706),
            .I(N__8688));
    InMux I__1969 (
            .O(N__8705),
            .I(N__8685));
    InMux I__1968 (
            .O(N__8704),
            .I(N__8682));
    InMux I__1967 (
            .O(N__8703),
            .I(N__8677));
    InMux I__1966 (
            .O(N__8702),
            .I(N__8671));
    InMux I__1965 (
            .O(N__8701),
            .I(N__8666));
    InMux I__1964 (
            .O(N__8700),
            .I(N__8666));
    InMux I__1963 (
            .O(N__8699),
            .I(N__8663));
    LocalMux I__1962 (
            .O(N__8696),
            .I(N__8655));
    LocalMux I__1961 (
            .O(N__8693),
            .I(N__8655));
    LocalMux I__1960 (
            .O(N__8688),
            .I(N__8655));
    LocalMux I__1959 (
            .O(N__8685),
            .I(N__8652));
    LocalMux I__1958 (
            .O(N__8682),
            .I(N__8649));
    InMux I__1957 (
            .O(N__8681),
            .I(N__8644));
    InMux I__1956 (
            .O(N__8680),
            .I(N__8644));
    LocalMux I__1955 (
            .O(N__8677),
            .I(N__8641));
    InMux I__1954 (
            .O(N__8676),
            .I(N__8636));
    InMux I__1953 (
            .O(N__8675),
            .I(N__8636));
    InMux I__1952 (
            .O(N__8674),
            .I(N__8633));
    LocalMux I__1951 (
            .O(N__8671),
            .I(N__8628));
    LocalMux I__1950 (
            .O(N__8666),
            .I(N__8628));
    LocalMux I__1949 (
            .O(N__8663),
            .I(N__8625));
    InMux I__1948 (
            .O(N__8662),
            .I(N__8622));
    Span4Mux_v I__1947 (
            .O(N__8655),
            .I(N__8617));
    Span4Mux_v I__1946 (
            .O(N__8652),
            .I(N__8617));
    Span4Mux_v I__1945 (
            .O(N__8649),
            .I(N__8614));
    LocalMux I__1944 (
            .O(N__8644),
            .I(N__8611));
    Span4Mux_v I__1943 (
            .O(N__8641),
            .I(N__8606));
    LocalMux I__1942 (
            .O(N__8636),
            .I(N__8606));
    LocalMux I__1941 (
            .O(N__8633),
            .I(N__8603));
    Span4Mux_v I__1940 (
            .O(N__8628),
            .I(N__8600));
    Span4Mux_h I__1939 (
            .O(N__8625),
            .I(N__8595));
    LocalMux I__1938 (
            .O(N__8622),
            .I(N__8595));
    Span4Mux_h I__1937 (
            .O(N__8617),
            .I(N__8584));
    Span4Mux_v I__1936 (
            .O(N__8614),
            .I(N__8584));
    Span4Mux_v I__1935 (
            .O(N__8611),
            .I(N__8584));
    Span4Mux_v I__1934 (
            .O(N__8606),
            .I(N__8584));
    Span4Mux_v I__1933 (
            .O(N__8603),
            .I(N__8584));
    Span4Mux_h I__1932 (
            .O(N__8600),
            .I(N__8579));
    Span4Mux_v I__1931 (
            .O(N__8595),
            .I(N__8579));
    Sp12to4 I__1930 (
            .O(N__8584),
            .I(N__8574));
    Sp12to4 I__1929 (
            .O(N__8579),
            .I(N__8574));
    Span12Mux_h I__1928 (
            .O(N__8574),
            .I(N__8571));
    Odrv12 I__1927 (
            .O(N__8571),
            .I(RESETn_c));
    IoInMux I__1926 (
            .O(N__8568),
            .I(N__8565));
    LocalMux I__1925 (
            .O(N__8565),
            .I(N__8562));
    Span12Mux_s3_v I__1924 (
            .O(N__8562),
            .I(N__8559));
    Odrv12 I__1923 (
            .O(N__8559),
            .I(RESETn_c_i));
    InMux I__1922 (
            .O(N__8556),
            .I(N__8552));
    InMux I__1921 (
            .O(N__8555),
            .I(N__8549));
    LocalMux I__1920 (
            .O(N__8552),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__1919 (
            .O(N__8549),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__1918 (
            .O(N__8544),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__1917 (
            .O(N__8541),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    CascadeMux I__1916 (
            .O(N__8538),
            .I(N__8535));
    InMux I__1915 (
            .O(N__8535),
            .I(N__8532));
    LocalMux I__1914 (
            .O(N__8532),
            .I(N__8528));
    InMux I__1913 (
            .O(N__8531),
            .I(N__8525));
    Span4Mux_h I__1912 (
            .O(N__8528),
            .I(N__8522));
    LocalMux I__1911 (
            .O(N__8525),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv4 I__1910 (
            .O(N__8522),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    SRMux I__1909 (
            .O(N__8517),
            .I(N__8514));
    LocalMux I__1908 (
            .O(N__8514),
            .I(N__8511));
    Odrv4 I__1907 (
            .O(N__8511),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    IoInMux I__1906 (
            .O(N__8508),
            .I(N__8505));
    LocalMux I__1905 (
            .O(N__8505),
            .I(N__8502));
    Span4Mux_s2_v I__1904 (
            .O(N__8502),
            .I(N__8499));
    Sp12to4 I__1903 (
            .O(N__8499),
            .I(N__8496));
    Span12Mux_h I__1902 (
            .O(N__8496),
            .I(N__8493));
    Odrv12 I__1901 (
            .O(N__8493),
            .I(un1_LDSn_i_0_0));
    InMux I__1900 (
            .O(N__8490),
            .I(N__8486));
    InMux I__1899 (
            .O(N__8489),
            .I(N__8483));
    LocalMux I__1898 (
            .O(N__8486),
            .I(N__8478));
    LocalMux I__1897 (
            .O(N__8483),
            .I(N__8478));
    Span4Mux_v I__1896 (
            .O(N__8478),
            .I(N__8475));
    Span4Mux_h I__1895 (
            .O(N__8475),
            .I(N__8471));
    InMux I__1894 (
            .O(N__8474),
            .I(N__8468));
    Odrv4 I__1893 (
            .O(N__8471),
            .I(DS_ENm));
    LocalMux I__1892 (
            .O(N__8468),
            .I(DS_ENm));
    InMux I__1891 (
            .O(N__8463),
            .I(N__8459));
    InMux I__1890 (
            .O(N__8462),
            .I(N__8456));
    LocalMux I__1889 (
            .O(N__8459),
            .I(N__8448));
    LocalMux I__1888 (
            .O(N__8456),
            .I(N__8448));
    InMux I__1887 (
            .O(N__8455),
            .I(N__8441));
    InMux I__1886 (
            .O(N__8454),
            .I(N__8441));
    InMux I__1885 (
            .O(N__8453),
            .I(N__8441));
    Span4Mux_v I__1884 (
            .O(N__8448),
            .I(N__8438));
    LocalMux I__1883 (
            .O(N__8441),
            .I(N__8435));
    Span4Mux_h I__1882 (
            .O(N__8438),
            .I(N__8430));
    Span4Mux_v I__1881 (
            .O(N__8435),
            .I(N__8430));
    Sp12to4 I__1880 (
            .O(N__8430),
            .I(N__8427));
    Odrv12 I__1879 (
            .O(N__8427),
            .I(A_c_0));
    InMux I__1878 (
            .O(N__8424),
            .I(N__8420));
    InMux I__1877 (
            .O(N__8423),
            .I(N__8417));
    LocalMux I__1876 (
            .O(N__8420),
            .I(N__8414));
    LocalMux I__1875 (
            .O(N__8417),
            .I(N__8408));
    Span4Mux_v I__1874 (
            .O(N__8414),
            .I(N__8408));
    InMux I__1873 (
            .O(N__8413),
            .I(N__8405));
    Span4Mux_h I__1872 (
            .O(N__8408),
            .I(N__8400));
    LocalMux I__1871 (
            .O(N__8405),
            .I(N__8400));
    Sp12to4 I__1870 (
            .O(N__8400),
            .I(N__8397));
    Span12Mux_v I__1869 (
            .O(N__8397),
            .I(N__8394));
    Odrv12 I__1868 (
            .O(N__8394),
            .I(SIZ_c_0));
    IoInMux I__1867 (
            .O(N__8391),
            .I(N__8388));
    LocalMux I__1866 (
            .O(N__8388),
            .I(N__8385));
    Span12Mux_s5_v I__1865 (
            .O(N__8385),
            .I(N__8382));
    Span12Mux_h I__1864 (
            .O(N__8382),
            .I(N__8379));
    Odrv12 I__1863 (
            .O(N__8379),
            .I(un1_UDSn_i_0_0));
    IoInMux I__1862 (
            .O(N__8376),
            .I(N__8373));
    LocalMux I__1861 (
            .O(N__8373),
            .I(N__8370));
    Span4Mux_s0_v I__1860 (
            .O(N__8370),
            .I(N__8367));
    Span4Mux_v I__1859 (
            .O(N__8367),
            .I(N__8364));
    Span4Mux_v I__1858 (
            .O(N__8364),
            .I(N__8361));
    Sp12to4 I__1857 (
            .O(N__8361),
            .I(N__8358));
    Odrv12 I__1856 (
            .O(N__8358),
            .I(RASn_c));
    IoInMux I__1855 (
            .O(N__8355),
            .I(N__8352));
    LocalMux I__1854 (
            .O(N__8352),
            .I(N__8349));
    Span4Mux_s2_v I__1853 (
            .O(N__8349),
            .I(N__8346));
    Sp12to4 I__1852 (
            .O(N__8346),
            .I(N__8343));
    Span12Mux_h I__1851 (
            .O(N__8343),
            .I(N__8340));
    Odrv12 I__1850 (
            .O(N__8340),
            .I(CRCSn_c));
    IoInMux I__1849 (
            .O(N__8337),
            .I(N__8334));
    LocalMux I__1848 (
            .O(N__8334),
            .I(N__8331));
    Span12Mux_s4_h I__1847 (
            .O(N__8331),
            .I(N__8328));
    Span12Mux_h I__1846 (
            .O(N__8328),
            .I(N__8325));
    Odrv12 I__1845 (
            .O(N__8325),
            .I(WEn_c));
    IoInMux I__1844 (
            .O(N__8322),
            .I(N__8319));
    LocalMux I__1843 (
            .O(N__8319),
            .I(N__8316));
    Span12Mux_s3_v I__1842 (
            .O(N__8316),
            .I(N__8313));
    Span12Mux_h I__1841 (
            .O(N__8313),
            .I(N__8310));
    Odrv12 I__1840 (
            .O(N__8310),
            .I(CASn_c));
    CascadeMux I__1839 (
            .O(N__8307),
            .I(N__8301));
    InMux I__1838 (
            .O(N__8306),
            .I(N__8297));
    InMux I__1837 (
            .O(N__8305),
            .I(N__8294));
    InMux I__1836 (
            .O(N__8304),
            .I(N__8291));
    InMux I__1835 (
            .O(N__8301),
            .I(N__8286));
    InMux I__1834 (
            .O(N__8300),
            .I(N__8286));
    LocalMux I__1833 (
            .O(N__8297),
            .I(N__8283));
    LocalMux I__1832 (
            .O(N__8294),
            .I(N__8279));
    LocalMux I__1831 (
            .O(N__8291),
            .I(N__8274));
    LocalMux I__1830 (
            .O(N__8286),
            .I(N__8274));
    Span4Mux_v I__1829 (
            .O(N__8283),
            .I(N__8271));
    InMux I__1828 (
            .O(N__8282),
            .I(N__8268));
    Span12Mux_h I__1827 (
            .O(N__8279),
            .I(N__8265));
    Span4Mux_v I__1826 (
            .O(N__8274),
            .I(N__8262));
    Span4Mux_v I__1825 (
            .O(N__8271),
            .I(N__8257));
    LocalMux I__1824 (
            .O(N__8268),
            .I(N__8257));
    Odrv12 I__1823 (
            .O(N__8265),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1822 (
            .O(N__8262),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1821 (
            .O(N__8257),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    InMux I__1820 (
            .O(N__8250),
            .I(N__8247));
    LocalMux I__1819 (
            .O(N__8247),
            .I(N__8243));
    InMux I__1818 (
            .O(N__8246),
            .I(N__8240));
    Span4Mux_h I__1817 (
            .O(N__8243),
            .I(N__8232));
    LocalMux I__1816 (
            .O(N__8240),
            .I(N__8232));
    CascadeMux I__1815 (
            .O(N__8239),
            .I(N__8228));
    CascadeMux I__1814 (
            .O(N__8238),
            .I(N__8225));
    CascadeMux I__1813 (
            .O(N__8237),
            .I(N__8222));
    Span4Mux_v I__1812 (
            .O(N__8232),
            .I(N__8216));
    InMux I__1811 (
            .O(N__8231),
            .I(N__8213));
    InMux I__1810 (
            .O(N__8228),
            .I(N__8208));
    InMux I__1809 (
            .O(N__8225),
            .I(N__8208));
    InMux I__1808 (
            .O(N__8222),
            .I(N__8200));
    InMux I__1807 (
            .O(N__8221),
            .I(N__8197));
    CascadeMux I__1806 (
            .O(N__8220),
            .I(N__8194));
    CascadeMux I__1805 (
            .O(N__8219),
            .I(N__8188));
    Sp12to4 I__1804 (
            .O(N__8216),
            .I(N__8180));
    LocalMux I__1803 (
            .O(N__8213),
            .I(N__8180));
    LocalMux I__1802 (
            .O(N__8208),
            .I(N__8180));
    InMux I__1801 (
            .O(N__8207),
            .I(N__8177));
    InMux I__1800 (
            .O(N__8206),
            .I(N__8174));
    InMux I__1799 (
            .O(N__8205),
            .I(N__8169));
    InMux I__1798 (
            .O(N__8204),
            .I(N__8169));
    InMux I__1797 (
            .O(N__8203),
            .I(N__8166));
    LocalMux I__1796 (
            .O(N__8200),
            .I(N__8159));
    LocalMux I__1795 (
            .O(N__8197),
            .I(N__8156));
    InMux I__1794 (
            .O(N__8194),
            .I(N__8151));
    InMux I__1793 (
            .O(N__8193),
            .I(N__8151));
    InMux I__1792 (
            .O(N__8192),
            .I(N__8148));
    InMux I__1791 (
            .O(N__8191),
            .I(N__8141));
    InMux I__1790 (
            .O(N__8188),
            .I(N__8141));
    InMux I__1789 (
            .O(N__8187),
            .I(N__8141));
    Span12Mux_h I__1788 (
            .O(N__8180),
            .I(N__8137));
    LocalMux I__1787 (
            .O(N__8177),
            .I(N__8132));
    LocalMux I__1786 (
            .O(N__8174),
            .I(N__8132));
    LocalMux I__1785 (
            .O(N__8169),
            .I(N__8127));
    LocalMux I__1784 (
            .O(N__8166),
            .I(N__8127));
    InMux I__1783 (
            .O(N__8165),
            .I(N__8118));
    InMux I__1782 (
            .O(N__8164),
            .I(N__8118));
    InMux I__1781 (
            .O(N__8163),
            .I(N__8118));
    InMux I__1780 (
            .O(N__8162),
            .I(N__8118));
    Span4Mux_v I__1779 (
            .O(N__8159),
            .I(N__8107));
    Span4Mux_h I__1778 (
            .O(N__8156),
            .I(N__8107));
    LocalMux I__1777 (
            .O(N__8151),
            .I(N__8107));
    LocalMux I__1776 (
            .O(N__8148),
            .I(N__8107));
    LocalMux I__1775 (
            .O(N__8141),
            .I(N__8107));
    InMux I__1774 (
            .O(N__8140),
            .I(N__8104));
    Odrv12 I__1773 (
            .O(N__8137),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1772 (
            .O(N__8132),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__1771 (
            .O(N__8127),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1770 (
            .O(N__8118),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1769 (
            .O(N__8107),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1768 (
            .O(N__8104),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    CascadeMux I__1767 (
            .O(N__8091),
            .I(N__8087));
    InMux I__1766 (
            .O(N__8090),
            .I(N__8084));
    InMux I__1765 (
            .O(N__8087),
            .I(N__8081));
    LocalMux I__1764 (
            .O(N__8084),
            .I(N__8075));
    LocalMux I__1763 (
            .O(N__8081),
            .I(N__8075));
    InMux I__1762 (
            .O(N__8080),
            .I(N__8072));
    Span12Mux_v I__1761 (
            .O(N__8075),
            .I(N__8068));
    LocalMux I__1760 (
            .O(N__8072),
            .I(N__8065));
    InMux I__1759 (
            .O(N__8071),
            .I(N__8062));
    Odrv12 I__1758 (
            .O(N__8068),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1757 (
            .O(N__8065),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1756 (
            .O(N__8062),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    InMux I__1755 (
            .O(N__8055),
            .I(N__8052));
    LocalMux I__1754 (
            .O(N__8052),
            .I(N__8049));
    Span4Mux_v I__1753 (
            .O(N__8049),
            .I(N__8043));
    InMux I__1752 (
            .O(N__8048),
            .I(N__8040));
    InMux I__1751 (
            .O(N__8047),
            .I(N__8035));
    InMux I__1750 (
            .O(N__8046),
            .I(N__8035));
    Sp12to4 I__1749 (
            .O(N__8043),
            .I(N__8029));
    LocalMux I__1748 (
            .O(N__8040),
            .I(N__8029));
    LocalMux I__1747 (
            .O(N__8035),
            .I(N__8025));
    CascadeMux I__1746 (
            .O(N__8034),
            .I(N__8022));
    Span12Mux_h I__1745 (
            .O(N__8029),
            .I(N__8019));
    InMux I__1744 (
            .O(N__8028),
            .I(N__8016));
    Span4Mux_h I__1743 (
            .O(N__8025),
            .I(N__8013));
    InMux I__1742 (
            .O(N__8022),
            .I(N__8010));
    Odrv12 I__1741 (
            .O(N__8019),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1740 (
            .O(N__8016),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1739 (
            .O(N__8013),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1738 (
            .O(N__8010),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1737 (
            .O(N__8001),
            .I(N__7998));
    LocalMux I__1736 (
            .O(N__7998),
            .I(N__7995));
    Span4Mux_s0_v I__1735 (
            .O(N__7995),
            .I(N__7992));
    Sp12to4 I__1734 (
            .O(N__7992),
            .I(N__7989));
    Span12Mux_h I__1733 (
            .O(N__7989),
            .I(N__7986));
    Odrv12 I__1732 (
            .O(N__7986),
            .I(CMA_c_10));
    InMux I__1731 (
            .O(N__7983),
            .I(N__7979));
    InMux I__1730 (
            .O(N__7982),
            .I(N__7976));
    LocalMux I__1729 (
            .O(N__7979),
            .I(N__7971));
    LocalMux I__1728 (
            .O(N__7976),
            .I(N__7971));
    Span4Mux_h I__1727 (
            .O(N__7971),
            .I(N__7966));
    InMux I__1726 (
            .O(N__7970),
            .I(N__7961));
    InMux I__1725 (
            .O(N__7969),
            .I(N__7961));
    Odrv4 I__1724 (
            .O(N__7966),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1723 (
            .O(N__7961),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    InMux I__1722 (
            .O(N__7956),
            .I(N__7950));
    InMux I__1721 (
            .O(N__7955),
            .I(N__7950));
    LocalMux I__1720 (
            .O(N__7950),
            .I(N__7947));
    Span4Mux_v I__1719 (
            .O(N__7947),
            .I(N__7944));
    Sp12to4 I__1718 (
            .O(N__7944),
            .I(N__7941));
    Span12Mux_h I__1717 (
            .O(N__7941),
            .I(N__7938));
    Span12Mux_v I__1716 (
            .O(N__7938),
            .I(N__7935));
    Odrv12 I__1715 (
            .O(N__7935),
            .I(A_c_14));
    CascadeMux I__1714 (
            .O(N__7932),
            .I(N__7927));
    CascadeMux I__1713 (
            .O(N__7931),
            .I(N__7916));
    InMux I__1712 (
            .O(N__7930),
            .I(N__7906));
    InMux I__1711 (
            .O(N__7927),
            .I(N__7906));
    InMux I__1710 (
            .O(N__7926),
            .I(N__7906));
    InMux I__1709 (
            .O(N__7925),
            .I(N__7903));
    CascadeMux I__1708 (
            .O(N__7924),
            .I(N__7899));
    CascadeMux I__1707 (
            .O(N__7923),
            .I(N__7896));
    CascadeMux I__1706 (
            .O(N__7922),
            .I(N__7893));
    CascadeMux I__1705 (
            .O(N__7921),
            .I(N__7890));
    InMux I__1704 (
            .O(N__7920),
            .I(N__7885));
    InMux I__1703 (
            .O(N__7919),
            .I(N__7882));
    InMux I__1702 (
            .O(N__7916),
            .I(N__7877));
    InMux I__1701 (
            .O(N__7915),
            .I(N__7874));
    InMux I__1700 (
            .O(N__7914),
            .I(N__7869));
    InMux I__1699 (
            .O(N__7913),
            .I(N__7869));
    LocalMux I__1698 (
            .O(N__7906),
            .I(N__7864));
    LocalMux I__1697 (
            .O(N__7903),
            .I(N__7864));
    CascadeMux I__1696 (
            .O(N__7902),
            .I(N__7861));
    InMux I__1695 (
            .O(N__7899),
            .I(N__7858));
    InMux I__1694 (
            .O(N__7896),
            .I(N__7849));
    InMux I__1693 (
            .O(N__7893),
            .I(N__7849));
    InMux I__1692 (
            .O(N__7890),
            .I(N__7849));
    InMux I__1691 (
            .O(N__7889),
            .I(N__7846));
    InMux I__1690 (
            .O(N__7888),
            .I(N__7841));
    LocalMux I__1689 (
            .O(N__7885),
            .I(N__7838));
    LocalMux I__1688 (
            .O(N__7882),
            .I(N__7835));
    InMux I__1687 (
            .O(N__7881),
            .I(N__7830));
    InMux I__1686 (
            .O(N__7880),
            .I(N__7830));
    LocalMux I__1685 (
            .O(N__7877),
            .I(N__7825));
    LocalMux I__1684 (
            .O(N__7874),
            .I(N__7825));
    LocalMux I__1683 (
            .O(N__7869),
            .I(N__7822));
    Span4Mux_v I__1682 (
            .O(N__7864),
            .I(N__7819));
    InMux I__1681 (
            .O(N__7861),
            .I(N__7816));
    LocalMux I__1680 (
            .O(N__7858),
            .I(N__7813));
    InMux I__1679 (
            .O(N__7857),
            .I(N__7808));
    InMux I__1678 (
            .O(N__7856),
            .I(N__7808));
    LocalMux I__1677 (
            .O(N__7849),
            .I(N__7803));
    LocalMux I__1676 (
            .O(N__7846),
            .I(N__7803));
    InMux I__1675 (
            .O(N__7845),
            .I(N__7798));
    InMux I__1674 (
            .O(N__7844),
            .I(N__7798));
    LocalMux I__1673 (
            .O(N__7841),
            .I(N__7793));
    Span4Mux_h I__1672 (
            .O(N__7838),
            .I(N__7793));
    Span4Mux_h I__1671 (
            .O(N__7835),
            .I(N__7784));
    LocalMux I__1670 (
            .O(N__7830),
            .I(N__7784));
    Span4Mux_v I__1669 (
            .O(N__7825),
            .I(N__7784));
    Span4Mux_h I__1668 (
            .O(N__7822),
            .I(N__7784));
    Odrv4 I__1667 (
            .O(N__7819),
            .I(CPU_CYCLEm));
    LocalMux I__1666 (
            .O(N__7816),
            .I(CPU_CYCLEm));
    Odrv4 I__1665 (
            .O(N__7813),
            .I(CPU_CYCLEm));
    LocalMux I__1664 (
            .O(N__7808),
            .I(CPU_CYCLEm));
    Odrv4 I__1663 (
            .O(N__7803),
            .I(CPU_CYCLEm));
    LocalMux I__1662 (
            .O(N__7798),
            .I(CPU_CYCLEm));
    Odrv4 I__1661 (
            .O(N__7793),
            .I(CPU_CYCLEm));
    Odrv4 I__1660 (
            .O(N__7784),
            .I(CPU_CYCLEm));
    InMux I__1659 (
            .O(N__7767),
            .I(N__7764));
    LocalMux I__1658 (
            .O(N__7764),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    InMux I__1657 (
            .O(N__7761),
            .I(N__7758));
    LocalMux I__1656 (
            .O(N__7758),
            .I(N__7755));
    Odrv4 I__1655 (
            .O(N__7755),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ));
    InMux I__1654 (
            .O(N__7752),
            .I(N__7748));
    InMux I__1653 (
            .O(N__7751),
            .I(N__7745));
    LocalMux I__1652 (
            .O(N__7748),
            .I(N__7740));
    LocalMux I__1651 (
            .O(N__7745),
            .I(N__7740));
    Odrv4 I__1650 (
            .O(N__7740),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__1649 (
            .O(N__7737),
            .I(bfn_11_11_0_));
    InMux I__1648 (
            .O(N__7734),
            .I(N__7730));
    InMux I__1647 (
            .O(N__7733),
            .I(N__7727));
    LocalMux I__1646 (
            .O(N__7730),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    LocalMux I__1645 (
            .O(N__7727),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    InMux I__1644 (
            .O(N__7722),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__1643 (
            .O(N__7719),
            .I(N__7715));
    InMux I__1642 (
            .O(N__7718),
            .I(N__7712));
    LocalMux I__1641 (
            .O(N__7715),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    LocalMux I__1640 (
            .O(N__7712),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    InMux I__1639 (
            .O(N__7707),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__1638 (
            .O(N__7704),
            .I(N__7701));
    LocalMux I__1637 (
            .O(N__7701),
            .I(N__7697));
    InMux I__1636 (
            .O(N__7700),
            .I(N__7694));
    Span4Mux_h I__1635 (
            .O(N__7697),
            .I(N__7691));
    LocalMux I__1634 (
            .O(N__7694),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    Odrv4 I__1633 (
            .O(N__7691),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__1632 (
            .O(N__7686),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    CascadeMux I__1631 (
            .O(N__7683),
            .I(N__7679));
    InMux I__1630 (
            .O(N__7682),
            .I(N__7676));
    InMux I__1629 (
            .O(N__7679),
            .I(N__7673));
    LocalMux I__1628 (
            .O(N__7676),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__1627 (
            .O(N__7673),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__1626 (
            .O(N__7668),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__1625 (
            .O(N__7665),
            .I(N__7661));
    InMux I__1624 (
            .O(N__7664),
            .I(N__7658));
    LocalMux I__1623 (
            .O(N__7661),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__1622 (
            .O(N__7658),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__1621 (
            .O(N__7653),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__1620 (
            .O(N__7650),
            .I(N__7647));
    LocalMux I__1619 (
            .O(N__7647),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i ));
    InMux I__1618 (
            .O(N__7644),
            .I(N__7641));
    LocalMux I__1617 (
            .O(N__7641),
            .I(N__7638));
    Span4Mux_h I__1616 (
            .O(N__7638),
            .I(N__7635));
    Odrv4 I__1615 (
            .O(N__7635),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__1614 (
            .O(N__7632),
            .I(N__7629));
    LocalMux I__1613 (
            .O(N__7629),
            .I(N__7626));
    Span12Mux_s4_v I__1612 (
            .O(N__7626),
            .I(N__7623));
    Odrv12 I__1611 (
            .O(N__7623),
            .I(CMA_c_2));
    IoInMux I__1610 (
            .O(N__7620),
            .I(N__7617));
    LocalMux I__1609 (
            .O(N__7617),
            .I(N__7614));
    IoSpan4Mux I__1608 (
            .O(N__7614),
            .I(N__7611));
    Sp12to4 I__1607 (
            .O(N__7611),
            .I(N__7608));
    Span12Mux_s7_h I__1606 (
            .O(N__7608),
            .I(N__7605));
    Span12Mux_v I__1605 (
            .O(N__7605),
            .I(N__7602));
    Odrv12 I__1604 (
            .O(N__7602),
            .I(CMA_c_7));
    InMux I__1603 (
            .O(N__7599),
            .I(N__7596));
    LocalMux I__1602 (
            .O(N__7596),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    IoInMux I__1601 (
            .O(N__7593),
            .I(N__7590));
    LocalMux I__1600 (
            .O(N__7590),
            .I(N__7587));
    IoSpan4Mux I__1599 (
            .O(N__7587),
            .I(N__7584));
    IoSpan4Mux I__1598 (
            .O(N__7584),
            .I(N__7581));
    Span4Mux_s3_h I__1597 (
            .O(N__7581),
            .I(N__7578));
    Sp12to4 I__1596 (
            .O(N__7578),
            .I(N__7575));
    Span12Mux_h I__1595 (
            .O(N__7575),
            .I(N__7572));
    Odrv12 I__1594 (
            .O(N__7572),
            .I(CMA_c_5));
    InMux I__1593 (
            .O(N__7569),
            .I(N__7566));
    LocalMux I__1592 (
            .O(N__7566),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__1591 (
            .O(N__7563),
            .I(N__7560));
    LocalMux I__1590 (
            .O(N__7560),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    InMux I__1589 (
            .O(N__7557),
            .I(N__7554));
    LocalMux I__1588 (
            .O(N__7554),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    InMux I__1587 (
            .O(N__7551),
            .I(N__7548));
    LocalMux I__1586 (
            .O(N__7548),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__1585 (
            .O(N__7545),
            .I(N__7542));
    LocalMux I__1584 (
            .O(N__7542),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    InMux I__1583 (
            .O(N__7539),
            .I(N__7536));
    LocalMux I__1582 (
            .O(N__7536),
            .I(N__7533));
    Odrv12 I__1581 (
            .O(N__7533),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    InMux I__1580 (
            .O(N__7530),
            .I(N__7527));
    LocalMux I__1579 (
            .O(N__7527),
            .I(N__7524));
    Span4Mux_v I__1578 (
            .O(N__7524),
            .I(N__7521));
    Sp12to4 I__1577 (
            .O(N__7521),
            .I(N__7518));
    Span12Mux_h I__1576 (
            .O(N__7518),
            .I(N__7515));
    Odrv12 I__1575 (
            .O(N__7515),
            .I(A_c_10));
    InMux I__1574 (
            .O(N__7512),
            .I(N__7509));
    LocalMux I__1573 (
            .O(N__7509),
            .I(N__7506));
    Span12Mux_v I__1572 (
            .O(N__7506),
            .I(N__7503));
    Span12Mux_h I__1571 (
            .O(N__7503),
            .I(N__7500));
    Odrv12 I__1570 (
            .O(N__7500),
            .I(A_c_3));
    InMux I__1569 (
            .O(N__7497),
            .I(N__7494));
    LocalMux I__1568 (
            .O(N__7494),
            .I(N__7491));
    Odrv4 I__1567 (
            .O(N__7491),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ));
    InMux I__1566 (
            .O(N__7488),
            .I(N__7485));
    LocalMux I__1565 (
            .O(N__7485),
            .I(N__7482));
    Span12Mux_v I__1564 (
            .O(N__7482),
            .I(N__7479));
    Span12Mux_h I__1563 (
            .O(N__7479),
            .I(N__7476));
    Odrv12 I__1562 (
            .O(N__7476),
            .I(A_c_12));
    InMux I__1561 (
            .O(N__7473),
            .I(N__7470));
    LocalMux I__1560 (
            .O(N__7470),
            .I(N__7467));
    Span4Mux_h I__1559 (
            .O(N__7467),
            .I(N__7464));
    Span4Mux_v I__1558 (
            .O(N__7464),
            .I(N__7461));
    Sp12to4 I__1557 (
            .O(N__7461),
            .I(N__7458));
    Odrv12 I__1556 (
            .O(N__7458),
            .I(A_c_5));
    InMux I__1555 (
            .O(N__7455),
            .I(N__7452));
    LocalMux I__1554 (
            .O(N__7452),
            .I(N__7449));
    Span4Mux_v I__1553 (
            .O(N__7449),
            .I(N__7446));
    Sp12to4 I__1552 (
            .O(N__7446),
            .I(N__7443));
    Span12Mux_h I__1551 (
            .O(N__7443),
            .I(N__7440));
    Span12Mux_v I__1550 (
            .O(N__7440),
            .I(N__7437));
    Odrv12 I__1549 (
            .O(N__7437),
            .I(A_c_2));
    InMux I__1548 (
            .O(N__7434),
            .I(N__7431));
    LocalMux I__1547 (
            .O(N__7431),
            .I(N__7428));
    Span12Mux_h I__1546 (
            .O(N__7428),
            .I(N__7425));
    Odrv12 I__1545 (
            .O(N__7425),
            .I(A_c_9));
    InMux I__1544 (
            .O(N__7422),
            .I(N__7419));
    LocalMux I__1543 (
            .O(N__7419),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    InMux I__1542 (
            .O(N__7416),
            .I(N__7413));
    LocalMux I__1541 (
            .O(N__7413),
            .I(N__7410));
    Sp12to4 I__1540 (
            .O(N__7410),
            .I(N__7407));
    Span12Mux_v I__1539 (
            .O(N__7407),
            .I(N__7404));
    Span12Mux_h I__1538 (
            .O(N__7404),
            .I(N__7401));
    Odrv12 I__1537 (
            .O(N__7401),
            .I(A_c_17));
    IoInMux I__1536 (
            .O(N__7398),
            .I(N__7395));
    LocalMux I__1535 (
            .O(N__7395),
            .I(N__7392));
    IoSpan4Mux I__1534 (
            .O(N__7392),
            .I(N__7389));
    IoSpan4Mux I__1533 (
            .O(N__7389),
            .I(N__7386));
    Span4Mux_s2_h I__1532 (
            .O(N__7386),
            .I(N__7383));
    Sp12to4 I__1531 (
            .O(N__7383),
            .I(N__7380));
    Span12Mux_s9_h I__1530 (
            .O(N__7380),
            .I(N__7377));
    Odrv12 I__1529 (
            .O(N__7377),
            .I(CMA_c_8));
    InMux I__1528 (
            .O(N__7374),
            .I(N__7371));
    LocalMux I__1527 (
            .O(N__7371),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__1526 (
            .O(N__7368),
            .I(N__7365));
    LocalMux I__1525 (
            .O(N__7365),
            .I(N__7362));
    Span12Mux_s5_h I__1524 (
            .O(N__7362),
            .I(N__7359));
    Span12Mux_h I__1523 (
            .O(N__7359),
            .I(N__7356));
    Odrv12 I__1522 (
            .O(N__7356),
            .I(CMA_c_6));
    IoInMux I__1521 (
            .O(N__7353),
            .I(N__7350));
    LocalMux I__1520 (
            .O(N__7350),
            .I(N__7347));
    Span4Mux_s3_v I__1519 (
            .O(N__7347),
            .I(N__7344));
    Span4Mux_v I__1518 (
            .O(N__7344),
            .I(N__7341));
    Span4Mux_v I__1517 (
            .O(N__7341),
            .I(N__7338));
    Span4Mux_h I__1516 (
            .O(N__7338),
            .I(N__7335));
    Odrv4 I__1515 (
            .O(N__7335),
            .I(CMA_c_0));
    InMux I__1514 (
            .O(N__7332),
            .I(N__7329));
    LocalMux I__1513 (
            .O(N__7329),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    InMux I__1512 (
            .O(N__7326),
            .I(N__7323));
    LocalMux I__1511 (
            .O(N__7323),
            .I(N__7320));
    Span4Mux_h I__1510 (
            .O(N__7320),
            .I(N__7317));
    Span4Mux_v I__1509 (
            .O(N__7317),
            .I(N__7314));
    Sp12to4 I__1508 (
            .O(N__7314),
            .I(N__7311));
    Odrv12 I__1507 (
            .O(N__7311),
            .I(A_c_7));
    CascadeMux I__1506 (
            .O(N__7308),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ));
    InMux I__1505 (
            .O(N__7305),
            .I(N__7302));
    LocalMux I__1504 (
            .O(N__7302),
            .I(\U712_CHIP_RAM.N_289 ));
    InMux I__1503 (
            .O(N__7299),
            .I(N__7296));
    LocalMux I__1502 (
            .O(N__7296),
            .I(N__7293));
    Odrv4 I__1501 (
            .O(N__7293),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    InMux I__1500 (
            .O(N__7290),
            .I(N__7287));
    LocalMux I__1499 (
            .O(N__7287),
            .I(N__7281));
    InMux I__1498 (
            .O(N__7286),
            .I(N__7276));
    InMux I__1497 (
            .O(N__7285),
            .I(N__7276));
    InMux I__1496 (
            .O(N__7284),
            .I(N__7272));
    Span4Mux_h I__1495 (
            .O(N__7281),
            .I(N__7269));
    LocalMux I__1494 (
            .O(N__7276),
            .I(N__7266));
    InMux I__1493 (
            .O(N__7275),
            .I(N__7263));
    LocalMux I__1492 (
            .O(N__7272),
            .I(\U712_CHIP_RAM.N_342 ));
    Odrv4 I__1491 (
            .O(N__7269),
            .I(\U712_CHIP_RAM.N_342 ));
    Odrv4 I__1490 (
            .O(N__7266),
            .I(\U712_CHIP_RAM.N_342 ));
    LocalMux I__1489 (
            .O(N__7263),
            .I(\U712_CHIP_RAM.N_342 ));
    CascadeMux I__1488 (
            .O(N__7254),
            .I(N__7247));
    CascadeMux I__1487 (
            .O(N__7253),
            .I(N__7240));
    CascadeMux I__1486 (
            .O(N__7252),
            .I(N__7234));
    CascadeMux I__1485 (
            .O(N__7251),
            .I(N__7231));
    InMux I__1484 (
            .O(N__7250),
            .I(N__7227));
    InMux I__1483 (
            .O(N__7247),
            .I(N__7224));
    InMux I__1482 (
            .O(N__7246),
            .I(N__7221));
    InMux I__1481 (
            .O(N__7245),
            .I(N__7218));
    InMux I__1480 (
            .O(N__7244),
            .I(N__7209));
    InMux I__1479 (
            .O(N__7243),
            .I(N__7209));
    InMux I__1478 (
            .O(N__7240),
            .I(N__7209));
    InMux I__1477 (
            .O(N__7239),
            .I(N__7204));
    InMux I__1476 (
            .O(N__7238),
            .I(N__7204));
    InMux I__1475 (
            .O(N__7237),
            .I(N__7197));
    InMux I__1474 (
            .O(N__7234),
            .I(N__7197));
    InMux I__1473 (
            .O(N__7231),
            .I(N__7197));
    InMux I__1472 (
            .O(N__7230),
            .I(N__7194));
    LocalMux I__1471 (
            .O(N__7227),
            .I(N__7191));
    LocalMux I__1470 (
            .O(N__7224),
            .I(N__7184));
    LocalMux I__1469 (
            .O(N__7221),
            .I(N__7184));
    LocalMux I__1468 (
            .O(N__7218),
            .I(N__7184));
    InMux I__1467 (
            .O(N__7217),
            .I(N__7181));
    InMux I__1466 (
            .O(N__7216),
            .I(N__7174));
    LocalMux I__1465 (
            .O(N__7209),
            .I(N__7169));
    LocalMux I__1464 (
            .O(N__7204),
            .I(N__7169));
    LocalMux I__1463 (
            .O(N__7197),
            .I(N__7164));
    LocalMux I__1462 (
            .O(N__7194),
            .I(N__7164));
    Span4Mux_v I__1461 (
            .O(N__7191),
            .I(N__7157));
    Span4Mux_v I__1460 (
            .O(N__7184),
            .I(N__7157));
    LocalMux I__1459 (
            .O(N__7181),
            .I(N__7157));
    InMux I__1458 (
            .O(N__7180),
            .I(N__7154));
    InMux I__1457 (
            .O(N__7179),
            .I(N__7149));
    InMux I__1456 (
            .O(N__7178),
            .I(N__7149));
    InMux I__1455 (
            .O(N__7177),
            .I(N__7146));
    LocalMux I__1454 (
            .O(N__7174),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1453 (
            .O(N__7169),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1452 (
            .O(N__7164),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1451 (
            .O(N__7157),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1450 (
            .O(N__7154),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1449 (
            .O(N__7149),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1448 (
            .O(N__7146),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__1447 (
            .O(N__7131),
            .I(N__7125));
    InMux I__1446 (
            .O(N__7130),
            .I(N__7122));
    InMux I__1445 (
            .O(N__7129),
            .I(N__7119));
    InMux I__1444 (
            .O(N__7128),
            .I(N__7116));
    LocalMux I__1443 (
            .O(N__7125),
            .I(N__7109));
    LocalMux I__1442 (
            .O(N__7122),
            .I(N__7104));
    LocalMux I__1441 (
            .O(N__7119),
            .I(N__7104));
    LocalMux I__1440 (
            .O(N__7116),
            .I(N__7101));
    InMux I__1439 (
            .O(N__7115),
            .I(N__7098));
    InMux I__1438 (
            .O(N__7114),
            .I(N__7092));
    InMux I__1437 (
            .O(N__7113),
            .I(N__7092));
    InMux I__1436 (
            .O(N__7112),
            .I(N__7089));
    Span4Mux_h I__1435 (
            .O(N__7109),
            .I(N__7086));
    Span4Mux_h I__1434 (
            .O(N__7104),
            .I(N__7083));
    Span4Mux_h I__1433 (
            .O(N__7101),
            .I(N__7078));
    LocalMux I__1432 (
            .O(N__7098),
            .I(N__7078));
    InMux I__1431 (
            .O(N__7097),
            .I(N__7075));
    LocalMux I__1430 (
            .O(N__7092),
            .I(\U712_CHIP_RAM.N_208 ));
    LocalMux I__1429 (
            .O(N__7089),
            .I(\U712_CHIP_RAM.N_208 ));
    Odrv4 I__1428 (
            .O(N__7086),
            .I(\U712_CHIP_RAM.N_208 ));
    Odrv4 I__1427 (
            .O(N__7083),
            .I(\U712_CHIP_RAM.N_208 ));
    Odrv4 I__1426 (
            .O(N__7078),
            .I(\U712_CHIP_RAM.N_208 ));
    LocalMux I__1425 (
            .O(N__7075),
            .I(\U712_CHIP_RAM.N_208 ));
    CEMux I__1424 (
            .O(N__7062),
            .I(N__7059));
    LocalMux I__1423 (
            .O(N__7059),
            .I(N__7056));
    Span4Mux_h I__1422 (
            .O(N__7056),
            .I(N__7053));
    Odrv4 I__1421 (
            .O(N__7053),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0 ));
    CascadeMux I__1420 (
            .O(N__7050),
            .I(N__7045));
    InMux I__1419 (
            .O(N__7049),
            .I(N__7035));
    InMux I__1418 (
            .O(N__7048),
            .I(N__7032));
    InMux I__1417 (
            .O(N__7045),
            .I(N__7026));
    InMux I__1416 (
            .O(N__7044),
            .I(N__7022));
    InMux I__1415 (
            .O(N__7043),
            .I(N__7010));
    InMux I__1414 (
            .O(N__7042),
            .I(N__7010));
    InMux I__1413 (
            .O(N__7041),
            .I(N__7010));
    InMux I__1412 (
            .O(N__7040),
            .I(N__7010));
    InMux I__1411 (
            .O(N__7039),
            .I(N__7010));
    InMux I__1410 (
            .O(N__7038),
            .I(N__7005));
    LocalMux I__1409 (
            .O(N__7035),
            .I(N__7000));
    LocalMux I__1408 (
            .O(N__7032),
            .I(N__7000));
    InMux I__1407 (
            .O(N__7031),
            .I(N__6997));
    InMux I__1406 (
            .O(N__7030),
            .I(N__6992));
    InMux I__1405 (
            .O(N__7029),
            .I(N__6992));
    LocalMux I__1404 (
            .O(N__7026),
            .I(N__6987));
    InMux I__1403 (
            .O(N__7025),
            .I(N__6984));
    LocalMux I__1402 (
            .O(N__7022),
            .I(N__6981));
    InMux I__1401 (
            .O(N__7021),
            .I(N__6978));
    LocalMux I__1400 (
            .O(N__7010),
            .I(N__6975));
    InMux I__1399 (
            .O(N__7009),
            .I(N__6972));
    InMux I__1398 (
            .O(N__7008),
            .I(N__6969));
    LocalMux I__1397 (
            .O(N__7005),
            .I(N__6960));
    Span4Mux_v I__1396 (
            .O(N__7000),
            .I(N__6960));
    LocalMux I__1395 (
            .O(N__6997),
            .I(N__6960));
    LocalMux I__1394 (
            .O(N__6992),
            .I(N__6960));
    InMux I__1393 (
            .O(N__6991),
            .I(N__6955));
    InMux I__1392 (
            .O(N__6990),
            .I(N__6955));
    Span4Mux_v I__1391 (
            .O(N__6987),
            .I(N__6950));
    LocalMux I__1390 (
            .O(N__6984),
            .I(N__6950));
    Odrv4 I__1389 (
            .O(N__6981),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1388 (
            .O(N__6978),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1387 (
            .O(N__6975),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1386 (
            .O(N__6972),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1385 (
            .O(N__6969),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1384 (
            .O(N__6960),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1383 (
            .O(N__6955),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1382 (
            .O(N__6950),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    CascadeMux I__1381 (
            .O(N__6933),
            .I(N__6926));
    InMux I__1380 (
            .O(N__6932),
            .I(N__6921));
    InMux I__1379 (
            .O(N__6931),
            .I(N__6917));
    InMux I__1378 (
            .O(N__6930),
            .I(N__6914));
    InMux I__1377 (
            .O(N__6929),
            .I(N__6907));
    InMux I__1376 (
            .O(N__6926),
            .I(N__6900));
    InMux I__1375 (
            .O(N__6925),
            .I(N__6900));
    InMux I__1374 (
            .O(N__6924),
            .I(N__6900));
    LocalMux I__1373 (
            .O(N__6921),
            .I(N__6897));
    InMux I__1372 (
            .O(N__6920),
            .I(N__6894));
    LocalMux I__1371 (
            .O(N__6917),
            .I(N__6891));
    LocalMux I__1370 (
            .O(N__6914),
            .I(N__6888));
    InMux I__1369 (
            .O(N__6913),
            .I(N__6885));
    CascadeMux I__1368 (
            .O(N__6912),
            .I(N__6881));
    CascadeMux I__1367 (
            .O(N__6911),
            .I(N__6877));
    InMux I__1366 (
            .O(N__6910),
            .I(N__6874));
    LocalMux I__1365 (
            .O(N__6907),
            .I(N__6869));
    LocalMux I__1364 (
            .O(N__6900),
            .I(N__6869));
    Span4Mux_v I__1363 (
            .O(N__6897),
            .I(N__6858));
    LocalMux I__1362 (
            .O(N__6894),
            .I(N__6858));
    Span4Mux_v I__1361 (
            .O(N__6891),
            .I(N__6858));
    Span4Mux_h I__1360 (
            .O(N__6888),
            .I(N__6858));
    LocalMux I__1359 (
            .O(N__6885),
            .I(N__6858));
    InMux I__1358 (
            .O(N__6884),
            .I(N__6853));
    InMux I__1357 (
            .O(N__6881),
            .I(N__6853));
    InMux I__1356 (
            .O(N__6880),
            .I(N__6848));
    InMux I__1355 (
            .O(N__6877),
            .I(N__6848));
    LocalMux I__1354 (
            .O(N__6874),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1353 (
            .O(N__6869),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1352 (
            .O(N__6858),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1351 (
            .O(N__6853),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1350 (
            .O(N__6848),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1349 (
            .O(N__6837),
            .I(N__6834));
    LocalMux I__1348 (
            .O(N__6834),
            .I(N__6831));
    Span4Mux_h I__1347 (
            .O(N__6831),
            .I(N__6828));
    Odrv4 I__1346 (
            .O(N__6828),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_a3_0 ));
    InMux I__1345 (
            .O(N__6825),
            .I(N__6822));
    LocalMux I__1344 (
            .O(N__6822),
            .I(N__6819));
    Span12Mux_v I__1343 (
            .O(N__6819),
            .I(N__6816));
    Span12Mux_h I__1342 (
            .O(N__6816),
            .I(N__6813));
    Odrv12 I__1341 (
            .O(N__6813),
            .I(A_c_16));
    InMux I__1340 (
            .O(N__6810),
            .I(N__6807));
    LocalMux I__1339 (
            .O(N__6807),
            .I(N__6804));
    Span12Mux_v I__1338 (
            .O(N__6804),
            .I(N__6801));
    Span12Mux_h I__1337 (
            .O(N__6801),
            .I(N__6798));
    Odrv12 I__1336 (
            .O(N__6798),
            .I(A_c_18));
    InMux I__1335 (
            .O(N__6795),
            .I(N__6791));
    InMux I__1334 (
            .O(N__6794),
            .I(N__6788));
    LocalMux I__1333 (
            .O(N__6791),
            .I(\U712_CHIP_RAM.N_303 ));
    LocalMux I__1332 (
            .O(N__6788),
            .I(\U712_CHIP_RAM.N_303 ));
    InMux I__1331 (
            .O(N__6783),
            .I(N__6777));
    InMux I__1330 (
            .O(N__6782),
            .I(N__6770));
    InMux I__1329 (
            .O(N__6781),
            .I(N__6770));
    InMux I__1328 (
            .O(N__6780),
            .I(N__6770));
    LocalMux I__1327 (
            .O(N__6777),
            .I(\U712_CHIP_RAM.N_241 ));
    LocalMux I__1326 (
            .O(N__6770),
            .I(\U712_CHIP_RAM.N_241 ));
    InMux I__1325 (
            .O(N__6765),
            .I(N__6761));
    InMux I__1324 (
            .O(N__6764),
            .I(N__6758));
    LocalMux I__1323 (
            .O(N__6761),
            .I(N__6751));
    LocalMux I__1322 (
            .O(N__6758),
            .I(N__6748));
    InMux I__1321 (
            .O(N__6757),
            .I(N__6745));
    InMux I__1320 (
            .O(N__6756),
            .I(N__6742));
    InMux I__1319 (
            .O(N__6755),
            .I(N__6739));
    InMux I__1318 (
            .O(N__6754),
            .I(N__6736));
    Span4Mux_v I__1317 (
            .O(N__6751),
            .I(N__6727));
    Span4Mux_h I__1316 (
            .O(N__6748),
            .I(N__6727));
    LocalMux I__1315 (
            .O(N__6745),
            .I(N__6727));
    LocalMux I__1314 (
            .O(N__6742),
            .I(N__6727));
    LocalMux I__1313 (
            .O(N__6739),
            .I(N__6724));
    LocalMux I__1312 (
            .O(N__6736),
            .I(N__6720));
    Span4Mux_v I__1311 (
            .O(N__6727),
            .I(N__6717));
    Span4Mux_h I__1310 (
            .O(N__6724),
            .I(N__6714));
    InMux I__1309 (
            .O(N__6723),
            .I(N__6711));
    Odrv12 I__1308 (
            .O(N__6720),
            .I(DMA_CYCLEm));
    Odrv4 I__1307 (
            .O(N__6717),
            .I(DMA_CYCLEm));
    Odrv4 I__1306 (
            .O(N__6714),
            .I(DMA_CYCLEm));
    LocalMux I__1305 (
            .O(N__6711),
            .I(DMA_CYCLEm));
    InMux I__1304 (
            .O(N__6702),
            .I(N__6698));
    InMux I__1303 (
            .O(N__6701),
            .I(N__6695));
    LocalMux I__1302 (
            .O(N__6698),
            .I(N__6692));
    LocalMux I__1301 (
            .O(N__6695),
            .I(N__6689));
    Span4Mux_v I__1300 (
            .O(N__6692),
            .I(N__6685));
    Span4Mux_v I__1299 (
            .O(N__6689),
            .I(N__6682));
    InMux I__1298 (
            .O(N__6688),
            .I(N__6679));
    Span4Mux_v I__1297 (
            .O(N__6685),
            .I(N__6676));
    Span4Mux_v I__1296 (
            .O(N__6682),
            .I(N__6671));
    LocalMux I__1295 (
            .O(N__6679),
            .I(N__6671));
    Span4Mux_v I__1294 (
            .O(N__6676),
            .I(N__6668));
    Span4Mux_v I__1293 (
            .O(N__6671),
            .I(N__6665));
    Sp12to4 I__1292 (
            .O(N__6668),
            .I(N__6660));
    Sp12to4 I__1291 (
            .O(N__6665),
            .I(N__6660));
    Span12Mux_h I__1290 (
            .O(N__6660),
            .I(N__6657));
    Odrv12 I__1289 (
            .O(N__6657),
            .I(AWEn_c));
    InMux I__1288 (
            .O(N__6654),
            .I(N__6651));
    LocalMux I__1287 (
            .O(N__6651),
            .I(N__6646));
    InMux I__1286 (
            .O(N__6650),
            .I(N__6643));
    InMux I__1285 (
            .O(N__6649),
            .I(N__6640));
    Span4Mux_v I__1284 (
            .O(N__6646),
            .I(N__6632));
    LocalMux I__1283 (
            .O(N__6643),
            .I(N__6632));
    LocalMux I__1282 (
            .O(N__6640),
            .I(N__6632));
    InMux I__1281 (
            .O(N__6639),
            .I(N__6629));
    Span4Mux_v I__1280 (
            .O(N__6632),
            .I(N__6626));
    LocalMux I__1279 (
            .O(N__6629),
            .I(N__6623));
    Span4Mux_v I__1278 (
            .O(N__6626),
            .I(N__6618));
    Span4Mux_v I__1277 (
            .O(N__6623),
            .I(N__6618));
    Sp12to4 I__1276 (
            .O(N__6618),
            .I(N__6615));
    Span12Mux_h I__1275 (
            .O(N__6615),
            .I(N__6612));
    Odrv12 I__1274 (
            .O(N__6612),
            .I(RnW_c));
    IoInMux I__1273 (
            .O(N__6609),
            .I(N__6606));
    LocalMux I__1272 (
            .O(N__6606),
            .I(N__6603));
    IoSpan4Mux I__1271 (
            .O(N__6603),
            .I(N__6600));
    Sp12to4 I__1270 (
            .O(N__6600),
            .I(N__6597));
    Span12Mux_s7_h I__1269 (
            .O(N__6597),
            .I(N__6594));
    Span12Mux_h I__1268 (
            .O(N__6594),
            .I(N__6591));
    Odrv12 I__1267 (
            .O(N__6591),
            .I(N_256));
    InMux I__1266 (
            .O(N__6588),
            .I(N__6585));
    LocalMux I__1265 (
            .O(N__6585),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    IoInMux I__1264 (
            .O(N__6582),
            .I(N__6579));
    LocalMux I__1263 (
            .O(N__6579),
            .I(N__6576));
    IoSpan4Mux I__1262 (
            .O(N__6576),
            .I(N__6573));
    Span4Mux_s2_v I__1261 (
            .O(N__6573),
            .I(N__6570));
    Span4Mux_v I__1260 (
            .O(N__6570),
            .I(N__6567));
    Span4Mux_v I__1259 (
            .O(N__6567),
            .I(N__6563));
    InMux I__1258 (
            .O(N__6566),
            .I(N__6560));
    Odrv4 I__1257 (
            .O(N__6563),
            .I(CONSTANT_ONE_NET));
    LocalMux I__1256 (
            .O(N__6560),
            .I(CONSTANT_ONE_NET));
    InMux I__1255 (
            .O(N__6555),
            .I(N__6552));
    LocalMux I__1254 (
            .O(N__6552),
            .I(N__6549));
    Span4Mux_h I__1253 (
            .O(N__6549),
            .I(N__6546));
    Sp12to4 I__1252 (
            .O(N__6546),
            .I(N__6543));
    Span12Mux_v I__1251 (
            .O(N__6543),
            .I(N__6540));
    Odrv12 I__1250 (
            .O(N__6540),
            .I(A_c_19));
    IoInMux I__1249 (
            .O(N__6537),
            .I(N__6534));
    LocalMux I__1248 (
            .O(N__6534),
            .I(N__6531));
    IoSpan4Mux I__1247 (
            .O(N__6531),
            .I(N__6528));
    Span4Mux_s1_h I__1246 (
            .O(N__6528),
            .I(N__6525));
    Span4Mux_v I__1245 (
            .O(N__6525),
            .I(N__6522));
    Sp12to4 I__1244 (
            .O(N__6522),
            .I(N__6519));
    Span12Mux_s10_h I__1243 (
            .O(N__6519),
            .I(N__6516));
    Odrv12 I__1242 (
            .O(N__6516),
            .I(CMA_c_9));
    InMux I__1241 (
            .O(N__6513),
            .I(N__6510));
    LocalMux I__1240 (
            .O(N__6510),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    IoInMux I__1239 (
            .O(N__6507),
            .I(N__6504));
    LocalMux I__1238 (
            .O(N__6504),
            .I(N__6501));
    Span12Mux_s6_h I__1237 (
            .O(N__6501),
            .I(N__6498));
    Span12Mux_h I__1236 (
            .O(N__6498),
            .I(N__6495));
    Odrv12 I__1235 (
            .O(N__6495),
            .I(CMA_c_4));
    IoInMux I__1234 (
            .O(N__6492),
            .I(N__6489));
    LocalMux I__1233 (
            .O(N__6489),
            .I(N__6486));
    Span4Mux_s3_v I__1232 (
            .O(N__6486),
            .I(N__6483));
    Sp12to4 I__1231 (
            .O(N__6483),
            .I(N__6480));
    Span12Mux_h I__1230 (
            .O(N__6480),
            .I(N__6477));
    Odrv12 I__1229 (
            .O(N__6477),
            .I(CMA_c_1));
    InMux I__1228 (
            .O(N__6474),
            .I(N__6471));
    LocalMux I__1227 (
            .O(N__6471),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    InMux I__1226 (
            .O(N__6468),
            .I(N__6465));
    LocalMux I__1225 (
            .O(N__6465),
            .I(N__6462));
    Span4Mux_h I__1224 (
            .O(N__6462),
            .I(N__6458));
    InMux I__1223 (
            .O(N__6461),
            .I(N__6455));
    Odrv4 I__1222 (
            .O(N__6458),
            .I(DBR_SYNCZ0Z_0));
    LocalMux I__1221 (
            .O(N__6455),
            .I(DBR_SYNCZ0Z_0));
    CascadeMux I__1220 (
            .O(N__6450),
            .I(N__6447));
    InMux I__1219 (
            .O(N__6447),
            .I(N__6444));
    LocalMux I__1218 (
            .O(N__6444),
            .I(N__6441));
    Span4Mux_h I__1217 (
            .O(N__6441),
            .I(N__6437));
    InMux I__1216 (
            .O(N__6440),
            .I(N__6434));
    Odrv4 I__1215 (
            .O(N__6437),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1214 (
            .O(N__6434),
            .I(DBR_SYNCZ0Z_1));
    InMux I__1213 (
            .O(N__6429),
            .I(N__6426));
    LocalMux I__1212 (
            .O(N__6426),
            .I(N__6422));
    InMux I__1211 (
            .O(N__6425),
            .I(N__6419));
    Span4Mux_v I__1210 (
            .O(N__6422),
            .I(N__6413));
    LocalMux I__1209 (
            .O(N__6419),
            .I(N__6413));
    InMux I__1208 (
            .O(N__6418),
            .I(N__6410));
    Span4Mux_h I__1207 (
            .O(N__6413),
            .I(N__6407));
    LocalMux I__1206 (
            .O(N__6410),
            .I(N__6404));
    Odrv4 I__1205 (
            .O(N__6407),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    Odrv4 I__1204 (
            .O(N__6404),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__1203 (
            .O(N__6399),
            .I(N__6396));
    LocalMux I__1202 (
            .O(N__6396),
            .I(N__6392));
    InMux I__1201 (
            .O(N__6395),
            .I(N__6387));
    Span4Mux_h I__1200 (
            .O(N__6392),
            .I(N__6384));
    InMux I__1199 (
            .O(N__6391),
            .I(N__6379));
    InMux I__1198 (
            .O(N__6390),
            .I(N__6379));
    LocalMux I__1197 (
            .O(N__6387),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    Odrv4 I__1196 (
            .O(N__6384),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1195 (
            .O(N__6379),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    CascadeMux I__1194 (
            .O(N__6372),
            .I(N__6369));
    InMux I__1193 (
            .O(N__6369),
            .I(N__6365));
    InMux I__1192 (
            .O(N__6368),
            .I(N__6362));
    LocalMux I__1191 (
            .O(N__6365),
            .I(N__6359));
    LocalMux I__1190 (
            .O(N__6362),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    Odrv4 I__1189 (
            .O(N__6359),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__1188 (
            .O(N__6354),
            .I(N__6351));
    LocalMux I__1187 (
            .O(N__6351),
            .I(N__6348));
    Span4Mux_v I__1186 (
            .O(N__6348),
            .I(N__6345));
    Sp12to4 I__1185 (
            .O(N__6345),
            .I(N__6342));
    Span12Mux_h I__1184 (
            .O(N__6342),
            .I(N__6339));
    Odrv12 I__1183 (
            .O(N__6339),
            .I(RAS1n_c));
    InMux I__1182 (
            .O(N__6336),
            .I(N__6330));
    InMux I__1181 (
            .O(N__6335),
            .I(N__6330));
    LocalMux I__1180 (
            .O(N__6330),
            .I(\U712_CHIP_RAM.REFRESH_SYNCZ0Z_0 ));
    InMux I__1179 (
            .O(N__6327),
            .I(N__6324));
    LocalMux I__1178 (
            .O(N__6324),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0 ));
    CascadeMux I__1177 (
            .O(N__6321),
            .I(N__6318));
    InMux I__1176 (
            .O(N__6318),
            .I(N__6315));
    LocalMux I__1175 (
            .O(N__6315),
            .I(N__6312));
    Odrv4 I__1174 (
            .O(N__6312),
            .I(\U712_CHIP_RAM.N_301 ));
    InMux I__1173 (
            .O(N__6309),
            .I(N__6306));
    LocalMux I__1172 (
            .O(N__6306),
            .I(N__6303));
    Span4Mux_h I__1171 (
            .O(N__6303),
            .I(N__6300));
    Odrv4 I__1170 (
            .O(N__6300),
            .I(\U712_CHIP_RAM.N_243 ));
    InMux I__1169 (
            .O(N__6297),
            .I(N__6294));
    LocalMux I__1168 (
            .O(N__6294),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1 ));
    InMux I__1167 (
            .O(N__6291),
            .I(N__6288));
    LocalMux I__1166 (
            .O(N__6288),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0 ));
    CEMux I__1165 (
            .O(N__6285),
            .I(N__6281));
    CEMux I__1164 (
            .O(N__6284),
            .I(N__6278));
    LocalMux I__1163 (
            .O(N__6281),
            .I(N__6275));
    LocalMux I__1162 (
            .O(N__6278),
            .I(N__6272));
    Span4Mux_v I__1161 (
            .O(N__6275),
            .I(N__6269));
    Span4Mux_v I__1160 (
            .O(N__6272),
            .I(N__6266));
    Span4Mux_h I__1159 (
            .O(N__6269),
            .I(N__6263));
    Span4Mux_h I__1158 (
            .O(N__6266),
            .I(N__6260));
    Odrv4 I__1157 (
            .O(N__6263),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ));
    Odrv4 I__1156 (
            .O(N__6260),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ));
    CascadeMux I__1155 (
            .O(N__6255),
            .I(N__6249));
    CascadeMux I__1154 (
            .O(N__6254),
            .I(N__6246));
    CascadeMux I__1153 (
            .O(N__6253),
            .I(N__6242));
    InMux I__1152 (
            .O(N__6252),
            .I(N__6235));
    InMux I__1151 (
            .O(N__6249),
            .I(N__6226));
    InMux I__1150 (
            .O(N__6246),
            .I(N__6226));
    InMux I__1149 (
            .O(N__6245),
            .I(N__6226));
    InMux I__1148 (
            .O(N__6242),
            .I(N__6226));
    InMux I__1147 (
            .O(N__6241),
            .I(N__6221));
    InMux I__1146 (
            .O(N__6240),
            .I(N__6221));
    InMux I__1145 (
            .O(N__6239),
            .I(N__6217));
    InMux I__1144 (
            .O(N__6238),
            .I(N__6214));
    LocalMux I__1143 (
            .O(N__6235),
            .I(N__6209));
    LocalMux I__1142 (
            .O(N__6226),
            .I(N__6209));
    LocalMux I__1141 (
            .O(N__6221),
            .I(N__6206));
    InMux I__1140 (
            .O(N__6220),
            .I(N__6203));
    LocalMux I__1139 (
            .O(N__6217),
            .I(N__6197));
    LocalMux I__1138 (
            .O(N__6214),
            .I(N__6188));
    Span4Mux_v I__1137 (
            .O(N__6209),
            .I(N__6188));
    Span4Mux_v I__1136 (
            .O(N__6206),
            .I(N__6188));
    LocalMux I__1135 (
            .O(N__6203),
            .I(N__6188));
    InMux I__1134 (
            .O(N__6202),
            .I(N__6181));
    InMux I__1133 (
            .O(N__6201),
            .I(N__6181));
    InMux I__1132 (
            .O(N__6200),
            .I(N__6181));
    Odrv12 I__1131 (
            .O(N__6197),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1130 (
            .O(N__6188),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1129 (
            .O(N__6181),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__1128 (
            .O(N__6174),
            .I(N__6171));
    InMux I__1127 (
            .O(N__6171),
            .I(N__6167));
    InMux I__1126 (
            .O(N__6170),
            .I(N__6164));
    LocalMux I__1125 (
            .O(N__6167),
            .I(N__6158));
    LocalMux I__1124 (
            .O(N__6164),
            .I(N__6158));
    InMux I__1123 (
            .O(N__6163),
            .I(N__6155));
    Span4Mux_v I__1122 (
            .O(N__6158),
            .I(N__6152));
    LocalMux I__1121 (
            .O(N__6155),
            .I(\U712_CHIP_RAM.N_209 ));
    Odrv4 I__1120 (
            .O(N__6152),
            .I(\U712_CHIP_RAM.N_209 ));
    InMux I__1119 (
            .O(N__6147),
            .I(N__6144));
    LocalMux I__1118 (
            .O(N__6144),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_1 ));
    CascadeMux I__1117 (
            .O(N__6141),
            .I(N__6136));
    CascadeMux I__1116 (
            .O(N__6140),
            .I(N__6133));
    CascadeMux I__1115 (
            .O(N__6139),
            .I(N__6130));
    InMux I__1114 (
            .O(N__6136),
            .I(N__6122));
    InMux I__1113 (
            .O(N__6133),
            .I(N__6111));
    InMux I__1112 (
            .O(N__6130),
            .I(N__6111));
    CascadeMux I__1111 (
            .O(N__6129),
            .I(N__6108));
    InMux I__1110 (
            .O(N__6128),
            .I(N__6104));
    InMux I__1109 (
            .O(N__6127),
            .I(N__6099));
    InMux I__1108 (
            .O(N__6126),
            .I(N__6099));
    InMux I__1107 (
            .O(N__6125),
            .I(N__6096));
    LocalMux I__1106 (
            .O(N__6122),
            .I(N__6093));
    InMux I__1105 (
            .O(N__6121),
            .I(N__6090));
    InMux I__1104 (
            .O(N__6120),
            .I(N__6083));
    InMux I__1103 (
            .O(N__6119),
            .I(N__6083));
    InMux I__1102 (
            .O(N__6118),
            .I(N__6083));
    CascadeMux I__1101 (
            .O(N__6117),
            .I(N__6078));
    InMux I__1100 (
            .O(N__6116),
            .I(N__6074));
    LocalMux I__1099 (
            .O(N__6111),
            .I(N__6071));
    InMux I__1098 (
            .O(N__6108),
            .I(N__6068));
    InMux I__1097 (
            .O(N__6107),
            .I(N__6065));
    LocalMux I__1096 (
            .O(N__6104),
            .I(N__6060));
    LocalMux I__1095 (
            .O(N__6099),
            .I(N__6060));
    LocalMux I__1094 (
            .O(N__6096),
            .I(N__6055));
    Span4Mux_v I__1093 (
            .O(N__6093),
            .I(N__6055));
    LocalMux I__1092 (
            .O(N__6090),
            .I(N__6050));
    LocalMux I__1091 (
            .O(N__6083),
            .I(N__6050));
    InMux I__1090 (
            .O(N__6082),
            .I(N__6047));
    InMux I__1089 (
            .O(N__6081),
            .I(N__6044));
    InMux I__1088 (
            .O(N__6078),
            .I(N__6039));
    InMux I__1087 (
            .O(N__6077),
            .I(N__6039));
    LocalMux I__1086 (
            .O(N__6074),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1085 (
            .O(N__6071),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1084 (
            .O(N__6068),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1083 (
            .O(N__6065),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1082 (
            .O(N__6060),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1081 (
            .O(N__6055),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1080 (
            .O(N__6050),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1079 (
            .O(N__6047),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1078 (
            .O(N__6044),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1077 (
            .O(N__6039),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1076 (
            .O(N__6018),
            .I(N__6015));
    LocalMux I__1075 (
            .O(N__6015),
            .I(\U712_CHIP_RAM.N_227 ));
    InMux I__1074 (
            .O(N__6012),
            .I(N__6009));
    LocalMux I__1073 (
            .O(N__6009),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_2 ));
    CascadeMux I__1072 (
            .O(N__6006),
            .I(\U712_CHIP_RAM.N_342_cascade_ ));
    InMux I__1071 (
            .O(N__6003),
            .I(N__6000));
    LocalMux I__1070 (
            .O(N__6000),
            .I(N__5997));
    Span4Mux_v I__1069 (
            .O(N__5997),
            .I(N__5994));
    Span4Mux_v I__1068 (
            .O(N__5994),
            .I(N__5991));
    Span4Mux_h I__1067 (
            .O(N__5991),
            .I(N__5988));
    Sp12to4 I__1066 (
            .O(N__5988),
            .I(N__5985));
    Odrv12 I__1065 (
            .O(N__5985),
            .I(A_c_20));
    CascadeMux I__1064 (
            .O(N__5982),
            .I(\U712_CHIP_RAM.N_352_cascade_ ));
    InMux I__1063 (
            .O(N__5979),
            .I(N__5972));
    InMux I__1062 (
            .O(N__5978),
            .I(N__5972));
    InMux I__1061 (
            .O(N__5977),
            .I(N__5969));
    LocalMux I__1060 (
            .O(N__5972),
            .I(\U712_CHIP_RAM.N_395 ));
    LocalMux I__1059 (
            .O(N__5969),
            .I(\U712_CHIP_RAM.N_395 ));
    InMux I__1058 (
            .O(N__5964),
            .I(N__5959));
    InMux I__1057 (
            .O(N__5963),
            .I(N__5956));
    InMux I__1056 (
            .O(N__5962),
            .I(N__5953));
    LocalMux I__1055 (
            .O(N__5959),
            .I(\U712_CHIP_RAM.N_352 ));
    LocalMux I__1054 (
            .O(N__5956),
            .I(\U712_CHIP_RAM.N_352 ));
    LocalMux I__1053 (
            .O(N__5953),
            .I(\U712_CHIP_RAM.N_352 ));
    CascadeMux I__1052 (
            .O(N__5946),
            .I(\U712_CHIP_RAM.N_293_cascade_ ));
    InMux I__1051 (
            .O(N__5943),
            .I(N__5938));
    InMux I__1050 (
            .O(N__5942),
            .I(N__5935));
    InMux I__1049 (
            .O(N__5941),
            .I(N__5932));
    LocalMux I__1048 (
            .O(N__5938),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    LocalMux I__1047 (
            .O(N__5935),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    LocalMux I__1046 (
            .O(N__5932),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    CascadeMux I__1045 (
            .O(N__5925),
            .I(\U712_CHIP_RAM.N_99_cascade_ ));
    InMux I__1044 (
            .O(N__5922),
            .I(N__5918));
    InMux I__1043 (
            .O(N__5921),
            .I(N__5915));
    LocalMux I__1042 (
            .O(N__5918),
            .I(\U712_CHIP_RAM.N_290 ));
    LocalMux I__1041 (
            .O(N__5915),
            .I(\U712_CHIP_RAM.N_290 ));
    IoInMux I__1040 (
            .O(N__5910),
            .I(N__5907));
    LocalMux I__1039 (
            .O(N__5907),
            .I(N__5904));
    Span4Mux_s3_v I__1038 (
            .O(N__5904),
            .I(N__5901));
    Span4Mux_v I__1037 (
            .O(N__5901),
            .I(N__5898));
    Span4Mux_v I__1036 (
            .O(N__5898),
            .I(N__5895));
    Span4Mux_h I__1035 (
            .O(N__5895),
            .I(N__5891));
    InMux I__1034 (
            .O(N__5894),
            .I(N__5888));
    Odrv4 I__1033 (
            .O(N__5891),
            .I(BANK0_c));
    LocalMux I__1032 (
            .O(N__5888),
            .I(BANK0_c));
    InMux I__1031 (
            .O(N__5883),
            .I(N__5880));
    LocalMux I__1030 (
            .O(N__5880),
            .I(N__5876));
    InMux I__1029 (
            .O(N__5879),
            .I(N__5873));
    Span4Mux_v I__1028 (
            .O(N__5876),
            .I(N__5870));
    LocalMux I__1027 (
            .O(N__5873),
            .I(N__5867));
    Span4Mux_h I__1026 (
            .O(N__5870),
            .I(N__5862));
    Span4Mux_v I__1025 (
            .O(N__5867),
            .I(N__5862));
    Sp12to4 I__1024 (
            .O(N__5862),
            .I(N__5859));
    Span12Mux_h I__1023 (
            .O(N__5859),
            .I(N__5856));
    Span12Mux_v I__1022 (
            .O(N__5856),
            .I(N__5853));
    Odrv12 I__1021 (
            .O(N__5853),
            .I(TSn_c));
    InMux I__1020 (
            .O(N__5850),
            .I(N__5847));
    LocalMux I__1019 (
            .O(N__5847),
            .I(N__5844));
    Span4Mux_v I__1018 (
            .O(N__5844),
            .I(N__5841));
    Sp12to4 I__1017 (
            .O(N__5841),
            .I(N__5838));
    Span12Mux_h I__1016 (
            .O(N__5838),
            .I(N__5835));
    Span12Mux_v I__1015 (
            .O(N__5835),
            .I(N__5832));
    Odrv12 I__1014 (
            .O(N__5832),
            .I(RAMSPACEn_c));
    InMux I__1013 (
            .O(N__5829),
            .I(N__5824));
    InMux I__1012 (
            .O(N__5828),
            .I(N__5821));
    InMux I__1011 (
            .O(N__5827),
            .I(N__5818));
    LocalMux I__1010 (
            .O(N__5824),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__1009 (
            .O(N__5821),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__1008 (
            .O(N__5818),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__1007 (
            .O(N__5811),
            .I(N__5806));
    InMux I__1006 (
            .O(N__5810),
            .I(N__5803));
    InMux I__1005 (
            .O(N__5809),
            .I(N__5800));
    LocalMux I__1004 (
            .O(N__5806),
            .I(N__5797));
    LocalMux I__1003 (
            .O(N__5803),
            .I(N__5794));
    LocalMux I__1002 (
            .O(N__5800),
            .I(N__5789));
    Span4Mux_v I__1001 (
            .O(N__5797),
            .I(N__5786));
    Span4Mux_h I__1000 (
            .O(N__5794),
            .I(N__5783));
    InMux I__999 (
            .O(N__5793),
            .I(N__5780));
    InMux I__998 (
            .O(N__5792),
            .I(N__5777));
    Odrv4 I__997 (
            .O(N__5789),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__996 (
            .O(N__5786),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__995 (
            .O(N__5783),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__994 (
            .O(N__5780),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__993 (
            .O(N__5777),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    CascadeMux I__992 (
            .O(N__5766),
            .I(N__5763));
    InMux I__991 (
            .O(N__5763),
            .I(N__5751));
    InMux I__990 (
            .O(N__5762),
            .I(N__5751));
    InMux I__989 (
            .O(N__5761),
            .I(N__5746));
    InMux I__988 (
            .O(N__5760),
            .I(N__5746));
    InMux I__987 (
            .O(N__5759),
            .I(N__5741));
    InMux I__986 (
            .O(N__5758),
            .I(N__5738));
    CascadeMux I__985 (
            .O(N__5757),
            .I(N__5734));
    InMux I__984 (
            .O(N__5756),
            .I(N__5730));
    LocalMux I__983 (
            .O(N__5751),
            .I(N__5725));
    LocalMux I__982 (
            .O(N__5746),
            .I(N__5725));
    InMux I__981 (
            .O(N__5745),
            .I(N__5720));
    InMux I__980 (
            .O(N__5744),
            .I(N__5720));
    LocalMux I__979 (
            .O(N__5741),
            .I(N__5715));
    LocalMux I__978 (
            .O(N__5738),
            .I(N__5715));
    InMux I__977 (
            .O(N__5737),
            .I(N__5712));
    InMux I__976 (
            .O(N__5734),
            .I(N__5709));
    InMux I__975 (
            .O(N__5733),
            .I(N__5706));
    LocalMux I__974 (
            .O(N__5730),
            .I(N__5701));
    Span4Mux_h I__973 (
            .O(N__5725),
            .I(N__5701));
    LocalMux I__972 (
            .O(N__5720),
            .I(N__5698));
    Span4Mux_h I__971 (
            .O(N__5715),
            .I(N__5695));
    LocalMux I__970 (
            .O(N__5712),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__969 (
            .O(N__5709),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__968 (
            .O(N__5706),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__967 (
            .O(N__5701),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__966 (
            .O(N__5698),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__965 (
            .O(N__5695),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__964 (
            .O(N__5682),
            .I(N__5678));
    CascadeMux I__963 (
            .O(N__5681),
            .I(N__5672));
    LocalMux I__962 (
            .O(N__5678),
            .I(N__5669));
    InMux I__961 (
            .O(N__5677),
            .I(N__5662));
    InMux I__960 (
            .O(N__5676),
            .I(N__5662));
    InMux I__959 (
            .O(N__5675),
            .I(N__5662));
    InMux I__958 (
            .O(N__5672),
            .I(N__5659));
    Odrv4 I__957 (
            .O(N__5669),
            .I(\U712_CHIP_RAM.N_359 ));
    LocalMux I__956 (
            .O(N__5662),
            .I(\U712_CHIP_RAM.N_359 ));
    LocalMux I__955 (
            .O(N__5659),
            .I(\U712_CHIP_RAM.N_359 ));
    IoInMux I__954 (
            .O(N__5652),
            .I(N__5649));
    LocalMux I__953 (
            .O(N__5649),
            .I(N__5646));
    IoSpan4Mux I__952 (
            .O(N__5646),
            .I(N__5643));
    Span4Mux_s3_v I__951 (
            .O(N__5643),
            .I(N__5639));
    CascadeMux I__950 (
            .O(N__5642),
            .I(N__5636));
    Sp12to4 I__949 (
            .O(N__5639),
            .I(N__5633));
    InMux I__948 (
            .O(N__5636),
            .I(N__5630));
    Odrv12 I__947 (
            .O(N__5633),
            .I(DBDIR_c));
    LocalMux I__946 (
            .O(N__5630),
            .I(DBDIR_c));
    InMux I__945 (
            .O(N__5625),
            .I(N__5622));
    LocalMux I__944 (
            .O(N__5622),
            .I(N__5619));
    Sp12to4 I__943 (
            .O(N__5619),
            .I(N__5616));
    Span12Mux_v I__942 (
            .O(N__5616),
            .I(N__5613));
    Span12Mux_h I__941 (
            .O(N__5613),
            .I(N__5610));
    Odrv12 I__940 (
            .O(N__5610),
            .I(A_c_6));
    InMux I__939 (
            .O(N__5607),
            .I(N__5604));
    LocalMux I__938 (
            .O(N__5604),
            .I(N__5601));
    Span4Mux_v I__937 (
            .O(N__5601),
            .I(N__5598));
    Sp12to4 I__936 (
            .O(N__5598),
            .I(N__5595));
    Odrv12 I__935 (
            .O(N__5595),
            .I(A_c_13));
    CascadeMux I__934 (
            .O(N__5592),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ));
    InMux I__933 (
            .O(N__5589),
            .I(N__5586));
    LocalMux I__932 (
            .O(N__5586),
            .I(N__5583));
    Span4Mux_h I__931 (
            .O(N__5583),
            .I(N__5580));
    Odrv4 I__930 (
            .O(N__5580),
            .I(\U712_CHIP_RAM.N_257 ));
    InMux I__929 (
            .O(N__5577),
            .I(N__5572));
    InMux I__928 (
            .O(N__5576),
            .I(N__5569));
    CascadeMux I__927 (
            .O(N__5575),
            .I(N__5566));
    LocalMux I__926 (
            .O(N__5572),
            .I(N__5560));
    LocalMux I__925 (
            .O(N__5569),
            .I(N__5560));
    InMux I__924 (
            .O(N__5566),
            .I(N__5554));
    InMux I__923 (
            .O(N__5565),
            .I(N__5554));
    Span4Mux_v I__922 (
            .O(N__5560),
            .I(N__5551));
    InMux I__921 (
            .O(N__5559),
            .I(N__5548));
    LocalMux I__920 (
            .O(N__5554),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__919 (
            .O(N__5551),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__918 (
            .O(N__5548),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    InMux I__917 (
            .O(N__5541),
            .I(N__5538));
    LocalMux I__916 (
            .O(N__5538),
            .I(\U712_CHIP_RAM.N_205 ));
    CascadeMux I__915 (
            .O(N__5535),
            .I(\U712_CHIP_RAM.N_205_cascade_ ));
    InMux I__914 (
            .O(N__5532),
            .I(N__5523));
    InMux I__913 (
            .O(N__5531),
            .I(N__5523));
    InMux I__912 (
            .O(N__5530),
            .I(N__5520));
    InMux I__911 (
            .O(N__5529),
            .I(N__5517));
    InMux I__910 (
            .O(N__5528),
            .I(N__5514));
    LocalMux I__909 (
            .O(N__5523),
            .I(N__5511));
    LocalMux I__908 (
            .O(N__5520),
            .I(\U712_CHIP_RAM.N_216 ));
    LocalMux I__907 (
            .O(N__5517),
            .I(\U712_CHIP_RAM.N_216 ));
    LocalMux I__906 (
            .O(N__5514),
            .I(\U712_CHIP_RAM.N_216 ));
    Odrv4 I__905 (
            .O(N__5511),
            .I(\U712_CHIP_RAM.N_216 ));
    InMux I__904 (
            .O(N__5502),
            .I(N__5499));
    LocalMux I__903 (
            .O(N__5499),
            .I(\U712_CHIP_RAM.N_291 ));
    CascadeMux I__902 (
            .O(N__5496),
            .I(\U712_CHIP_RAM.N_291_cascade_ ));
    CascadeMux I__901 (
            .O(N__5493),
            .I(N__5490));
    InMux I__900 (
            .O(N__5490),
            .I(N__5487));
    LocalMux I__899 (
            .O(N__5487),
            .I(N__5484));
    Odrv4 I__898 (
            .O(N__5484),
            .I(\U712_CHIP_RAM.N_204 ));
    InMux I__897 (
            .O(N__5481),
            .I(N__5478));
    LocalMux I__896 (
            .O(N__5478),
            .I(N__5475));
    Span4Mux_h I__895 (
            .O(N__5475),
            .I(N__5472));
    Odrv4 I__894 (
            .O(N__5472),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ));
    IoInMux I__893 (
            .O(N__5469),
            .I(N__5466));
    LocalMux I__892 (
            .O(N__5466),
            .I(N__5462));
    InMux I__891 (
            .O(N__5465),
            .I(N__5459));
    Span4Mux_s3_v I__890 (
            .O(N__5462),
            .I(N__5455));
    LocalMux I__889 (
            .O(N__5459),
            .I(N__5452));
    InMux I__888 (
            .O(N__5458),
            .I(N__5449));
    Span4Mux_h I__887 (
            .O(N__5455),
            .I(N__5445));
    Span4Mux_h I__886 (
            .O(N__5452),
            .I(N__5440));
    LocalMux I__885 (
            .O(N__5449),
            .I(N__5440));
    InMux I__884 (
            .O(N__5448),
            .I(N__5437));
    Sp12to4 I__883 (
            .O(N__5445),
            .I(N__5433));
    Sp12to4 I__882 (
            .O(N__5440),
            .I(N__5428));
    LocalMux I__881 (
            .O(N__5437),
            .I(N__5428));
    InMux I__880 (
            .O(N__5436),
            .I(N__5425));
    Odrv12 I__879 (
            .O(N__5433),
            .I(DBENn_c));
    Odrv12 I__878 (
            .O(N__5428),
            .I(DBENn_c));
    LocalMux I__877 (
            .O(N__5425),
            .I(DBENn_c));
    InMux I__876 (
            .O(N__5418),
            .I(N__5415));
    LocalMux I__875 (
            .O(N__5415),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0 ));
    CascadeMux I__874 (
            .O(N__5412),
            .I(N__5409));
    InMux I__873 (
            .O(N__5409),
            .I(N__5404));
    InMux I__872 (
            .O(N__5408),
            .I(N__5401));
    InMux I__871 (
            .O(N__5407),
            .I(N__5398));
    LocalMux I__870 (
            .O(N__5404),
            .I(\U712_BYTE_ENABLE.N_319 ));
    LocalMux I__869 (
            .O(N__5401),
            .I(\U712_BYTE_ENABLE.N_319 ));
    LocalMux I__868 (
            .O(N__5398),
            .I(\U712_BYTE_ENABLE.N_319 ));
    InMux I__867 (
            .O(N__5391),
            .I(N__5388));
    LocalMux I__866 (
            .O(N__5388),
            .I(\U712_BYTE_ENABLE.N_322 ));
    CascadeMux I__865 (
            .O(N__5385),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_cascade_ ));
    InMux I__864 (
            .O(N__5382),
            .I(N__5378));
    InMux I__863 (
            .O(N__5381),
            .I(N__5375));
    LocalMux I__862 (
            .O(N__5378),
            .I(N__5372));
    LocalMux I__861 (
            .O(N__5375),
            .I(N__5368));
    Span4Mux_v I__860 (
            .O(N__5372),
            .I(N__5365));
    InMux I__859 (
            .O(N__5371),
            .I(N__5362));
    Span12Mux_h I__858 (
            .O(N__5368),
            .I(N__5359));
    Sp12to4 I__857 (
            .O(N__5365),
            .I(N__5354));
    LocalMux I__856 (
            .O(N__5362),
            .I(N__5354));
    Span12Mux_h I__855 (
            .O(N__5359),
            .I(N__5351));
    Span12Mux_h I__854 (
            .O(N__5354),
            .I(N__5348));
    Span12Mux_v I__853 (
            .O(N__5351),
            .I(N__5345));
    Span12Mux_v I__852 (
            .O(N__5348),
            .I(N__5342));
    Odrv12 I__851 (
            .O(N__5345),
            .I(CASLn_c));
    Odrv12 I__850 (
            .O(N__5342),
            .I(CASLn_c));
    IoInMux I__849 (
            .O(N__5337),
            .I(N__5334));
    LocalMux I__848 (
            .O(N__5334),
            .I(N__5331));
    IoSpan4Mux I__847 (
            .O(N__5331),
            .I(N__5328));
    Span4Mux_s0_h I__846 (
            .O(N__5328),
            .I(N__5325));
    Span4Mux_h I__845 (
            .O(N__5325),
            .I(N__5322));
    Sp12to4 I__844 (
            .O(N__5322),
            .I(N__5319));
    Span12Mux_v I__843 (
            .O(N__5319),
            .I(N__5316));
    Span12Mux_h I__842 (
            .O(N__5316),
            .I(N__5313));
    Odrv12 I__841 (
            .O(N__5313),
            .I(N_42_i));
    InMux I__840 (
            .O(N__5310),
            .I(N__5307));
    LocalMux I__839 (
            .O(N__5307),
            .I(N__5303));
    InMux I__838 (
            .O(N__5306),
            .I(N__5300));
    Span4Mux_v I__837 (
            .O(N__5303),
            .I(N__5296));
    LocalMux I__836 (
            .O(N__5300),
            .I(N__5293));
    InMux I__835 (
            .O(N__5299),
            .I(N__5290));
    Span4Mux_v I__834 (
            .O(N__5296),
            .I(N__5285));
    Span4Mux_v I__833 (
            .O(N__5293),
            .I(N__5285));
    LocalMux I__832 (
            .O(N__5290),
            .I(N__5282));
    Odrv4 I__831 (
            .O(N__5285),
            .I(REG_CYCLEm));
    Odrv4 I__830 (
            .O(N__5282),
            .I(REG_CYCLEm));
    IoInMux I__829 (
            .O(N__5277),
            .I(N__5274));
    LocalMux I__828 (
            .O(N__5274),
            .I(N__5271));
    IoSpan4Mux I__827 (
            .O(N__5271),
            .I(N__5268));
    IoSpan4Mux I__826 (
            .O(N__5268),
            .I(N__5265));
    Span4Mux_s3_v I__825 (
            .O(N__5265),
            .I(N__5262));
    Sp12to4 I__824 (
            .O(N__5262),
            .I(N__5259));
    Span12Mux_s11_v I__823 (
            .O(N__5259),
            .I(N__5256));
    Odrv12 I__822 (
            .O(N__5256),
            .I(DRDENn_c));
    InMux I__821 (
            .O(N__5253),
            .I(N__5250));
    LocalMux I__820 (
            .O(N__5250),
            .I(N__5247));
    Span4Mux_h I__819 (
            .O(N__5247),
            .I(N__5244));
    Sp12to4 I__818 (
            .O(N__5244),
            .I(N__5241));
    Span12Mux_v I__817 (
            .O(N__5241),
            .I(N__5238));
    Odrv12 I__816 (
            .O(N__5238),
            .I(A_c_8));
    InMux I__815 (
            .O(N__5235),
            .I(N__5232));
    LocalMux I__814 (
            .O(N__5232),
            .I(N__5229));
    Span4Mux_v I__813 (
            .O(N__5229),
            .I(N__5226));
    Span4Mux_v I__812 (
            .O(N__5226),
            .I(N__5223));
    Sp12to4 I__811 (
            .O(N__5223),
            .I(N__5220));
    Odrv12 I__810 (
            .O(N__5220),
            .I(A_c_15));
    IoInMux I__809 (
            .O(N__5217),
            .I(N__5214));
    LocalMux I__808 (
            .O(N__5214),
            .I(N__5211));
    IoSpan4Mux I__807 (
            .O(N__5211),
            .I(N__5208));
    Sp12to4 I__806 (
            .O(N__5208),
            .I(N__5205));
    Span12Mux_s7_h I__805 (
            .O(N__5205),
            .I(N__5202));
    Span12Mux_h I__804 (
            .O(N__5202),
            .I(N__5199));
    Odrv12 I__803 (
            .O(N__5199),
            .I(CLK_EN_c));
    InMux I__802 (
            .O(N__5196),
            .I(N__5193));
    LocalMux I__801 (
            .O(N__5193),
            .I(N__5190));
    Span4Mux_v I__800 (
            .O(N__5190),
            .I(N__5187));
    Odrv4 I__799 (
            .O(N__5187),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    InMux I__798 (
            .O(N__5184),
            .I(N__5181));
    LocalMux I__797 (
            .O(N__5181),
            .I(N__5178));
    Odrv4 I__796 (
            .O(N__5178),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0 ));
    CEMux I__795 (
            .O(N__5175),
            .I(N__5172));
    LocalMux I__794 (
            .O(N__5172),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0 ));
    CascadeMux I__793 (
            .O(N__5169),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_ ));
    InMux I__792 (
            .O(N__5166),
            .I(N__5161));
    InMux I__791 (
            .O(N__5165),
            .I(N__5158));
    InMux I__790 (
            .O(N__5164),
            .I(N__5155));
    LocalMux I__789 (
            .O(N__5161),
            .I(\U712_CHIP_RAM.N_393 ));
    LocalMux I__788 (
            .O(N__5158),
            .I(\U712_CHIP_RAM.N_393 ));
    LocalMux I__787 (
            .O(N__5155),
            .I(\U712_CHIP_RAM.N_393 ));
    InMux I__786 (
            .O(N__5148),
            .I(N__5145));
    LocalMux I__785 (
            .O(N__5145),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0 ));
    InMux I__784 (
            .O(N__5142),
            .I(N__5139));
    LocalMux I__783 (
            .O(N__5139),
            .I(\U712_CHIP_RAM.REFRESH_SYNCZ0Z_1 ));
    CascadeMux I__782 (
            .O(N__5136),
            .I(\U712_CHIP_RAM.N_227_cascade_ ));
    InMux I__781 (
            .O(N__5133),
            .I(N__5130));
    LocalMux I__780 (
            .O(N__5130),
            .I(N__5127));
    Odrv4 I__779 (
            .O(N__5127),
            .I(\U712_CHIP_RAM.N_226 ));
    InMux I__778 (
            .O(N__5124),
            .I(N__5121));
    LocalMux I__777 (
            .O(N__5121),
            .I(\U712_CHIP_RAM.N_245 ));
    CascadeMux I__776 (
            .O(N__5118),
            .I(\U712_CHIP_RAM.N_181_cascade_ ));
    InMux I__775 (
            .O(N__5115),
            .I(N__5112));
    LocalMux I__774 (
            .O(N__5112),
            .I(N__5109));
    Span4Mux_h I__773 (
            .O(N__5109),
            .I(N__5106));
    Odrv4 I__772 (
            .O(N__5106),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_a4_0_a3_0 ));
    CascadeMux I__771 (
            .O(N__5103),
            .I(\U712_CHIP_RAM.N_216_cascade_ ));
    InMux I__770 (
            .O(N__5100),
            .I(N__5097));
    LocalMux I__769 (
            .O(N__5097),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_0 ));
    InMux I__768 (
            .O(N__5094),
            .I(N__5091));
    LocalMux I__767 (
            .O(N__5091),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    CascadeMux I__766 (
            .O(N__5088),
            .I(N__5081));
    InMux I__765 (
            .O(N__5087),
            .I(N__5070));
    InMux I__764 (
            .O(N__5086),
            .I(N__5070));
    InMux I__763 (
            .O(N__5085),
            .I(N__5070));
    InMux I__762 (
            .O(N__5084),
            .I(N__5070));
    InMux I__761 (
            .O(N__5081),
            .I(N__5067));
    InMux I__760 (
            .O(N__5080),
            .I(N__5062));
    InMux I__759 (
            .O(N__5079),
            .I(N__5062));
    LocalMux I__758 (
            .O(N__5070),
            .I(N__5059));
    LocalMux I__757 (
            .O(N__5067),
            .I(\U712_CHIP_RAM.N_181 ));
    LocalMux I__756 (
            .O(N__5062),
            .I(\U712_CHIP_RAM.N_181 ));
    Odrv4 I__755 (
            .O(N__5059),
            .I(\U712_CHIP_RAM.N_181 ));
    CEMux I__754 (
            .O(N__5052),
            .I(N__5048));
    CEMux I__753 (
            .O(N__5051),
            .I(N__5045));
    LocalMux I__752 (
            .O(N__5048),
            .I(N__5040));
    LocalMux I__751 (
            .O(N__5045),
            .I(N__5040));
    Span4Mux_v I__750 (
            .O(N__5040),
            .I(N__5037));
    Span4Mux_h I__749 (
            .O(N__5037),
            .I(N__5034));
    Odrv4 I__748 (
            .O(N__5034),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    CascadeMux I__747 (
            .O(N__5031),
            .I(\U712_CHIP_RAM.N_204_cascade_ ));
    InMux I__746 (
            .O(N__5028),
            .I(N__5025));
    LocalMux I__745 (
            .O(N__5025),
            .I(N__5022));
    Odrv4 I__744 (
            .O(N__5022),
            .I(\U712_CHIP_RAM.N_279_1 ));
    CascadeMux I__743 (
            .O(N__5019),
            .I(\U712_CHIP_RAM.N_279_1_cascade_ ));
    InMux I__742 (
            .O(N__5016),
            .I(N__5012));
    InMux I__741 (
            .O(N__5015),
            .I(N__5009));
    LocalMux I__740 (
            .O(N__5012),
            .I(\U712_CHIP_RAM.N_398 ));
    LocalMux I__739 (
            .O(N__5009),
            .I(\U712_CHIP_RAM.N_398 ));
    CascadeMux I__738 (
            .O(N__5004),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_1_cascade_ ));
    IoInMux I__737 (
            .O(N__5001),
            .I(N__4998));
    LocalMux I__736 (
            .O(N__4998),
            .I(N__4995));
    Span12Mux_s5_v I__735 (
            .O(N__4995),
            .I(N__4992));
    Odrv12 I__734 (
            .O(N__4992),
            .I(VBENn_c));
    CascadeMux I__733 (
            .O(N__4989),
            .I(\U712_CHIP_RAM.N_209_cascade_ ));
    CascadeMux I__732 (
            .O(N__4986),
            .I(\U712_CHIP_RAM.N_359_cascade_ ));
    CascadeMux I__731 (
            .O(N__4983),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0_cascade_ ));
    CascadeMux I__730 (
            .O(N__4980),
            .I(\U712_CHIP_RAM.N_290_cascade_ ));
    InMux I__729 (
            .O(N__4977),
            .I(N__4972));
    InMux I__728 (
            .O(N__4976),
            .I(N__4969));
    CascadeMux I__727 (
            .O(N__4975),
            .I(N__4966));
    LocalMux I__726 (
            .O(N__4972),
            .I(N__4963));
    LocalMux I__725 (
            .O(N__4969),
            .I(N__4960));
    InMux I__724 (
            .O(N__4966),
            .I(N__4957));
    Span4Mux_v I__723 (
            .O(N__4963),
            .I(N__4952));
    Span4Mux_v I__722 (
            .O(N__4960),
            .I(N__4952));
    LocalMux I__721 (
            .O(N__4957),
            .I(N__4949));
    Sp12to4 I__720 (
            .O(N__4952),
            .I(N__4946));
    Span12Mux_v I__719 (
            .O(N__4949),
            .I(N__4943));
    Span12Mux_h I__718 (
            .O(N__4946),
            .I(N__4940));
    Span12Mux_h I__717 (
            .O(N__4943),
            .I(N__4935));
    Span12Mux_v I__716 (
            .O(N__4940),
            .I(N__4935));
    Odrv12 I__715 (
            .O(N__4935),
            .I(CASUn_c));
    CascadeMux I__714 (
            .O(N__4932),
            .I(\U712_BYTE_ENABLE.N_319_cascade_ ));
    IoInMux I__713 (
            .O(N__4929),
            .I(N__4926));
    LocalMux I__712 (
            .O(N__4926),
            .I(N__4923));
    IoSpan4Mux I__711 (
            .O(N__4923),
            .I(N__4920));
    Sp12to4 I__710 (
            .O(N__4920),
            .I(N__4917));
    Span12Mux_s9_h I__709 (
            .O(N__4917),
            .I(N__4914));
    Span12Mux_h I__708 (
            .O(N__4914),
            .I(N__4911));
    Odrv12 I__707 (
            .O(N__4911),
            .I(N_43_i));
    InMux I__706 (
            .O(N__4908),
            .I(N__4905));
    LocalMux I__705 (
            .O(N__4905),
            .I(N__4901));
    InMux I__704 (
            .O(N__4904),
            .I(N__4898));
    Span4Mux_v I__703 (
            .O(N__4901),
            .I(N__4895));
    LocalMux I__702 (
            .O(N__4898),
            .I(N__4892));
    Span4Mux_v I__701 (
            .O(N__4895),
            .I(N__4889));
    Span12Mux_h I__700 (
            .O(N__4892),
            .I(N__4886));
    Span4Mux_v I__699 (
            .O(N__4889),
            .I(N__4883));
    Span12Mux_v I__698 (
            .O(N__4886),
            .I(N__4880));
    Sp12to4 I__697 (
            .O(N__4883),
            .I(N__4877));
    Odrv12 I__696 (
            .O(N__4880),
            .I(SIZ_c_1));
    Odrv12 I__695 (
            .O(N__4877),
            .I(SIZ_c_1));
    InMux I__694 (
            .O(N__4872),
            .I(N__4869));
    LocalMux I__693 (
            .O(N__4869),
            .I(N__4865));
    InMux I__692 (
            .O(N__4868),
            .I(N__4862));
    Odrv4 I__691 (
            .O(N__4865),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0 ));
    LocalMux I__690 (
            .O(N__4862),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0 ));
    InMux I__689 (
            .O(N__4857),
            .I(N__4854));
    LocalMux I__688 (
            .O(N__4854),
            .I(\U712_BYTE_ENABLE.N_321 ));
    InMux I__687 (
            .O(N__4851),
            .I(N__4848));
    LocalMux I__686 (
            .O(N__4848),
            .I(N__4844));
    InMux I__685 (
            .O(N__4847),
            .I(N__4841));
    Span4Mux_v I__684 (
            .O(N__4844),
            .I(N__4836));
    LocalMux I__683 (
            .O(N__4841),
            .I(N__4836));
    Span4Mux_h I__682 (
            .O(N__4836),
            .I(N__4831));
    InMux I__681 (
            .O(N__4835),
            .I(N__4826));
    InMux I__680 (
            .O(N__4834),
            .I(N__4826));
    Span4Mux_v I__679 (
            .O(N__4831),
            .I(N__4823));
    LocalMux I__678 (
            .O(N__4826),
            .I(N__4820));
    Span4Mux_v I__677 (
            .O(N__4823),
            .I(N__4817));
    Sp12to4 I__676 (
            .O(N__4820),
            .I(N__4814));
    Sp12to4 I__675 (
            .O(N__4817),
            .I(N__4809));
    Span12Mux_v I__674 (
            .O(N__4814),
            .I(N__4809));
    Odrv12 I__673 (
            .O(N__4809),
            .I(A_c_1));
    InMux I__672 (
            .O(N__4806),
            .I(N__4803));
    LocalMux I__671 (
            .O(N__4803),
            .I(\U712_BYTE_ENABLE.un1_CLMBEn_i_0Z0Z_0 ));
    InMux I__670 (
            .O(N__4800),
            .I(N__4797));
    LocalMux I__669 (
            .O(N__4797),
            .I(N__4794));
    Span4Mux_v I__668 (
            .O(N__4794),
            .I(N__4791));
    Span4Mux_h I__667 (
            .O(N__4791),
            .I(N__4788));
    Span4Mux_v I__666 (
            .O(N__4788),
            .I(N__4785));
    Odrv4 I__665 (
            .O(N__4785),
            .I(TACK_EN_i_ess));
    InMux I__664 (
            .O(N__4782),
            .I(N__4777));
    InMux I__663 (
            .O(N__4781),
            .I(N__4774));
    InMux I__662 (
            .O(N__4780),
            .I(N__4771));
    LocalMux I__661 (
            .O(N__4777),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__660 (
            .O(N__4774),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__659 (
            .O(N__4771),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CascadeMux I__658 (
            .O(N__4764),
            .I(N__4760));
    CascadeMux I__657 (
            .O(N__4763),
            .I(N__4757));
    InMux I__656 (
            .O(N__4760),
            .I(N__4754));
    InMux I__655 (
            .O(N__4757),
            .I(N__4751));
    LocalMux I__654 (
            .O(N__4754),
            .I(N__4748));
    LocalMux I__653 (
            .O(N__4751),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    Odrv4 I__652 (
            .O(N__4748),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    InMux I__651 (
            .O(N__4743),
            .I(N__4738));
    InMux I__650 (
            .O(N__4742),
            .I(N__4735));
    InMux I__649 (
            .O(N__4741),
            .I(N__4732));
    LocalMux I__648 (
            .O(N__4738),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__647 (
            .O(N__4735),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__646 (
            .O(N__4732),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__645 (
            .O(N__4725),
            .I(\U712_CYCLE_TERM.N_233_i_0_en_cascade_ ));
    CEMux I__644 (
            .O(N__4722),
            .I(N__4719));
    LocalMux I__643 (
            .O(N__4719),
            .I(\U712_CYCLE_TERM.N_233_i_0_en_0 ));
    InMux I__642 (
            .O(N__4716),
            .I(N__4713));
    LocalMux I__641 (
            .O(N__4713),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ));
    InMux I__640 (
            .O(N__4710),
            .I(N__4707));
    LocalMux I__639 (
            .O(N__4707),
            .I(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ));
    CascadeMux I__638 (
            .O(N__4704),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_i_2_cascade_ ));
    InMux I__637 (
            .O(N__4701),
            .I(N__4697));
    InMux I__636 (
            .O(N__4700),
            .I(N__4694));
    LocalMux I__635 (
            .O(N__4697),
            .I(N__4691));
    LocalMux I__634 (
            .O(N__4694),
            .I(CPU_TACKm));
    Odrv4 I__633 (
            .O(N__4691),
            .I(CPU_TACKm));
    InMux I__632 (
            .O(N__4686),
            .I(N__4682));
    InMux I__631 (
            .O(N__4685),
            .I(N__4679));
    LocalMux I__630 (
            .O(N__4682),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__629 (
            .O(N__4679),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__628 (
            .O(N__4674),
            .I(N__4670));
    InMux I__627 (
            .O(N__4673),
            .I(N__4667));
    LocalMux I__626 (
            .O(N__4670),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__625 (
            .O(N__4667),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__624 (
            .O(N__4662),
            .I(N__4658));
    InMux I__623 (
            .O(N__4661),
            .I(N__4655));
    InMux I__622 (
            .O(N__4658),
            .I(N__4652));
    LocalMux I__621 (
            .O(N__4655),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__620 (
            .O(N__4652),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__619 (
            .O(N__4647),
            .I(N__4643));
    InMux I__618 (
            .O(N__4646),
            .I(N__4640));
    LocalMux I__617 (
            .O(N__4643),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__616 (
            .O(N__4640),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__615 (
            .O(N__4635),
            .I(N__4632));
    LocalMux I__614 (
            .O(N__4632),
            .I(\U712_CHIP_RAM.N_218 ));
    CascadeMux I__613 (
            .O(N__4629),
            .I(\U712_CHIP_RAM.N_208_cascade_ ));
    CascadeMux I__612 (
            .O(N__4626),
            .I(\U712_CHIP_RAM.N_245_cascade_ ));
    InMux I__611 (
            .O(N__4623),
            .I(N__4620));
    LocalMux I__610 (
            .O(N__4620),
            .I(\U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a3_0_2 ));
    InMux I__609 (
            .O(N__4617),
            .I(N__4614));
    LocalMux I__608 (
            .O(N__4614),
            .I(N__4611));
    Span4Mux_v I__607 (
            .O(N__4611),
            .I(N__4608));
    Sp12to4 I__606 (
            .O(N__4608),
            .I(N__4605));
    Odrv12 I__605 (
            .O(N__4605),
            .I(A_c_4));
    InMux I__604 (
            .O(N__4602),
            .I(N__4599));
    LocalMux I__603 (
            .O(N__4599),
            .I(N__4596));
    Sp12to4 I__602 (
            .O(N__4596),
            .I(N__4593));
    Span12Mux_v I__601 (
            .O(N__4593),
            .I(N__4590));
    Odrv12 I__600 (
            .O(N__4590),
            .I(A_c_11));
    CascadeMux I__599 (
            .O(N__4587),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ));
    InMux I__598 (
            .O(N__4584),
            .I(N__4581));
    LocalMux I__597 (
            .O(N__4581),
            .I(\U712_BYTE_ENABLE.N_327 ));
    InMux I__596 (
            .O(N__4578),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__595 (
            .O(N__4575),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__594 (
            .O(N__4572),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__593 (
            .O(N__4569),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__592 (
            .O(N__4566),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    CascadeMux I__591 (
            .O(N__4563),
            .I(\U712_CHIP_RAM.N_282_cascade_ ));
    CascadeMux I__590 (
            .O(N__4560),
            .I(\U712_CHIP_RAM.N_265_cascade_ ));
    InMux I__589 (
            .O(N__4557),
            .I(N__4553));
    InMux I__588 (
            .O(N__4556),
            .I(N__4550));
    LocalMux I__587 (
            .O(N__4553),
            .I(REG_TACK));
    LocalMux I__586 (
            .O(N__4550),
            .I(REG_TACK));
    CascadeMux I__585 (
            .O(N__4545),
            .I(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ));
    InMux I__584 (
            .O(N__4542),
            .I(N__4539));
    LocalMux I__583 (
            .O(N__4539),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_2 ));
    IoInMux I__582 (
            .O(N__4536),
            .I(N__4533));
    LocalMux I__581 (
            .O(N__4533),
            .I(N__4530));
    Span4Mux_s1_h I__580 (
            .O(N__4530),
            .I(N__4527));
    Sp12to4 I__579 (
            .O(N__4527),
            .I(N__4524));
    Span12Mux_v I__578 (
            .O(N__4524),
            .I(N__4520));
    InMux I__577 (
            .O(N__4523),
            .I(N__4517));
    Odrv12 I__576 (
            .O(N__4520),
            .I(TACK_OUTn));
    LocalMux I__575 (
            .O(N__4517),
            .I(TACK_OUTn));
    InMux I__574 (
            .O(N__4512),
            .I(N__4508));
    InMux I__573 (
            .O(N__4511),
            .I(N__4505));
    LocalMux I__572 (
            .O(N__4508),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    LocalMux I__571 (
            .O(N__4505),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__570 (
            .O(N__4500),
            .I(N__4496));
    InMux I__569 (
            .O(N__4499),
            .I(N__4493));
    LocalMux I__568 (
            .O(N__4496),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__567 (
            .O(N__4493),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__566 (
            .O(N__4488),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__565 (
            .O(N__4485),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    CascadeMux I__564 (
            .O(N__4482),
            .I(N__4479));
    InMux I__563 (
            .O(N__4479),
            .I(N__4474));
    InMux I__562 (
            .O(N__4478),
            .I(N__4469));
    InMux I__561 (
            .O(N__4477),
            .I(N__4469));
    LocalMux I__560 (
            .O(N__4474),
            .I(N__4460));
    LocalMux I__559 (
            .O(N__4469),
            .I(N__4460));
    InMux I__558 (
            .O(N__4468),
            .I(N__4451));
    InMux I__557 (
            .O(N__4467),
            .I(N__4451));
    InMux I__556 (
            .O(N__4466),
            .I(N__4451));
    InMux I__555 (
            .O(N__4465),
            .I(N__4451));
    Odrv4 I__554 (
            .O(N__4460),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__553 (
            .O(N__4451),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    InMux I__552 (
            .O(N__4446),
            .I(N__4438));
    InMux I__551 (
            .O(N__4445),
            .I(N__4438));
    InMux I__550 (
            .O(N__4444),
            .I(N__4435));
    InMux I__549 (
            .O(N__4443),
            .I(N__4432));
    LocalMux I__548 (
            .O(N__4438),
            .I(N__4429));
    LocalMux I__547 (
            .O(N__4435),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__546 (
            .O(N__4432),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv4 I__545 (
            .O(N__4429),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    InMux I__544 (
            .O(N__4422),
            .I(N__4419));
    LocalMux I__543 (
            .O(N__4419),
            .I(\U712_REG_SM.STATE_COUNT_srsts_i_i_0_0_3 ));
    InMux I__542 (
            .O(N__4416),
            .I(N__4410));
    InMux I__541 (
            .O(N__4415),
            .I(N__4406));
    InMux I__540 (
            .O(N__4414),
            .I(N__4403));
    InMux I__539 (
            .O(N__4413),
            .I(N__4400));
    LocalMux I__538 (
            .O(N__4410),
            .I(N__4397));
    InMux I__537 (
            .O(N__4409),
            .I(N__4394));
    LocalMux I__536 (
            .O(N__4406),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__535 (
            .O(N__4403),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__534 (
            .O(N__4400),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    Odrv4 I__533 (
            .O(N__4397),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__532 (
            .O(N__4394),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    CascadeMux I__531 (
            .O(N__4383),
            .I(N__4377));
    CascadeMux I__530 (
            .O(N__4382),
            .I(N__4371));
    InMux I__529 (
            .O(N__4381),
            .I(N__4367));
    InMux I__528 (
            .O(N__4380),
            .I(N__4364));
    InMux I__527 (
            .O(N__4377),
            .I(N__4361));
    InMux I__526 (
            .O(N__4376),
            .I(N__4356));
    InMux I__525 (
            .O(N__4375),
            .I(N__4356));
    InMux I__524 (
            .O(N__4374),
            .I(N__4349));
    InMux I__523 (
            .O(N__4371),
            .I(N__4349));
    InMux I__522 (
            .O(N__4370),
            .I(N__4349));
    LocalMux I__521 (
            .O(N__4367),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__520 (
            .O(N__4364),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__519 (
            .O(N__4361),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__518 (
            .O(N__4356),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__517 (
            .O(N__4349),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    IoInMux I__516 (
            .O(N__4338),
            .I(N__4335));
    LocalMux I__515 (
            .O(N__4335),
            .I(N__4332));
    IoSpan4Mux I__514 (
            .O(N__4332),
            .I(N__4329));
    Sp12to4 I__513 (
            .O(N__4329),
            .I(N__4326));
    Span12Mux_s7_v I__512 (
            .O(N__4326),
            .I(N__4323));
    Odrv12 I__511 (
            .O(N__4323),
            .I(N_40_i));
    InMux I__510 (
            .O(N__4320),
            .I(N__4317));
    LocalMux I__509 (
            .O(N__4317),
            .I(\U712_REG_SM.N_261 ));
    CascadeMux I__508 (
            .O(N__4314),
            .I(N__4307));
    InMux I__507 (
            .O(N__4313),
            .I(N__4304));
    InMux I__506 (
            .O(N__4312),
            .I(N__4301));
    InMux I__505 (
            .O(N__4311),
            .I(N__4298));
    InMux I__504 (
            .O(N__4310),
            .I(N__4293));
    InMux I__503 (
            .O(N__4307),
            .I(N__4293));
    LocalMux I__502 (
            .O(N__4304),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__501 (
            .O(N__4301),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__500 (
            .O(N__4298),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__499 (
            .O(N__4293),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    CascadeMux I__498 (
            .O(N__4284),
            .I(N__4280));
    InMux I__497 (
            .O(N__4283),
            .I(N__4275));
    InMux I__496 (
            .O(N__4280),
            .I(N__4272));
    InMux I__495 (
            .O(N__4279),
            .I(N__4267));
    InMux I__494 (
            .O(N__4278),
            .I(N__4267));
    LocalMux I__493 (
            .O(N__4275),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__492 (
            .O(N__4272),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__491 (
            .O(N__4267),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    InMux I__490 (
            .O(N__4260),
            .I(N__4257));
    LocalMux I__489 (
            .O(N__4257),
            .I(N__4249));
    InMux I__488 (
            .O(N__4256),
            .I(N__4246));
    InMux I__487 (
            .O(N__4255),
            .I(N__4243));
    InMux I__486 (
            .O(N__4254),
            .I(N__4240));
    InMux I__485 (
            .O(N__4253),
            .I(N__4237));
    InMux I__484 (
            .O(N__4252),
            .I(N__4234));
    Odrv4 I__483 (
            .O(N__4249),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__482 (
            .O(N__4246),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__481 (
            .O(N__4243),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__480 (
            .O(N__4240),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__479 (
            .O(N__4237),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__478 (
            .O(N__4234),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    IoInMux I__477 (
            .O(N__4221),
            .I(N__4218));
    LocalMux I__476 (
            .O(N__4218),
            .I(N__4215));
    Span12Mux_s10_h I__475 (
            .O(N__4215),
            .I(N__4212));
    Span12Mux_h I__474 (
            .O(N__4212),
            .I(N__4209));
    Span12Mux_v I__473 (
            .O(N__4209),
            .I(N__4206));
    Odrv12 I__472 (
            .O(N__4206),
            .I(N_41_i));
    InMux I__471 (
            .O(N__4203),
            .I(N__4200));
    LocalMux I__470 (
            .O(N__4200),
            .I(\U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_0 ));
    CascadeMux I__469 (
            .O(N__4197),
            .I(N__4194));
    InMux I__468 (
            .O(N__4194),
            .I(N__4191));
    LocalMux I__467 (
            .O(N__4191),
            .I(\U712_REG_SM.DS_EN_RNOZ0Z_0 ));
    InMux I__466 (
            .O(N__4188),
            .I(N__4185));
    LocalMux I__465 (
            .O(N__4185),
            .I(N__4182));
    Odrv4 I__464 (
            .O(N__4182),
            .I(\U712_REG_SM.N_314 ));
    InMux I__463 (
            .O(N__4179),
            .I(N__4173));
    InMux I__462 (
            .O(N__4178),
            .I(N__4170));
    InMux I__461 (
            .O(N__4177),
            .I(N__4167));
    InMux I__460 (
            .O(N__4176),
            .I(N__4164));
    LocalMux I__459 (
            .O(N__4173),
            .I(\U712_REG_SM.N_225 ));
    LocalMux I__458 (
            .O(N__4170),
            .I(\U712_REG_SM.N_225 ));
    LocalMux I__457 (
            .O(N__4167),
            .I(\U712_REG_SM.N_225 ));
    LocalMux I__456 (
            .O(N__4164),
            .I(\U712_REG_SM.N_225 ));
    CascadeMux I__455 (
            .O(N__4155),
            .I(\U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_1_1_3_cascade_ ));
    CascadeMux I__454 (
            .O(N__4152),
            .I(N__4149));
    InMux I__453 (
            .O(N__4149),
            .I(N__4146));
    LocalMux I__452 (
            .O(N__4146),
            .I(\U712_REG_SM.N_259 ));
    CascadeMux I__451 (
            .O(N__4143),
            .I(\U712_REG_SM.N_259_cascade_ ));
    InMux I__450 (
            .O(N__4140),
            .I(N__4137));
    LocalMux I__449 (
            .O(N__4137),
            .I(N__4133));
    InMux I__448 (
            .O(N__4136),
            .I(N__4130));
    Odrv4 I__447 (
            .O(N__4133),
            .I(\U712_REG_SM.N_236 ));
    LocalMux I__446 (
            .O(N__4130),
            .I(\U712_REG_SM.N_236 ));
    InMux I__445 (
            .O(N__4125),
            .I(N__4115));
    InMux I__444 (
            .O(N__4124),
            .I(N__4115));
    InMux I__443 (
            .O(N__4123),
            .I(N__4110));
    InMux I__442 (
            .O(N__4122),
            .I(N__4110));
    InMux I__441 (
            .O(N__4121),
            .I(N__4105));
    InMux I__440 (
            .O(N__4120),
            .I(N__4105));
    LocalMux I__439 (
            .O(N__4115),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__438 (
            .O(N__4110),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__437 (
            .O(N__4105),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    IoInMux I__436 (
            .O(N__4098),
            .I(N__4095));
    LocalMux I__435 (
            .O(N__4095),
            .I(N__4092));
    Span12Mux_s7_v I__434 (
            .O(N__4092),
            .I(N__4088));
    InMux I__433 (
            .O(N__4091),
            .I(N__4084));
    Span12Mux_v I__432 (
            .O(N__4088),
            .I(N__4081));
    InMux I__431 (
            .O(N__4087),
            .I(N__4078));
    LocalMux I__430 (
            .O(N__4084),
            .I(N__4075));
    Odrv12 I__429 (
            .O(N__4081),
            .I(REGENn_c));
    LocalMux I__428 (
            .O(N__4078),
            .I(REGENn_c));
    Odrv12 I__427 (
            .O(N__4075),
            .I(REGENn_c));
    InMux I__426 (
            .O(N__4068),
            .I(N__4065));
    LocalMux I__425 (
            .O(N__4065),
            .I(\U712_REG_SM.N_307 ));
    CascadeMux I__424 (
            .O(N__4062),
            .I(N__4059));
    InMux I__423 (
            .O(N__4059),
            .I(N__4055));
    InMux I__422 (
            .O(N__4058),
            .I(N__4052));
    LocalMux I__421 (
            .O(N__4055),
            .I(\U712_REG_SM.N_219 ));
    LocalMux I__420 (
            .O(N__4052),
            .I(\U712_REG_SM.N_219 ));
    CascadeMux I__419 (
            .O(N__4047),
            .I(N__4044));
    InMux I__418 (
            .O(N__4044),
            .I(N__4041));
    LocalMux I__417 (
            .O(N__4041),
            .I(\U712_REG_SM.REG_TACK_RNOZ0Z_0 ));
    CascadeMux I__416 (
            .O(N__4038),
            .I(N__4034));
    InMux I__415 (
            .O(N__4037),
            .I(N__4031));
    InMux I__414 (
            .O(N__4034),
            .I(N__4028));
    LocalMux I__413 (
            .O(N__4031),
            .I(\U712_REG_SM.N_235 ));
    LocalMux I__412 (
            .O(N__4028),
            .I(\U712_REG_SM.N_235 ));
    CascadeMux I__411 (
            .O(N__4023),
            .I(\U712_CHIP_RAM.un5_DMA_CYCLE_START_0_cascade_ ));
    CascadeMux I__410 (
            .O(N__4020),
            .I(\U712_REG_SM.N_219_cascade_ ));
    InMux I__409 (
            .O(N__4017),
            .I(N__4014));
    LocalMux I__408 (
            .O(N__4014),
            .I(\U712_REG_SM.N_304 ));
    CascadeMux I__407 (
            .O(N__4011),
            .I(\U712_REG_SM.N_304_cascade_ ));
    CascadeMux I__406 (
            .O(N__4008),
            .I(N__4005));
    InMux I__405 (
            .O(N__4005),
            .I(N__4002));
    LocalMux I__404 (
            .O(N__4002),
            .I(N__3999));
    Odrv4 I__403 (
            .O(N__3999),
            .I(\U712_REG_SM.STATE_COUNT_srsts_i_0_i_0_1 ));
    InMux I__402 (
            .O(N__3996),
            .I(N__3993));
    LocalMux I__401 (
            .O(N__3993),
            .I(N__3989));
    IoInMux I__400 (
            .O(N__3992),
            .I(N__3986));
    Span4Mux_v I__399 (
            .O(N__3989),
            .I(N__3983));
    LocalMux I__398 (
            .O(N__3986),
            .I(N__3980));
    Sp12to4 I__397 (
            .O(N__3983),
            .I(N__3977));
    IoSpan4Mux I__396 (
            .O(N__3980),
            .I(N__3974));
    Span12Mux_h I__395 (
            .O(N__3977),
            .I(N__3971));
    IoSpan4Mux I__394 (
            .O(N__3974),
            .I(N__3968));
    Span12Mux_v I__393 (
            .O(N__3971),
            .I(N__3965));
    IoSpan4Mux I__392 (
            .O(N__3968),
            .I(N__3962));
    Odrv12 I__391 (
            .O(N__3965),
            .I(C3_c));
    Odrv4 I__390 (
            .O(N__3962),
            .I(C3_c));
    InMux I__389 (
            .O(N__3957),
            .I(N__3954));
    LocalMux I__388 (
            .O(N__3954),
            .I(N__3950));
    IoInMux I__387 (
            .O(N__3953),
            .I(N__3947));
    Span4Mux_v I__386 (
            .O(N__3950),
            .I(N__3944));
    LocalMux I__385 (
            .O(N__3947),
            .I(N__3941));
    Sp12to4 I__384 (
            .O(N__3944),
            .I(N__3938));
    Span4Mux_s3_h I__383 (
            .O(N__3941),
            .I(N__3935));
    Span12Mux_h I__382 (
            .O(N__3938),
            .I(N__3930));
    Sp12to4 I__381 (
            .O(N__3935),
            .I(N__3930));
    Span12Mux_v I__380 (
            .O(N__3930),
            .I(N__3927));
    Odrv12 I__379 (
            .O(N__3927),
            .I(C1_c));
    CascadeMux I__378 (
            .O(N__3924),
            .I(N__3921));
    InMux I__377 (
            .O(N__3921),
            .I(N__3918));
    LocalMux I__376 (
            .O(N__3918),
            .I(N__3915));
    Span4Mux_h I__375 (
            .O(N__3915),
            .I(N__3912));
    Span4Mux_v I__374 (
            .O(N__3912),
            .I(N__3909));
    Span4Mux_v I__373 (
            .O(N__3909),
            .I(N__3906));
    Span4Mux_v I__372 (
            .O(N__3906),
            .I(N__3903));
    Odrv4 I__371 (
            .O(N__3903),
            .I(REGSPACEn_c));
    InMux I__370 (
            .O(N__3900),
            .I(N__3896));
    InMux I__369 (
            .O(N__3899),
            .I(N__3893));
    LocalMux I__368 (
            .O(N__3896),
            .I(N__3890));
    LocalMux I__367 (
            .O(N__3893),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    Odrv4 I__366 (
            .O(N__3890),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    IoInMux I__365 (
            .O(N__3885),
            .I(N__3882));
    LocalMux I__364 (
            .O(N__3882),
            .I(N__3879));
    IoSpan4Mux I__363 (
            .O(N__3879),
            .I(N__3876));
    IoSpan4Mux I__362 (
            .O(N__3876),
            .I(N__3873));
    Span4Mux_s3_h I__361 (
            .O(N__3873),
            .I(N__3870));
    Odrv4 I__360 (
            .O(N__3870),
            .I(N_991_i));
    IoInMux I__359 (
            .O(N__3867),
            .I(N__3864));
    LocalMux I__358 (
            .O(N__3864),
            .I(N__3861));
    IoSpan4Mux I__357 (
            .O(N__3861),
            .I(N__3858));
    Span4Mux_s2_v I__356 (
            .O(N__3858),
            .I(N__3855));
    Span4Mux_v I__355 (
            .O(N__3855),
            .I(N__3852));
    Odrv4 I__354 (
            .O(N__3852),
            .I(CLK80_PLL_i_i));
    IoInMux I__353 (
            .O(N__3849),
            .I(N__3846));
    LocalMux I__352 (
            .O(N__3846),
            .I(N__3843));
    Span4Mux_s3_v I__351 (
            .O(N__3843),
            .I(N__3840));
    Span4Mux_h I__350 (
            .O(N__3840),
            .I(N__3837));
    Span4Mux_h I__349 (
            .O(N__3837),
            .I(N__3834));
    Sp12to4 I__348 (
            .O(N__3834),
            .I(N__3831));
    Span12Mux_s8_v I__347 (
            .O(N__3831),
            .I(N__3828));
    Span12Mux_h I__346 (
            .O(N__3828),
            .I(N__3824));
    InMux I__345 (
            .O(N__3827),
            .I(N__3821));
    Odrv12 I__344 (
            .O(N__3824),
            .I(ASn_c));
    LocalMux I__343 (
            .O(N__3821),
            .I(ASn_c));
    CascadeMux I__342 (
            .O(N__3816),
            .I(\U712_REG_SM.N_238_cascade_ ));
    InMux I__341 (
            .O(N__3813),
            .I(N__3809));
    InMux I__340 (
            .O(N__3812),
            .I(N__3806));
    LocalMux I__339 (
            .O(N__3809),
            .I(\U712_REG_SM.N_238 ));
    LocalMux I__338 (
            .O(N__3806),
            .I(\U712_REG_SM.N_238 ));
    InMux I__337 (
            .O(N__3801),
            .I(N__3797));
    InMux I__336 (
            .O(N__3800),
            .I(N__3794));
    LocalMux I__335 (
            .O(N__3797),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__334 (
            .O(N__3794),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    CascadeMux I__333 (
            .O(N__3789),
            .I(N__3785));
    InMux I__332 (
            .O(N__3788),
            .I(N__3780));
    InMux I__331 (
            .O(N__3785),
            .I(N__3780));
    LocalMux I__330 (
            .O(N__3780),
            .I(\U712_REG_SM.ASn_0_sqmuxa_1 ));
    IoInMux I__329 (
            .O(N__3777),
            .I(N__3774));
    LocalMux I__328 (
            .O(N__3774),
            .I(N__3771));
    IoSpan4Mux I__327 (
            .O(N__3771),
            .I(N__3768));
    Span4Mux_s2_v I__326 (
            .O(N__3768),
            .I(N__3765));
    Sp12to4 I__325 (
            .O(N__3765),
            .I(N__3762));
    Span12Mux_v I__324 (
            .O(N__3762),
            .I(N__3759));
    Odrv12 I__323 (
            .O(N__3759),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__8863));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__8865));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__8866));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__8867));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .I(N__8868));
    INV \INVU712_CHIP_RAM.DMA_A20C  (
            .O(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .I(N__8864));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__8568),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__3953),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__3992),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam TACKn_obuft_RNO_LC_1_14_3.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_1_14_3.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_1_14_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_obuft_RNO_LC_1_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4800),
            .lcout(N_991_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_5_1_4.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_5_1_4.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_5_1_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_5_1_4 (
            .in0(N__9105),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_LC_5_7_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_5_7_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_5_7_0 .LUT_INIT=16'b1111101111110000;
    LogicCell40 \U712_REG_SM.REGENn_LC_5_7_0  (
            .in0(N__3812),
            .in1(N__3801),
            .in2(N__3789),
            .in3(N__4087),
            .lcout(REGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9092),
            .ce(),
            .sr(N__9997));
    defparam \U712_REG_SM.ASn_LC_5_7_3 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_LC_5_7_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_LC_5_7_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U712_REG_SM.ASn_LC_5_7_3  (
            .in0(N__3827),
            .in1(N__3788),
            .in2(_gnd_net_),
            .in3(N__4140),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9092),
            .ce(),
            .sr(N__9997));
    defparam \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_5_8_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_5_8_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(N__4176),
            .in2(_gnd_net_),
            .in3(N__3900),
            .lcout(\U712_REG_SM.N_238 ),
            .ltout(\U712_REG_SM.N_238_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_5_8_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_5_8_1 .LUT_INIT=16'b1101010111110111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_5_8_1  (
            .in0(N__8709),
            .in1(N__3800),
            .in2(N__3816),
            .in3(N__4254),
            .lcout(\U712_REG_SM.STATE_COUNT_srsts_i_0_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_5_8_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_5_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_5_8_2 .LUT_INIT=16'b0001001100010001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_5_8_2  (
            .in0(N__8708),
            .in1(N__4017),
            .in2(N__4038),
            .in3(N__3813),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9096),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_5_8_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_5_8_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_5_8_5  (
            .in0(_gnd_net_),
            .in1(N__4413),
            .in2(_gnd_net_),
            .in3(N__4058),
            .lcout(\U712_REG_SM.ASn_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_5_9_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_5_9_1 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_5_9_1  (
            .in0(N__4278),
            .in1(N__4370),
            .in2(N__4314),
            .in3(N__4120),
            .lcout(\U712_REG_SM.N_225 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_5_9_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_5_9_3 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_5_9_3  (
            .in0(N__4124),
            .in1(N__4253),
            .in2(N__4383),
            .in3(N__8880),
            .lcout(\U712_REG_SM.N_236 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_5_9_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_5_9_4 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_5_9_4  (
            .in0(N__4121),
            .in1(N__4279),
            .in2(N__4382),
            .in3(N__4310),
            .lcout(\U712_REG_SM.N_219 ),
            .ltout(\U712_REG_SM.N_219_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIEMV42_4_LC_5_9_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIEMV42_4_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIEMV42_4_LC_5_9_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIEMV42_4_LC_5_9_5  (
            .in0(_gnd_net_),
            .in1(N__8707),
            .in2(N__4020),
            .in3(N__4414),
            .lcout(\U712_REG_SM.N_304 ),
            .ltout(\U712_REG_SM.N_304_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_5_9_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_5_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_5_9_6 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_5_9_6  (
            .in0(N__8706),
            .in1(N__4444),
            .in2(N__4011),
            .in3(N__4178),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9098),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_5_9_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_5_9_7 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_5_9_7  (
            .in0(N__4125),
            .in1(N__4374),
            .in2(N__4008),
            .in3(N__8881),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9098),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_0_LC_5_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_5_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_5_10_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_5_10_0  (
            .in0(N__3996),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9099),
            .ce(),
            .sr(N__9990));
    defparam \U712_REG_SM.C1_SYNC_1_LC_5_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_5_10_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_5_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4313),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9099),
            .ce(),
            .sr(N__9990));
    defparam \U712_REG_SM.C1_SYNC_0_LC_5_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_5_10_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_5_10_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_5_10_3  (
            .in0(N__3957),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9099),
            .ce(),
            .sr(N__9990));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_5_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_5_10_4 .LUT_INIT=16'b0000010111001101;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_5_10_4  (
            .in0(N__5879),
            .in1(N__3899),
            .in2(N__3924),
            .in3(N__5299),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9099),
            .ce(),
            .sr(N__9990));
    defparam \U712_REG_SM.C3_SYNC_1_LC_5_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_5_10_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_5_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4381),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9099),
            .ce(),
            .sr(N__9990));
    defparam DBR_SYNC_0_LC_5_11_6.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_5_11_6.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_5_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_5_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8923),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9101),
            .ce(),
            .sr(N__9982));
    defparam \U712_REG_SM.REG_CYCLE_LC_5_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_5_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_5_13_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_5_13_2  (
            .in0(N__8705),
            .in1(N__8911),
            .in2(_gnd_net_),
            .in3(N__4091),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10136),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_6_7_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_6_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6429),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9085),
            .ce(),
            .sr(N__9996));
    defparam \U712_REG_SM.REG_TACK_LC_6_7_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_6_7_5 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_6_7_5  (
            .in0(N__4037),
            .in1(N__4068),
            .in2(N__4047),
            .in3(N__4557),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9085),
            .ce(),
            .sr(N__9996));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_6_8_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_6_8_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_6_8_0  (
            .in0(N__4478),
            .in1(N__4256),
            .in2(_gnd_net_),
            .in3(N__4177),
            .lcout(\U712_REG_SM.N_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_6_8_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_6_8_4 .LUT_INIT=16'b1010111000000100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_6_8_4  (
            .in0(N__6654),
            .in1(N__4409),
            .in2(N__4062),
            .in3(N__4446),
            .lcout(\U712_REG_SM.REG_TACK_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_6_8_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_6_8_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_6_8_5  (
            .in0(N__4445),
            .in1(N__4252),
            .in2(_gnd_net_),
            .in3(N__4477),
            .lcout(\U712_REG_SM.N_235 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_6_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_6_9_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__4499),
            .in2(_gnd_net_),
            .in3(N__4511),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un5_DMA_CYCLE_START_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_6_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_6_9_2 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_6_9_2  (
            .in0(N__5737),
            .in1(N__4542),
            .in2(N__4023),
            .in3(N__6755),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9093),
            .ce(),
            .sr(N__9987));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_6_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_6_9_3 .LUT_INIT=16'b0010101000100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_6_9_3  (
            .in0(N__8702),
            .in1(N__6201),
            .in2(N__5757),
            .in3(N__5811),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_a4_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_6_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_6_9_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_6_9_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_6_9_5  (
            .in0(N__4977),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5382),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9093),
            .ce(),
            .sr(N__9987));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_6_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_6_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_6_9_6 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_6_9_6  (
            .in0(N__6202),
            .in1(N__6880),
            .in2(_gnd_net_),
            .in3(N__5481),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9093),
            .ce(),
            .sr(N__9987));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOO5O1_LC_6_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOO5O1_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOO5O1_LC_6_9_7 .LUT_INIT=16'b0000001001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOO5O1_LC_6_9_7  (
            .in0(N__7025),
            .in1(N__6200),
            .in2(N__6911),
            .in3(N__7177),
            .lcout(\U712_CHIP_RAM.N_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_6_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_6_10_0 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_6_10_0  (
            .in0(N__4422),
            .in1(N__4179),
            .in2(N__4152),
            .in3(N__4468),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9097),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI07K21_1_LC_6_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI07K21_1_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI07K21_1_LC_6_10_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI07K21_1_LC_6_10_1  (
            .in0(N__4376),
            .in1(N__4123),
            .in2(N__6450),
            .in3(N__6461),
            .lcout(),
            .ltout(\U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_1_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI35EO1_1_LC_6_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI35EO1_1_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI35EO1_1_LC_6_10_2 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI35EO1_1_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(N__4283),
            .in2(N__4155),
            .in3(N__4311),
            .lcout(\U712_REG_SM.N_259 ),
            .ltout(\U712_REG_SM.N_259_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_6_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_6_10_3 .LUT_INIT=16'b1000000011000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_6_10_3  (
            .in0(N__4467),
            .in1(N__8700),
            .in2(N__4143),
            .in3(N__4136),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9097),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_3_LC_6_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_3_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_3_LC_6_10_4 .LUT_INIT=16'b0111011111101110;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_3_LC_6_10_4  (
            .in0(N__4122),
            .in1(N__4465),
            .in2(_gnd_net_),
            .in3(N__4375),
            .lcout(\U712_REG_SM.N_261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_6_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_6_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_6_10_5  (
            .in0(N__6650),
            .in1(N__6702),
            .in2(_gnd_net_),
            .in3(N__5733),
            .lcout(\U712_CHIP_RAM.N_257 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_6_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_6_10_6 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_1_LC_6_10_6  (
            .in0(N__4255),
            .in1(N__4415),
            .in2(N__4482),
            .in3(N__8882),
            .lcout(\U712_REG_SM.N_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_6_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_6_10_7 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_6_10_7  (
            .in0(N__4466),
            .in1(N__8701),
            .in2(_gnd_net_),
            .in3(N__4443),
            .lcout(\U712_REG_SM.STATE_COUNT_srsts_i_i_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_6_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_6_11_2 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_6_11_2  (
            .in0(N__6649),
            .in1(N__4416),
            .in2(_gnd_net_),
            .in3(N__4380),
            .lcout(\U712_REG_SM.DS_EN_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_40_i_LC_6_11_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_40_i_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_40_i_LC_6_11_3 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \U712_BYTE_ENABLE.N_40_i_LC_6_11_3  (
            .in0(N__4847),
            .in1(N__4872),
            .in2(N__5412),
            .in3(N__4584),
            .lcout(N_40_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_6_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_6_11_4 .LUT_INIT=16'b1010101010111111;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_2_LC_6_11_4  (
            .in0(N__4320),
            .in1(N__4312),
            .in2(N__4284),
            .in3(N__4260),
            .lcout(\U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_6_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_6_11_5 .LUT_INIT=16'b0000100000001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_6_11_5  (
            .in0(N__5756),
            .in1(N__6239),
            .in2(N__6141),
            .in3(N__5810),
            .lcout(\U712_CHIP_RAM.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_41_i_LC_6_12_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_41_i_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_41_i_LC_6_12_0 .LUT_INIT=16'b0011001000110011;
    LogicCell40 \U712_BYTE_ENABLE.N_41_i_LC_6_12_0  (
            .in0(N__5465),
            .in1(N__4806),
            .in2(N__4975),
            .in3(N__6764),
            .lcout(N_41_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_LC_6_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_6_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_6_12_7 .LUT_INIT=16'b1100110010001101;
    LogicCell40 \U712_REG_SM.DS_EN_LC_6_12_7  (
            .in0(N__4203),
            .in1(N__8474),
            .in2(N__4197),
            .in3(N__4188),
            .lcout(DS_ENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9100),
            .ce(),
            .sr(N__9959));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_7_7_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_7_7_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_7_7_1  (
            .in0(N__4701),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4556),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_7_7_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_7_7_2 .LUT_INIT=16'b1100111110001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_7_7_2  (
            .in0(N__8817),
            .in1(N__6391),
            .in2(N__4545),
            .in3(N__4742),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9082),
            .ce(),
            .sr(N__9994));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_7_7_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_7_7_5 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_7_7_5 .LUT_INIT=16'b0101010001010000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_7_7_5  (
            .in0(N__6390),
            .in1(N__4716),
            .in2(N__4763),
            .in3(N__4781),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9082),
            .ce(),
            .sr(N__9994));
    defparam \U712_CHIP_RAM.CAS_SYNC_2_LC_7_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_2_LC_7_8_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_2_LC_7_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_2_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4500),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9086),
            .ce(),
            .sr(N__9988));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_7_8_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_7_8_5 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_7_8_5 .LUT_INIT=16'b1111111111000100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_7_8_5  (
            .in0(N__6395),
            .in1(N__4523),
            .in2(N__8826),
            .in3(N__6425),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9086),
            .ce(),
            .sr(N__9988));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_7_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_7_8_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_7_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4512),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9086),
            .ce(),
            .sr(N__9988));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_9_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_9_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__6125),
            .in2(_gnd_net_),
            .in3(N__6238),
            .lcout(\U712_CHIP_RAM.N_243 ),
            .ltout(),
            .carryin(bfn_7_9_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_9_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_9_1  (
            .in0(N__5084),
            .in1(N__6920),
            .in2(_gnd_net_),
            .in3(N__4488),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__9089),
            .ce(N__5052),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_9_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(N__7038),
            .in2(_gnd_net_),
            .in3(N__4485),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_9_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_9_3  (
            .in0(N__5085),
            .in1(N__7216),
            .in2(_gnd_net_),
            .in3(N__4578),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__9089),
            .ce(N__5052),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_9_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_9_4  (
            .in0(N__5079),
            .in1(N__4661),
            .in2(_gnd_net_),
            .in3(N__4575),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__9089),
            .ce(N__5052),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_9_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_9_5  (
            .in0(N__5086),
            .in1(N__4674),
            .in2(_gnd_net_),
            .in3(N__4572),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__9089),
            .ce(N__5052),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_9_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_9_6  (
            .in0(N__5080),
            .in1(N__4686),
            .in2(_gnd_net_),
            .in3(N__4569),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__9089),
            .ce(N__5052),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_9_7  (
            .in0(N__5087),
            .in1(N__4647),
            .in2(_gnd_net_),
            .in3(N__4566),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9089),
            .ce(N__5052),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_10_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_10_0  (
            .in0(N__5166),
            .in1(N__7920),
            .in2(N__7251),
            .in3(N__7113),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_282_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_10_1 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_10_1  (
            .in0(N__7114),
            .in1(N__4623),
            .in2(N__4563),
            .in3(N__6116),
            .lcout(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_7_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_7_10_2 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_7_10_2  (
            .in0(N__7290),
            .in1(N__6910),
            .in2(N__7252),
            .in3(N__5577),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_265_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_10_3 .LUT_INIT=16'b1111111111111001;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_10_3  (
            .in0(N__7049),
            .in1(N__7237),
            .in2(N__4560),
            .in3(N__6795),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_7_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_7_10_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_7_10_4  (
            .in0(N__4700),
            .in1(N__4710),
            .in2(N__4704),
            .in3(N__5530),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9094),
            .ce(),
            .sr(N__9969));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_7_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_7_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_7_10_5  (
            .in0(N__4685),
            .in1(N__4673),
            .in2(N__4662),
            .in3(N__4646),
            .lcout(\U712_CHIP_RAM.N_208 ),
            .ltout(\U712_CHIP_RAM.N_208_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_7_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_7_10_6 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(N__4635),
            .in2(N__4629),
            .in3(N__6082),
            .lcout(\U712_CHIP_RAM.N_398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIP7DI_LC_7_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIP7DI_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIP7DI_LC_7_11_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIP7DI_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__5576),
            .in2(_gnd_net_),
            .in3(N__7230),
            .lcout(\U712_CHIP_RAM.N_245 ),
            .ltout(\U712_CHIP_RAM.N_245_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_7_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_7_11_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_7_11_3  (
            .in0(N__6929),
            .in1(N__7048),
            .in2(N__4626),
            .in3(N__7913),
            .lcout(\U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_7_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_7_11_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_7_11_5  (
            .in0(N__4617),
            .in1(N__4602),
            .in2(_gnd_net_),
            .in3(N__8206),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_7_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_7_11_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_7_11_6  (
            .in0(N__7914),
            .in1(N__8207),
            .in2(N__4587),
            .in3(N__9330),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_LC_7_12_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_LC_7_12_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_LC_7_12_1  (
            .in0(N__4851),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4868),
            .lcout(\U712_BYTE_ENABLE.N_322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_7_12_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_7_12_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_7_12_3  (
            .in0(N__5458),
            .in1(N__5381),
            .in2(_gnd_net_),
            .in3(N__6757),
            .lcout(\U712_BYTE_ENABLE.N_327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_7_12_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_7_12_4 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_7_12_4  (
            .in0(N__7925),
            .in1(N__8413),
            .in2(_gnd_net_),
            .in3(N__4904),
            .lcout(\U712_BYTE_ENABLE.N_319 ),
            .ltout(\U712_BYTE_ENABLE.N_319_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_43_i_LC_7_12_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_43_i_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_43_i_LC_7_12_5 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \U712_BYTE_ENABLE.N_43_i_LC_7_12_5  (
            .in0(N__4976),
            .in1(N__5418),
            .in2(N__4932),
            .in3(N__4857),
            .lcout(N_43_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_1_LC_7_13_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_1_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_1_LC_7_13_1 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_1_LC_7_13_1  (
            .in0(N__4908),
            .in1(N__8453),
            .in2(_gnd_net_),
            .in3(N__7926),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_1_LC_7_13_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_1_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_1_LC_7_13_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_1_LC_7_13_5  (
            .in0(N__4835),
            .in1(N__8455),
            .in2(_gnd_net_),
            .in3(N__7930),
            .lcout(\U712_BYTE_ENABLE.N_321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_0_LC_7_13_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_0_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_0_LC_7_13_6 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_0_0_LC_7_13_6  (
            .in0(N__8454),
            .in1(N__4834),
            .in2(N__7932),
            .in3(N__5408),
            .lcout(\U712_BYTE_ENABLE.un1_CLMBEn_i_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_6_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_6_4 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_6_4 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_6_4  (
            .in0(N__8703),
            .in1(N__4743),
            .in2(_gnd_net_),
            .in3(N__4782),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9079),
            .ce(N__4722),
            .sr(N__9995));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_7_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_7_2 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_7_2  (
            .in0(N__8699),
            .in1(N__4780),
            .in2(N__4764),
            .in3(N__4741),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_233_i_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_7_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_7_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4725),
            .in3(N__10020),
            .lcout(\U712_CYCLE_TERM.N_233_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_7_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_7_4 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_7_4  (
            .in0(N__6418),
            .in1(_gnd_net_),
            .in2(N__6372),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a3_0_a3_LC_8_7_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a3_0_a3_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a3_0_a3_LC_8_7_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a3_0_a3_LC_8_7_5  (
            .in0(N__5310),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7919),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_8_8_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__7180),
            .in2(_gnd_net_),
            .in3(N__7008),
            .lcout(\U712_CHIP_RAM.N_209 ),
            .ltout(\U712_CHIP_RAM.N_209_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_8_8_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_8_8_1  (
            .in0(N__6240),
            .in1(N__7275),
            .in2(N__4989),
            .in3(N__7115),
            .lcout(\U712_CHIP_RAM.N_359 ),
            .ltout(\U712_CHIP_RAM.N_359_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_8_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_8_8_2 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_8_8_2  (
            .in0(N__5761),
            .in1(_gnd_net_),
            .in2(N__4986),
            .in3(N__5921),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_8_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_8_8_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_8_8_3 .LUT_INIT=16'b1010110011111100;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_8_8_3  (
            .in0(N__6128),
            .in1(N__5436),
            .in2(N__4983),
            .in3(N__9345),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9083),
            .ce(),
            .sr(N__9979));
    defparam \U712_CHIP_RAM.REFRESH_RNILCLN6_LC_8_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNILCLN6_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNILCLN6_LC_8_8_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNILCLN6_LC_8_8_4  (
            .in0(N__5760),
            .in1(N__5809),
            .in2(N__5681),
            .in3(N__5028),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_8_5 .LUT_INIT=16'b1000100011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_8_5  (
            .in0(N__6241),
            .in1(N__7021),
            .in2(_gnd_net_),
            .in3(N__6163),
            .lcout(\U712_CHIP_RAM.N_226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_8_9_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_8_9_0  (
            .in0(N__7239),
            .in1(N__5541),
            .in2(N__6129),
            .in3(N__5529),
            .lcout(\U712_CHIP_RAM.N_290 ),
            .ltout(\U712_CHIP_RAM.N_290_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_8_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_8_9_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_8_9_1  (
            .in0(N__5962),
            .in1(N__8681),
            .in2(N__4980),
            .in3(N__5016),
            .lcout(\U712_CHIP_RAM.N_181 ),
            .ltout(\U712_CHIP_RAM.N_181_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_9_2 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_9_2  (
            .in0(N__5964),
            .in1(N__5196),
            .in2(N__5118),
            .in3(N__5115),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9087),
            .ce(N__5051),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_9_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__6220),
            .in2(_gnd_net_),
            .in3(N__7097),
            .lcout(\U712_CHIP_RAM.N_216 ),
            .ltout(\U712_CHIP_RAM.N_216_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_8_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_8_9_4 .LUT_INIT=16'b0000111000001100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_8_9_4  (
            .in0(N__7238),
            .in1(N__5148),
            .in2(N__5103),
            .in3(N__5100),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_2_LC_8_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_2_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_2_LC_8_9_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_2_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__5559),
            .in2(_gnd_net_),
            .in3(N__5164),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_9_7 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_9_7  (
            .in0(N__5094),
            .in1(N__8680),
            .in2(N__5088),
            .in3(N__5941),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9087),
            .ce(N__5051),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_SYNC_RNI2HJQ_1_LC_8_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_RNI2HJQ_1_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_RNI2HJQ_1_LC_8_10_0 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_SYNC_RNI2HJQ_1_LC_8_10_0  (
            .in0(N__5142),
            .in1(N__6335),
            .in2(_gnd_net_),
            .in3(N__6440),
            .lcout(\U712_CHIP_RAM.N_204 ),
            .ltout(\U712_CHIP_RAM.N_204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIRS4M1_LC_8_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIRS4M1_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIRS4M1_LC_8_10_1 .LUT_INIT=16'b0000110011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIRS4M1_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__8675),
            .in2(N__5031),
            .in3(N__5827),
            .lcout(\U712_CHIP_RAM.N_279_1 ),
            .ltout(\U712_CHIP_RAM.N_279_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIGKJ14_LC_8_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIGKJ14_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIGKJ14_LC_8_10_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIGKJ14_LC_8_10_2  (
            .in0(N__5793),
            .in1(N__5758),
            .in2(N__5019),
            .in3(N__5165),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIAQERA_LC_8_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIAQERA_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIAQERA_LC_8_10_3 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIAQERA_LC_8_10_3  (
            .in0(N__5531),
            .in1(N__5015),
            .in2(N__5004),
            .in3(N__8676),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI2B8VE_3_LC_8_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI2B8VE_3_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI2B8VE_3_LC_8_10_4 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI2B8VE_3_LC_8_10_4  (
            .in0(N__7179),
            .in1(N__5532),
            .in2(N__5169),
            .in3(N__6837),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_LC_8_10_5 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_LC_8_10_5  (
            .in0(N__6990),
            .in1(_gnd_net_),
            .in2(N__6912),
            .in3(N__6077),
            .lcout(\U712_CHIP_RAM.N_393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_8_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_8_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_8_10_6  (
            .in0(N__7178),
            .in1(N__6991),
            .in2(N__6117),
            .in3(N__6884),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_SYNC_1_LC_8_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_1_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_1_LC_8_10_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_SYNC_1_LC_8_10_7  (
            .in0(N__6336),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.REFRESH_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9090),
            .ce(),
            .sr(N__9960));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_11_1 .LUT_INIT=16'b1000111110001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_11_1  (
            .in0(N__7043),
            .in1(N__7286),
            .in2(N__6255),
            .in3(N__7244),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_11_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_11_2  (
            .in0(N__7243),
            .in1(N__6245),
            .in2(N__6933),
            .in3(N__7042),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIJC372_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIJC372_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIJC372_LC_8_11_3 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIJC372_LC_8_11_3  (
            .in0(N__7039),
            .in1(N__6925),
            .in2(N__6253),
            .in3(N__7285),
            .lcout(\U712_CHIP_RAM.N_227 ),
            .ltout(\U712_CHIP_RAM.N_227_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_11_4 .LUT_INIT=16'b1111111011111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_11_4  (
            .in0(N__6783),
            .in1(N__6121),
            .in2(N__5136),
            .in3(N__5133),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9095),
            .ce(N__6284),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_11_5 .LUT_INIT=16'b1101110001010100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_11_5  (
            .in0(N__7041),
            .in1(N__6120),
            .in2(N__6254),
            .in3(N__5124),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_0_LC_8_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_0_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_0_LC_8_11_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_0_LC_8_11_6  (
            .in0(N__6119),
            .in1(N__7112),
            .in2(N__7253),
            .in3(N__7040),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__6924),
            .in2(_gnd_net_),
            .in3(N__6118),
            .lcout(\U712_CHIP_RAM.N_303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_0_0_LC_8_12_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_0_0_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_0_0_LC_8_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_0_0_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__5448),
            .in2(_gnd_net_),
            .in3(N__6756),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0 ),
            .ltout(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_42_i_LC_8_12_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_42_i_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_42_i_LC_8_12_4 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_42_i_LC_8_12_4  (
            .in0(N__5407),
            .in1(N__5391),
            .in2(N__5385),
            .in3(N__5371),
            .lcout(N_42_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_8_15_4 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_8_15_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__6765),
            .in2(_gnd_net_),
            .in3(N__5306),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_5_3  (
            .in0(N__5253),
            .in1(N__5235),
            .in2(_gnd_net_),
            .in3(N__8203),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_9_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_9_6_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_9_6_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_LC_9_6_0  (
            .in0(N__6127),
            .in1(N__7246),
            .in2(N__7050),
            .in3(N__7128),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9076),
            .ce(N__5175),
            .sr(N__9989));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__6566),
            .in2(_gnd_net_),
            .in3(N__6126),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_LC_9_7_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(N__10019),
            .in2(_gnd_net_),
            .in3(N__5184),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_7_5  (
            .in0(N__5625),
            .in1(N__5607),
            .in2(_gnd_net_),
            .in3(N__8204),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_9_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_9_7_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_9_7_6  (
            .in0(N__8205),
            .in1(N__7888),
            .in2(N__5592),
            .in3(N__9387),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_8_0 .LUT_INIT=16'b0101010111110000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_9_8_0  (
            .in0(N__5589),
            .in1(_gnd_net_),
            .in2(N__5575),
            .in3(N__5943),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9080),
            .ce(),
            .sr(N__9970));
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_9_8_2 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_LC_9_8_2  (
            .in0(N__6723),
            .in1(N__5677),
            .in2(N__5766),
            .in3(N__5502),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9080),
            .ce(),
            .sr(N__9970));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICREN6_LC_9_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICREN6_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICREN6_LC_9_8_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICREN6_LC_9_8_3  (
            .in0(N__5676),
            .in1(N__5762),
            .in2(_gnd_net_),
            .in3(N__5978),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIMTA11_LC_9_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIMTA11_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIMTA11_LC_9_8_4 .LUT_INIT=16'b1100110000100010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIMTA11_LC_9_8_4  (
            .in0(N__5565),
            .in1(N__7009),
            .in2(_gnd_net_),
            .in3(N__6931),
            .lcout(\U712_CHIP_RAM.N_205 ),
            .ltout(\U712_CHIP_RAM.N_205_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_0_LC_9_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_0_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_0_LC_9_8_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_0_LC_9_8_5  (
            .in0(N__7245),
            .in1(N__6107),
            .in2(N__5535),
            .in3(N__5528),
            .lcout(\U712_CHIP_RAM.N_291 ),
            .ltout(\U712_CHIP_RAM.N_291_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_8_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_8_6  (
            .in0(N__5979),
            .in1(N__5675),
            .in2(N__5496),
            .in3(N__10018),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI06U42_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI06U42_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI06U42_LC_9_9_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI06U42_LC_9_9_1  (
            .in0(N__5792),
            .in1(N__5828),
            .in2(N__5493),
            .in3(N__5744),
            .lcout(\U712_CHIP_RAM.N_395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_1_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_1_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_1_LC_9_9_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_1_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__6913),
            .in2(_gnd_net_),
            .in3(N__6081),
            .lcout(\U712_CHIP_RAM.N_342 ),
            .ltout(\U712_CHIP_RAM.N_342_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_9_9_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_9_9_3  (
            .in0(N__7217),
            .in1(N__7031),
            .in2(N__6006),
            .in3(N__7129),
            .lcout(\U712_CHIP_RAM.N_352 ),
            .ltout(\U712_CHIP_RAM.N_352_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_9_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_1_LC_9_9_4  (
            .in0(N__10358),
            .in1(N__6003),
            .in2(N__5982),
            .in3(N__5977),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_293_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_9_9_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_0_LC_9_9_5  (
            .in0(N__5963),
            .in1(N__5745),
            .in2(N__5946),
            .in3(N__8952),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.BANK0_LC_9_9_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \U712_CHIP_RAM.BANK0_LC_9_9_6  (
            .in0(N__5894),
            .in1(N__5942),
            .in2(N__5925),
            .in3(N__5922),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9084),
            .ce(),
            .sr(N__9961));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_10_0 .LUT_INIT=16'b0001111100010001;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_10_0  (
            .in0(N__5883),
            .in1(N__5850),
            .in2(N__7902),
            .in3(N__5829),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9088),
            .ce(),
            .sr(N__9953));
    defparam \U712_CHIP_RAM.REFRESH_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_9_10_1 .LUT_INIT=16'b1111001111111011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_9_10_1  (
            .in0(N__7704),
            .in1(N__7761),
            .in2(N__8538),
            .in3(N__7422),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9088),
            .ce(),
            .sr(N__9953));
    defparam \U712_CHIP_RAM.DBDIR_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_10_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_10_2 .LUT_INIT=16'b0111010011110000;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_9_10_2  (
            .in0(N__6701),
            .in1(N__5759),
            .in2(N__5642),
            .in3(N__5682),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9088),
            .ce(),
            .sr(N__9953));
    defparam DBR_SYNC_1_LC_9_10_3.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_9_10_3.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_9_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_9_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6468),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9088),
            .ce(),
            .sr(N__9953));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_10_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6368),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9088),
            .ce(),
            .sr(N__9953));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_10_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__8825),
            .in2(_gnd_net_),
            .in3(N__6399),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9088),
            .ce(),
            .sr(N__9953));
    defparam \U712_CHIP_RAM.REFRESH_SYNC_0_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_0_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_0_LC_9_10_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.REFRESH_SYNC_0_LC_9_10_7  (
            .in0(N__9264),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6354),
            .lcout(\U712_CHIP_RAM.REFRESH_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9088),
            .ce(),
            .sr(N__9953));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_11_2  (
            .in0(N__6327),
            .in1(N__6147),
            .in2(N__6321),
            .in3(N__6781),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9091),
            .ce(N__6285),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_11_5 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_11_5  (
            .in0(N__6782),
            .in1(N__6309),
            .in2(N__6174),
            .in3(N__6012),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9091),
            .ce(N__6285),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_11_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_11_6  (
            .in0(N__6297),
            .in1(N__6291),
            .in2(_gnd_net_),
            .in3(N__6780),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9091),
            .ce(N__6285),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_12_2 .LUT_INIT=16'b0000111111110001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_12_2  (
            .in0(N__6252),
            .in1(N__6932),
            .in2(N__6139),
            .in3(N__6170),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_12_4 .LUT_INIT=16'b1111111110010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_12_4  (
            .in0(N__7250),
            .in1(N__7044),
            .in2(N__6140),
            .in3(N__6018),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR4F93_1_LC_9_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR4F93_1_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR4F93_1_LC_9_12_5 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIR4F93_1_LC_9_12_5  (
            .in0(N__8674),
            .in1(N__6794),
            .in2(_gnd_net_),
            .in3(N__7131),
            .lcout(\U712_CHIP_RAM.N_241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_9_16_7 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_9_16_7 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_9_16_7  (
            .in0(N__6754),
            .in1(N__6688),
            .in2(_gnd_net_),
            .in3(N__6639),
            .lcout(N_256),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_5_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_5_4  (
            .in0(N__7915),
            .in1(N__6588),
            .in2(N__8237),
            .in3(N__9408),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_10_5_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_5_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_5_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_10_6_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_10_6_0  (
            .in0(N__7983),
            .in1(N__6555),
            .in2(N__7931),
            .in3(N__9234),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9075),
            .ce(N__8988),
            .sr(N__9980));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_10_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_10_7_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_10_7_2  (
            .in0(N__9221),
            .in1(N__9678),
            .in2(N__9189),
            .in3(N__6513),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9077),
            .ce(N__8983),
            .sr(N__9971));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_7_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_10_7_3  (
            .in0(N__7299),
            .in1(N__6474),
            .in2(_gnd_net_),
            .in3(N__7332),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9077),
            .ce(N__8983),
            .sr(N__9971));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_8_0 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_8_0  (
            .in0(N__7845),
            .in1(N__7497),
            .in2(N__8219),
            .in3(N__9357),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_8_1 .LUT_INIT=16'b0000111101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_8_1  (
            .in0(N__7881),
            .in1(N__9419),
            .in2(N__8220),
            .in3(N__9162),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_8_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_8_2  (
            .in0(N__7844),
            .in1(N__7326),
            .in2(_gnd_net_),
            .in3(N__9396),
            .lcout(\U712_CHIP_RAM.N_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_10_8_3 .LUT_INIT=16'b0000001100110001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_10_8_3  (
            .in0(N__8047),
            .in1(N__8080),
            .in2(N__8307),
            .in3(N__8187),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_10_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_10_8_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_10_8_4  (
            .in0(_gnd_net_),
            .in1(N__8300),
            .in2(_gnd_net_),
            .in3(N__8046),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_5 .LUT_INIT=16'b0011111100110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(N__8191),
            .in2(N__7308),
            .in3(N__7305),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_8_6 .LUT_INIT=16'b0011111100111011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_8_6  (
            .in0(N__9420),
            .in1(N__8193),
            .in2(N__9178),
            .in3(N__7880),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_9_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_9_0  (
            .in0(N__7030),
            .in1(N__7284),
            .in2(N__7254),
            .in3(N__7130),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9081),
            .ce(N__7062),
            .sr(N__9954));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJOND1_1_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJOND1_1_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJOND1_1_LC_10_9_1 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIJOND1_1_LC_10_9_1  (
            .in0(N__8662),
            .in1(N__7029),
            .in2(_gnd_net_),
            .in3(N__6930),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_9_3  (
            .in0(N__6825),
            .in1(N__6810),
            .in2(_gnd_net_),
            .in3(N__8192),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_10_0 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_10_0  (
            .in0(N__8164),
            .in1(N__8304),
            .in2(_gnd_net_),
            .in3(N__8028),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_10_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_10_3  (
            .in0(N__7530),
            .in1(N__7512),
            .in2(_gnd_net_),
            .in3(N__8163),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_4  (
            .in0(N__8165),
            .in1(N__7488),
            .in2(_gnd_net_),
            .in3(N__7473),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_10_6  (
            .in0(N__8162),
            .in1(N__7455),
            .in2(_gnd_net_),
            .in3(N__7434),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_11_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_11_2  (
            .in0(N__8071),
            .in1(N__8140),
            .in2(N__8034),
            .in3(N__8282),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_11_3 .LUT_INIT=16'b0001111100111111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_11_3  (
            .in0(N__7751),
            .in1(N__7718),
            .in2(N__7683),
            .in3(N__7733),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_11_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_11_6_0 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_11_6_0  (
            .in0(N__9528),
            .in1(N__7982),
            .in2(N__7924),
            .in3(N__7416),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9070),
            .ce(N__8984),
            .sr(N__9972));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_6_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_11_6_4  (
            .in0(N__9218),
            .in1(N__9789),
            .in2(N__9192),
            .in3(N__7374),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9070),
            .ce(N__8984),
            .sr(N__9972));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_6_6 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_11_6_6  (
            .in0(N__9217),
            .in1(N__9642),
            .in2(N__9191),
            .in3(N__7539),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9070),
            .ce(N__8984),
            .sr(N__9972));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_7_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__10017),
            .in2(_gnd_net_),
            .in3(N__7650),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_7_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__7889),
            .in2(_gnd_net_),
            .in3(N__8221),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_8_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_11_8_3  (
            .in0(N__9219),
            .in1(N__9732),
            .in2(N__9188),
            .in3(N__7644),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9078),
            .ce(N__8993),
            .sr(N__9955));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_8_6 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_11_8_6  (
            .in0(N__9177),
            .in1(N__9220),
            .in2(N__9846),
            .in3(N__7563),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9078),
            .ce(N__8993),
            .sr(N__9955));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_11_8_7  (
            .in0(N__7551),
            .in1(N__7767),
            .in2(_gnd_net_),
            .in3(N__7599),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9078),
            .ce(N__8993),
            .sr(N__9955));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_9_2 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_9_2  (
            .in0(N__7857),
            .in1(N__7569),
            .in2(N__8239),
            .in3(N__9366),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_9_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_9_3  (
            .in0(N__8231),
            .in1(N__7557),
            .in2(N__7923),
            .in3(N__9318),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_9_5 .LUT_INIT=16'b1101111111010101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_9_5  (
            .in0(N__7969),
            .in1(N__7956),
            .in2(N__7921),
            .in3(N__10152),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_9_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_9_6  (
            .in0(N__7856),
            .in1(N__7545),
            .in2(N__8238),
            .in3(N__9375),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_9_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_9_7  (
            .in0(N__7970),
            .in1(N__7955),
            .in2(N__7922),
            .in3(N__10151),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_10_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__8555),
            .in2(_gnd_net_),
            .in3(N__7664),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_11_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_11_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__7752),
            .in2(_gnd_net_),
            .in3(N__7737),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__8862),
            .ce(),
            .sr(N__8517));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_11_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_11_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__7734),
            .in2(_gnd_net_),
            .in3(N__7722),
            .lcout(\U712_CHIP_RAM.REFRESH5lto1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__8862),
            .ce(),
            .sr(N__8517));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_11_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_11_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__7719),
            .in2(_gnd_net_),
            .in3(N__7707),
            .lcout(\U712_CHIP_RAM.REFRESH5lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__8862),
            .ce(),
            .sr(N__8517));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_11_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_11_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__7700),
            .in2(_gnd_net_),
            .in3(N__7686),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__8862),
            .ce(),
            .sr(N__8517));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_11_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_11_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__7682),
            .in2(_gnd_net_),
            .in3(N__7668),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__8862),
            .ce(),
            .sr(N__8517));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_11_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_11_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__7665),
            .in2(_gnd_net_),
            .in3(N__7653),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__8862),
            .ce(),
            .sr(N__8517));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_11_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_11_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__8556),
            .in2(_gnd_net_),
            .in3(N__8544),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__8862),
            .ce(),
            .sr(N__8517));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_11_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_11_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(N__8531),
            .in2(_gnd_net_),
            .in3(N__8541),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8862),
            .ce(),
            .sr(N__8517));
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_11_14_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_11_14_2 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_11_14_2  (
            .in0(N__8489),
            .in1(N__8463),
            .in2(_gnd_net_),
            .in3(N__8423),
            .lcout(un1_LDSn_i_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_11_15_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_11_15_6 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_11_15_6  (
            .in0(N__8490),
            .in1(N__8462),
            .in2(_gnd_net_),
            .in3(N__8424),
            .lcout(un1_UDSn_i_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RASn_LC_12_3_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_12_3_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_12_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8305),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9066),
            .ce(),
            .sr(N__9986));
    defparam \U712_CHIP_RAM.CRCSn_LC_12_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_12_4_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_12_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_12_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8090),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9067),
            .ce(),
            .sr(N__9978));
    defparam \U712_CHIP_RAM.WEn_LC_12_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_12_5_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_12_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8048),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9068),
            .ce(),
            .sr(N__9968));
    defparam \U712_CHIP_RAM.CASn_LC_12_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_12_5_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_12_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_12_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8250),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9068),
            .ce(),
            .sr(N__9968));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_6_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_12_6_1  (
            .in0(N__8306),
            .in1(N__8246),
            .in2(N__8091),
            .in3(N__8055),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9069),
            .ce(N__8989),
            .sr(N__9958));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_7_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_7_3  (
            .in0(N__9629),
            .in1(N__10359),
            .in2(_gnd_net_),
            .in3(N__9260),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10132),
            .ce(N__10086),
            .sr(N__9952));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_8_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_12_8_7  (
            .in0(N__9222),
            .in1(N__9777),
            .in2(N__9190),
            .in3(N__9126),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9071),
            .ce(N__8994),
            .sr(N__9949));
    defparam \U712_CHIP_RAM.DMA_A20_LC_12_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A20_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A20_LC_12_9_2 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A20_LC_12_9_2  (
            .in0(N__10346),
            .in1(N__8937),
            .in2(N__9628),
            .in3(N__8951),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .ce(),
            .sr(N__9947));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS10_LC_12_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS10_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS10_LC_12_10_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS10_LC_12_10_1  (
            .in0(N__8924),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10140),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10 ),
            .ltout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_12_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_12_10_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8931),
            .in3(N__10015),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_10_7 .LUT_INIT=16'b1010111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_10_7  (
            .in0(N__10016),
            .in1(_gnd_net_),
            .in2(N__8928),
            .in3(N__8883),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pll_RNI8MQ3_LC_12_11_4.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_12_11_4.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_12_11_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 pll_RNI8MQ3_LC_12_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8821),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_5.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_5.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8704),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_7  (
            .in0(N__10338),
            .in1(N__9576),
            .in2(_gnd_net_),
            .in3(N__9829),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__9306),
            .sr(N__9962));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_7  (
            .in0(N__10411),
            .in1(N__10347),
            .in2(_gnd_net_),
            .in3(N__9828),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__9305),
            .sr(N__9956));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_0  (
            .in0(N__10412),
            .in1(N__10342),
            .in2(_gnd_net_),
            .in3(N__10198),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__9291),
            .sr(N__9950));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_9_4  (
            .in0(N__9472),
            .in1(N__10340),
            .in2(_gnd_net_),
            .in3(N__9515),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__9291),
            .sr(N__9950));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_5  (
            .in0(N__9556),
            .in1(_gnd_net_),
            .in2(N__10357),
            .in3(N__9618),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__9291),
            .sr(N__9950));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_6  (
            .in0(N__9768),
            .in1(N__10341),
            .in2(_gnd_net_),
            .in3(N__9516),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__9291),
            .sr(N__9950));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0  (
            .in0(N__9473),
            .in1(_gnd_net_),
            .in2(N__9666),
            .in3(N__10339),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__9290),
            .sr(N__9948));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_11_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_11_1  (
            .in0(N__9720),
            .in1(N__10303),
            .in2(_gnd_net_),
            .in3(N__9764),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__9292),
            .sr(N__9946));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_4  (
            .in0(N__10304),
            .in1(N__9721),
            .in2(_gnd_net_),
            .in3(N__10188),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__9292),
            .sr(N__9946));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_1  (
            .in0(N__10299),
            .in1(N__9575),
            .in2(_gnd_net_),
            .in3(N__9831),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10133),
            .ce(N__10090),
            .sr(N__9973));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_3  (
            .in0(N__10298),
            .in1(N__10413),
            .in2(_gnd_net_),
            .in3(N__9830),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10133),
            .ce(N__10090),
            .sr(N__9973));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_0  (
            .in0(N__10296),
            .in1(N__9723),
            .in2(_gnd_net_),
            .in3(N__9763),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10130),
            .ce(N__10092),
            .sr(N__9963));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_8_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_8_3  (
            .in0(N__9762),
            .in1(N__10295),
            .in2(_gnd_net_),
            .in3(N__9514),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10130),
            .ce(N__10092),
            .sr(N__9963));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_9_4  (
            .in0(N__10200),
            .in1(N__10353),
            .in2(_gnd_net_),
            .in3(N__9722),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10129),
            .ce(N__10091),
            .sr(N__9957));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_10_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_10_0  (
            .in0(N__9465),
            .in1(N__10294),
            .in2(_gnd_net_),
            .in3(N__9662),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10128),
            .ce(N__10064),
            .sr(N__9951));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_0  (
            .in0(N__10297),
            .in1(N__9630),
            .in2(_gnd_net_),
            .in3(N__9574),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10135),
            .ce(N__10098),
            .sr(N__9981));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_3  (
            .in0(N__10352),
            .in1(N__9508),
            .in2(_gnd_net_),
            .in3(N__9477),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10134),
            .ce(N__10093),
            .sr(N__9974));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_9_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_9_1  (
            .in0(N__10404),
            .in1(N__10351),
            .in2(_gnd_net_),
            .in3(N__10199),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10131),
            .ce(N__10097),
            .sr(N__9964));
endmodule // U712_TOP

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     May 8 2025 19:59:06

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    CMA,
    DRA,
    DA,
    A,
    DBRn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    TCIn,
    TBIn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    input [1:0] SIZ;
    output [10:0] CMA;
    input [9:0] DRA;
    output [2:0] DA;
    input [20:0] A;
    input DBRn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    output TCIn;
    output TBIn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__12817;
    wire N__12816;
    wire N__12815;
    wire N__12808;
    wire N__12807;
    wire N__12806;
    wire N__12799;
    wire N__12798;
    wire N__12797;
    wire N__12790;
    wire N__12789;
    wire N__12788;
    wire N__12781;
    wire N__12780;
    wire N__12779;
    wire N__12772;
    wire N__12771;
    wire N__12770;
    wire N__12763;
    wire N__12762;
    wire N__12761;
    wire N__12754;
    wire N__12753;
    wire N__12752;
    wire N__12745;
    wire N__12744;
    wire N__12743;
    wire N__12736;
    wire N__12735;
    wire N__12734;
    wire N__12727;
    wire N__12726;
    wire N__12725;
    wire N__12718;
    wire N__12717;
    wire N__12716;
    wire N__12709;
    wire N__12708;
    wire N__12707;
    wire N__12700;
    wire N__12699;
    wire N__12698;
    wire N__12691;
    wire N__12690;
    wire N__12689;
    wire N__12682;
    wire N__12681;
    wire N__12680;
    wire N__12673;
    wire N__12672;
    wire N__12671;
    wire N__12664;
    wire N__12663;
    wire N__12662;
    wire N__12655;
    wire N__12654;
    wire N__12653;
    wire N__12646;
    wire N__12645;
    wire N__12644;
    wire N__12637;
    wire N__12636;
    wire N__12635;
    wire N__12628;
    wire N__12627;
    wire N__12626;
    wire N__12619;
    wire N__12618;
    wire N__12617;
    wire N__12610;
    wire N__12609;
    wire N__12608;
    wire N__12601;
    wire N__12600;
    wire N__12599;
    wire N__12592;
    wire N__12591;
    wire N__12590;
    wire N__12583;
    wire N__12582;
    wire N__12581;
    wire N__12574;
    wire N__12573;
    wire N__12572;
    wire N__12565;
    wire N__12564;
    wire N__12563;
    wire N__12556;
    wire N__12555;
    wire N__12554;
    wire N__12547;
    wire N__12546;
    wire N__12545;
    wire N__12538;
    wire N__12537;
    wire N__12536;
    wire N__12529;
    wire N__12528;
    wire N__12527;
    wire N__12520;
    wire N__12519;
    wire N__12518;
    wire N__12511;
    wire N__12510;
    wire N__12509;
    wire N__12502;
    wire N__12501;
    wire N__12500;
    wire N__12493;
    wire N__12492;
    wire N__12491;
    wire N__12484;
    wire N__12483;
    wire N__12482;
    wire N__12475;
    wire N__12474;
    wire N__12473;
    wire N__12466;
    wire N__12465;
    wire N__12464;
    wire N__12457;
    wire N__12456;
    wire N__12455;
    wire N__12448;
    wire N__12447;
    wire N__12446;
    wire N__12439;
    wire N__12438;
    wire N__12437;
    wire N__12430;
    wire N__12429;
    wire N__12428;
    wire N__12421;
    wire N__12420;
    wire N__12419;
    wire N__12412;
    wire N__12411;
    wire N__12410;
    wire N__12403;
    wire N__12402;
    wire N__12401;
    wire N__12394;
    wire N__12393;
    wire N__12392;
    wire N__12385;
    wire N__12384;
    wire N__12383;
    wire N__12376;
    wire N__12375;
    wire N__12374;
    wire N__12367;
    wire N__12366;
    wire N__12365;
    wire N__12358;
    wire N__12357;
    wire N__12356;
    wire N__12349;
    wire N__12348;
    wire N__12347;
    wire N__12340;
    wire N__12339;
    wire N__12338;
    wire N__12331;
    wire N__12330;
    wire N__12329;
    wire N__12322;
    wire N__12321;
    wire N__12320;
    wire N__12313;
    wire N__12312;
    wire N__12311;
    wire N__12304;
    wire N__12303;
    wire N__12302;
    wire N__12295;
    wire N__12294;
    wire N__12293;
    wire N__12286;
    wire N__12285;
    wire N__12284;
    wire N__12277;
    wire N__12276;
    wire N__12275;
    wire N__12268;
    wire N__12267;
    wire N__12266;
    wire N__12259;
    wire N__12258;
    wire N__12257;
    wire N__12250;
    wire N__12249;
    wire N__12248;
    wire N__12241;
    wire N__12240;
    wire N__12239;
    wire N__12232;
    wire N__12231;
    wire N__12230;
    wire N__12223;
    wire N__12222;
    wire N__12221;
    wire N__12214;
    wire N__12213;
    wire N__12212;
    wire N__12205;
    wire N__12204;
    wire N__12203;
    wire N__12196;
    wire N__12195;
    wire N__12194;
    wire N__12187;
    wire N__12186;
    wire N__12185;
    wire N__12178;
    wire N__12177;
    wire N__12176;
    wire N__12169;
    wire N__12168;
    wire N__12167;
    wire N__12160;
    wire N__12159;
    wire N__12158;
    wire N__12151;
    wire N__12150;
    wire N__12149;
    wire N__12142;
    wire N__12141;
    wire N__12140;
    wire N__12133;
    wire N__12132;
    wire N__12131;
    wire N__12124;
    wire N__12123;
    wire N__12122;
    wire N__12115;
    wire N__12114;
    wire N__12113;
    wire N__12106;
    wire N__12105;
    wire N__12104;
    wire N__12097;
    wire N__12096;
    wire N__12095;
    wire N__12088;
    wire N__12087;
    wire N__12086;
    wire N__12079;
    wire N__12078;
    wire N__12077;
    wire N__12070;
    wire N__12069;
    wire N__12068;
    wire N__12061;
    wire N__12060;
    wire N__12059;
    wire N__12052;
    wire N__12051;
    wire N__12050;
    wire N__12043;
    wire N__12042;
    wire N__12041;
    wire N__12034;
    wire N__12033;
    wire N__12032;
    wire N__12025;
    wire N__12024;
    wire N__12023;
    wire N__12016;
    wire N__12015;
    wire N__12014;
    wire N__12007;
    wire N__12006;
    wire N__12005;
    wire N__11998;
    wire N__11997;
    wire N__11996;
    wire N__11989;
    wire N__11988;
    wire N__11987;
    wire N__11980;
    wire N__11979;
    wire N__11978;
    wire N__11971;
    wire N__11970;
    wire N__11969;
    wire N__11952;
    wire N__11951;
    wire N__11950;
    wire N__11947;
    wire N__11944;
    wire N__11941;
    wire N__11938;
    wire N__11933;
    wire N__11928;
    wire N__11927;
    wire N__11924;
    wire N__11923;
    wire N__11920;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11910;
    wire N__11907;
    wire N__11904;
    wire N__11901;
    wire N__11896;
    wire N__11891;
    wire N__11888;
    wire N__11885;
    wire N__11882;
    wire N__11879;
    wire N__11874;
    wire N__11873;
    wire N__11872;
    wire N__11869;
    wire N__11868;
    wire N__11865;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11851;
    wire N__11850;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11836;
    wire N__11835;
    wire N__11830;
    wire N__11827;
    wire N__11824;
    wire N__11819;
    wire N__11816;
    wire N__11811;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11792;
    wire N__11787;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11767;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11755;
    wire N__11752;
    wire N__11747;
    wire N__11744;
    wire N__11741;
    wire N__11738;
    wire N__11733;
    wire N__11732;
    wire N__11731;
    wire N__11730;
    wire N__11727;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11707;
    wire N__11702;
    wire N__11699;
    wire N__11696;
    wire N__11693;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11673;
    wire N__11670;
    wire N__11669;
    wire N__11668;
    wire N__11667;
    wire N__11664;
    wire N__11661;
    wire N__11658;
    wire N__11655;
    wire N__11650;
    wire N__11647;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11622;
    wire N__11619;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11611;
    wire N__11610;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11587;
    wire N__11584;
    wire N__11579;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11565;
    wire N__11562;
    wire N__11559;
    wire N__11556;
    wire N__11553;
    wire N__11552;
    wire N__11549;
    wire N__11548;
    wire N__11545;
    wire N__11540;
    wire N__11539;
    wire N__11536;
    wire N__11535;
    wire N__11534;
    wire N__11533;
    wire N__11532;
    wire N__11531;
    wire N__11530;
    wire N__11529;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11501;
    wire N__11500;
    wire N__11497;
    wire N__11496;
    wire N__11495;
    wire N__11494;
    wire N__11491;
    wire N__11490;
    wire N__11487;
    wire N__11484;
    wire N__11481;
    wire N__11472;
    wire N__11471;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11455;
    wire N__11452;
    wire N__11447;
    wire N__11446;
    wire N__11445;
    wire N__11440;
    wire N__11435;
    wire N__11430;
    wire N__11419;
    wire N__11414;
    wire N__11409;
    wire N__11406;
    wire N__11403;
    wire N__11400;
    wire N__11397;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11383;
    wire N__11378;
    wire N__11373;
    wire N__11372;
    wire N__11371;
    wire N__11368;
    wire N__11365;
    wire N__11364;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11352;
    wire N__11349;
    wire N__11346;
    wire N__11339;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11321;
    wire N__11318;
    wire N__11315;
    wire N__11310;
    wire N__11307;
    wire N__11304;
    wire N__11301;
    wire N__11298;
    wire N__11295;
    wire N__11292;
    wire N__11289;
    wire N__11286;
    wire N__11285;
    wire N__11284;
    wire N__11283;
    wire N__11282;
    wire N__11281;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11261;
    wire N__11260;
    wire N__11259;
    wire N__11258;
    wire N__11257;
    wire N__11256;
    wire N__11255;
    wire N__11254;
    wire N__11253;
    wire N__11252;
    wire N__11251;
    wire N__11226;
    wire N__11223;
    wire N__11220;
    wire N__11219;
    wire N__11218;
    wire N__11217;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11197;
    wire N__11196;
    wire N__11195;
    wire N__11194;
    wire N__11193;
    wire N__11192;
    wire N__11191;
    wire N__11190;
    wire N__11189;
    wire N__11188;
    wire N__11187;
    wire N__11186;
    wire N__11185;
    wire N__11184;
    wire N__11181;
    wire N__11178;
    wire N__11177;
    wire N__11176;
    wire N__11175;
    wire N__11174;
    wire N__11173;
    wire N__11172;
    wire N__11171;
    wire N__11170;
    wire N__11169;
    wire N__11168;
    wire N__11167;
    wire N__11164;
    wire N__11163;
    wire N__11162;
    wire N__11161;
    wire N__11160;
    wire N__11159;
    wire N__11158;
    wire N__11157;
    wire N__11156;
    wire N__11155;
    wire N__11154;
    wire N__11151;
    wire N__11150;
    wire N__11149;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11046;
    wire N__11043;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11027;
    wire N__11024;
    wire N__11021;
    wire N__11016;
    wire N__11013;
    wire N__11010;
    wire N__11009;
    wire N__11008;
    wire N__11007;
    wire N__11006;
    wire N__11005;
    wire N__11004;
    wire N__11003;
    wire N__11002;
    wire N__11001;
    wire N__11000;
    wire N__10999;
    wire N__10998;
    wire N__10997;
    wire N__10996;
    wire N__10993;
    wire N__10990;
    wire N__10987;
    wire N__10982;
    wire N__10977;
    wire N__10972;
    wire N__10969;
    wire N__10966;
    wire N__10963;
    wire N__10962;
    wire N__10961;
    wire N__10960;
    wire N__10959;
    wire N__10958;
    wire N__10957;
    wire N__10956;
    wire N__10955;
    wire N__10954;
    wire N__10949;
    wire N__10948;
    wire N__10947;
    wire N__10944;
    wire N__10943;
    wire N__10942;
    wire N__10941;
    wire N__10938;
    wire N__10923;
    wire N__10920;
    wire N__10917;
    wire N__10914;
    wire N__10909;
    wire N__10902;
    wire N__10897;
    wire N__10894;
    wire N__10891;
    wire N__10888;
    wire N__10881;
    wire N__10878;
    wire N__10877;
    wire N__10876;
    wire N__10875;
    wire N__10870;
    wire N__10863;
    wire N__10860;
    wire N__10855;
    wire N__10844;
    wire N__10841;
    wire N__10840;
    wire N__10835;
    wire N__10834;
    wire N__10829;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10801;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10785;
    wire N__10782;
    wire N__10779;
    wire N__10776;
    wire N__10773;
    wire N__10770;
    wire N__10767;
    wire N__10766;
    wire N__10765;
    wire N__10764;
    wire N__10763;
    wire N__10762;
    wire N__10761;
    wire N__10760;
    wire N__10759;
    wire N__10758;
    wire N__10757;
    wire N__10756;
    wire N__10755;
    wire N__10754;
    wire N__10753;
    wire N__10752;
    wire N__10751;
    wire N__10750;
    wire N__10749;
    wire N__10748;
    wire N__10747;
    wire N__10746;
    wire N__10745;
    wire N__10744;
    wire N__10743;
    wire N__10742;
    wire N__10741;
    wire N__10740;
    wire N__10739;
    wire N__10738;
    wire N__10737;
    wire N__10736;
    wire N__10735;
    wire N__10734;
    wire N__10733;
    wire N__10732;
    wire N__10731;
    wire N__10730;
    wire N__10729;
    wire N__10728;
    wire N__10725;
    wire N__10724;
    wire N__10723;
    wire N__10722;
    wire N__10721;
    wire N__10720;
    wire N__10719;
    wire N__10718;
    wire N__10623;
    wire N__10620;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10600;
    wire N__10597;
    wire N__10594;
    wire N__10591;
    wire N__10584;
    wire N__10583;
    wire N__10580;
    wire N__10579;
    wire N__10576;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10563;
    wire N__10560;
    wire N__10557;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10545;
    wire N__10542;
    wire N__10539;
    wire N__10536;
    wire N__10531;
    wire N__10528;
    wire N__10525;
    wire N__10522;
    wire N__10517;
    wire N__10512;
    wire N__10509;
    wire N__10508;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10500;
    wire N__10499;
    wire N__10498;
    wire N__10495;
    wire N__10492;
    wire N__10489;
    wire N__10486;
    wire N__10479;
    wire N__10478;
    wire N__10471;
    wire N__10468;
    wire N__10465;
    wire N__10464;
    wire N__10463;
    wire N__10460;
    wire N__10455;
    wire N__10450;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10422;
    wire N__10421;
    wire N__10420;
    wire N__10417;
    wire N__10416;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10405;
    wire N__10402;
    wire N__10399;
    wire N__10398;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10365;
    wire N__10362;
    wire N__10359;
    wire N__10356;
    wire N__10353;
    wire N__10348;
    wire N__10345;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10329;
    wire N__10326;
    wire N__10323;
    wire N__10320;
    wire N__10317;
    wire N__10314;
    wire N__10311;
    wire N__10308;
    wire N__10305;
    wire N__10304;
    wire N__10303;
    wire N__10300;
    wire N__10297;
    wire N__10296;
    wire N__10293;
    wire N__10288;
    wire N__10285;
    wire N__10282;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10260;
    wire N__10257;
    wire N__10254;
    wire N__10251;
    wire N__10248;
    wire N__10245;
    wire N__10242;
    wire N__10241;
    wire N__10240;
    wire N__10235;
    wire N__10232;
    wire N__10231;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10212;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10195;
    wire N__10194;
    wire N__10189;
    wire N__10186;
    wire N__10183;
    wire N__10180;
    wire N__10175;
    wire N__10170;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10152;
    wire N__10149;
    wire N__10148;
    wire N__10147;
    wire N__10144;
    wire N__10139;
    wire N__10134;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10104;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10078;
    wire N__10073;
    wire N__10072;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10062;
    wire N__10059;
    wire N__10050;
    wire N__10047;
    wire N__10044;
    wire N__10041;
    wire N__10038;
    wire N__10035;
    wire N__10032;
    wire N__10029;
    wire N__10028;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10017;
    wire N__10014;
    wire N__10011;
    wire N__10008;
    wire N__10005;
    wire N__9996;
    wire N__9993;
    wire N__9990;
    wire N__9987;
    wire N__9984;
    wire N__9981;
    wire N__9978;
    wire N__9975;
    wire N__9972;
    wire N__9969;
    wire N__9966;
    wire N__9963;
    wire N__9960;
    wire N__9957;
    wire N__9954;
    wire N__9951;
    wire N__9948;
    wire N__9945;
    wire N__9942;
    wire N__9939;
    wire N__9936;
    wire N__9933;
    wire N__9930;
    wire N__9927;
    wire N__9924;
    wire N__9921;
    wire N__9920;
    wire N__9917;
    wire N__9912;
    wire N__9909;
    wire N__9906;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9882;
    wire N__9879;
    wire N__9876;
    wire N__9873;
    wire N__9872;
    wire N__9871;
    wire N__9870;
    wire N__9869;
    wire N__9868;
    wire N__9867;
    wire N__9860;
    wire N__9855;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9835;
    wire N__9832;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9807;
    wire N__9804;
    wire N__9801;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9793;
    wire N__9792;
    wire N__9791;
    wire N__9790;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9776;
    wire N__9775;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9747;
    wire N__9744;
    wire N__9735;
    wire N__9732;
    wire N__9729;
    wire N__9728;
    wire N__9725;
    wire N__9724;
    wire N__9721;
    wire N__9720;
    wire N__9717;
    wire N__9714;
    wire N__9711;
    wire N__9708;
    wire N__9699;
    wire N__9696;
    wire N__9693;
    wire N__9690;
    wire N__9687;
    wire N__9684;
    wire N__9681;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9669;
    wire N__9668;
    wire N__9667;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9645;
    wire N__9642;
    wire N__9639;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9621;
    wire N__9620;
    wire N__9619;
    wire N__9618;
    wire N__9617;
    wire N__9614;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9606;
    wire N__9605;
    wire N__9602;
    wire N__9601;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9593;
    wire N__9592;
    wire N__9591;
    wire N__9588;
    wire N__9583;
    wire N__9578;
    wire N__9577;
    wire N__9574;
    wire N__9569;
    wire N__9564;
    wire N__9557;
    wire N__9550;
    wire N__9547;
    wire N__9534;
    wire N__9533;
    wire N__9530;
    wire N__9529;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9501;
    wire N__9498;
    wire N__9495;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9483;
    wire N__9480;
    wire N__9477;
    wire N__9474;
    wire N__9471;
    wire N__9468;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9455;
    wire N__9454;
    wire N__9453;
    wire N__9452;
    wire N__9451;
    wire N__9450;
    wire N__9449;
    wire N__9448;
    wire N__9447;
    wire N__9446;
    wire N__9443;
    wire N__9442;
    wire N__9441;
    wire N__9440;
    wire N__9439;
    wire N__9438;
    wire N__9425;
    wire N__9420;
    wire N__9419;
    wire N__9418;
    wire N__9417;
    wire N__9414;
    wire N__9411;
    wire N__9410;
    wire N__9409;
    wire N__9408;
    wire N__9407;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9391;
    wire N__9386;
    wire N__9381;
    wire N__9378;
    wire N__9375;
    wire N__9372;
    wire N__9369;
    wire N__9366;
    wire N__9363;
    wire N__9360;
    wire N__9357;
    wire N__9356;
    wire N__9345;
    wire N__9344;
    wire N__9339;
    wire N__9336;
    wire N__9333;
    wire N__9330;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9303;
    wire N__9288;
    wire N__9285;
    wire N__9282;
    wire N__9279;
    wire N__9276;
    wire N__9273;
    wire N__9270;
    wire N__9267;
    wire N__9264;
    wire N__9261;
    wire N__9258;
    wire N__9255;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9236;
    wire N__9235;
    wire N__9234;
    wire N__9229;
    wire N__9228;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9210;
    wire N__9209;
    wire N__9206;
    wire N__9201;
    wire N__9200;
    wire N__9199;
    wire N__9198;
    wire N__9197;
    wire N__9196;
    wire N__9195;
    wire N__9194;
    wire N__9193;
    wire N__9192;
    wire N__9189;
    wire N__9182;
    wire N__9181;
    wire N__9174;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9147;
    wire N__9146;
    wire N__9145;
    wire N__9144;
    wire N__9143;
    wire N__9140;
    wire N__9139;
    wire N__9136;
    wire N__9133;
    wire N__9130;
    wire N__9127;
    wire N__9122;
    wire N__9119;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9101;
    wire N__9098;
    wire N__9097;
    wire N__9096;
    wire N__9093;
    wire N__9090;
    wire N__9087;
    wire N__9084;
    wire N__9081;
    wire N__9078;
    wire N__9071;
    wire N__9068;
    wire N__9063;
    wire N__9060;
    wire N__9057;
    wire N__9056;
    wire N__9055;
    wire N__9052;
    wire N__9051;
    wire N__9048;
    wire N__9047;
    wire N__9046;
    wire N__9045;
    wire N__9044;
    wire N__9043;
    wire N__9040;
    wire N__9039;
    wire N__9038;
    wire N__9037;
    wire N__9036;
    wire N__9035;
    wire N__9034;
    wire N__9029;
    wire N__9026;
    wire N__9025;
    wire N__9018;
    wire N__9013;
    wire N__9012;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9004;
    wire N__9003;
    wire N__8996;
    wire N__8991;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8970;
    wire N__8967;
    wire N__8964;
    wire N__8959;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8940;
    wire N__8937;
    wire N__8936;
    wire N__8935;
    wire N__8934;
    wire N__8931;
    wire N__8922;
    wire N__8919;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8901;
    wire N__8896;
    wire N__8883;
    wire N__8880;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8862;
    wire N__8859;
    wire N__8856;
    wire N__8853;
    wire N__8850;
    wire N__8849;
    wire N__8848;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8838;
    wire N__8835;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8819;
    wire N__8814;
    wire N__8813;
    wire N__8812;
    wire N__8807;
    wire N__8804;
    wire N__8803;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8787;
    wire N__8784;
    wire N__8781;
    wire N__8780;
    wire N__8779;
    wire N__8778;
    wire N__8775;
    wire N__8772;
    wire N__8767;
    wire N__8766;
    wire N__8763;
    wire N__8758;
    wire N__8755;
    wire N__8752;
    wire N__8749;
    wire N__8746;
    wire N__8745;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8724;
    wire N__8723;
    wire N__8722;
    wire N__8721;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8709;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8697;
    wire N__8694;
    wire N__8691;
    wire N__8686;
    wire N__8683;
    wire N__8680;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8663;
    wire N__8660;
    wire N__8659;
    wire N__8656;
    wire N__8653;
    wire N__8650;
    wire N__8643;
    wire N__8640;
    wire N__8637;
    wire N__8634;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8622;
    wire N__8619;
    wire N__8616;
    wire N__8615;
    wire N__8614;
    wire N__8611;
    wire N__8608;
    wire N__8605;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8587;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8562;
    wire N__8561;
    wire N__8560;
    wire N__8557;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8539;
    wire N__8536;
    wire N__8533;
    wire N__8530;
    wire N__8527;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8515;
    wire N__8514;
    wire N__8511;
    wire N__8506;
    wire N__8503;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8460;
    wire N__8457;
    wire N__8454;
    wire N__8451;
    wire N__8448;
    wire N__8447;
    wire N__8446;
    wire N__8443;
    wire N__8440;
    wire N__8437;
    wire N__8430;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8418;
    wire N__8415;
    wire N__8412;
    wire N__8409;
    wire N__8406;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8390;
    wire N__8389;
    wire N__8388;
    wire N__8385;
    wire N__8382;
    wire N__8379;
    wire N__8378;
    wire N__8377;
    wire N__8376;
    wire N__8375;
    wire N__8374;
    wire N__8373;
    wire N__8370;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8356;
    wire N__8351;
    wire N__8346;
    wire N__8343;
    wire N__8340;
    wire N__8337;
    wire N__8322;
    wire N__8319;
    wire N__8316;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8304;
    wire N__8301;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8293;
    wire N__8292;
    wire N__8291;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8265;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8241;
    wire N__8238;
    wire N__8235;
    wire N__8232;
    wire N__8229;
    wire N__8226;
    wire N__8225;
    wire N__8222;
    wire N__8219;
    wire N__8214;
    wire N__8211;
    wire N__8208;
    wire N__8205;
    wire N__8202;
    wire N__8199;
    wire N__8196;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8171;
    wire N__8166;
    wire N__8163;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8153;
    wire N__8148;
    wire N__8145;
    wire N__8142;
    wire N__8139;
    wire N__8136;
    wire N__8133;
    wire N__8130;
    wire N__8127;
    wire N__8124;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8099;
    wire N__8094;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8082;
    wire N__8079;
    wire N__8076;
    wire N__8073;
    wire N__8070;
    wire N__8067;
    wire N__8064;
    wire N__8061;
    wire N__8058;
    wire N__8055;
    wire N__8052;
    wire N__8049;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8037;
    wire N__8034;
    wire N__8031;
    wire N__8028;
    wire N__8025;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8013;
    wire N__8012;
    wire N__8011;
    wire N__8010;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7997;
    wire N__7996;
    wire N__7991;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7971;
    wire N__7968;
    wire N__7965;
    wire N__7962;
    wire N__7959;
    wire N__7956;
    wire N__7953;
    wire N__7950;
    wire N__7949;
    wire N__7948;
    wire N__7945;
    wire N__7942;
    wire N__7939;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7917;
    wire N__7914;
    wire N__7911;
    wire N__7910;
    wire N__7909;
    wire N__7906;
    wire N__7905;
    wire N__7904;
    wire N__7903;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7887;
    wire N__7884;
    wire N__7875;
    wire N__7872;
    wire N__7869;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7861;
    wire N__7858;
    wire N__7855;
    wire N__7852;
    wire N__7849;
    wire N__7846;
    wire N__7843;
    wire N__7840;
    wire N__7837;
    wire N__7834;
    wire N__7831;
    wire N__7828;
    wire N__7825;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7815;
    wire N__7812;
    wire N__7807;
    wire N__7804;
    wire N__7797;
    wire N__7796;
    wire N__7793;
    wire N__7790;
    wire N__7787;
    wire N__7784;
    wire N__7781;
    wire N__7778;
    wire N__7775;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7761;
    wire N__7758;
    wire N__7755;
    wire N__7754;
    wire N__7753;
    wire N__7750;
    wire N__7747;
    wire N__7746;
    wire N__7745;
    wire N__7744;
    wire N__7743;
    wire N__7742;
    wire N__7741;
    wire N__7740;
    wire N__7739;
    wire N__7738;
    wire N__7737;
    wire N__7734;
    wire N__7731;
    wire N__7730;
    wire N__7727;
    wire N__7720;
    wire N__7719;
    wire N__7714;
    wire N__7711;
    wire N__7710;
    wire N__7709;
    wire N__7708;
    wire N__7707;
    wire N__7702;
    wire N__7699;
    wire N__7698;
    wire N__7697;
    wire N__7696;
    wire N__7695;
    wire N__7694;
    wire N__7693;
    wire N__7692;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7674;
    wire N__7671;
    wire N__7666;
    wire N__7661;
    wire N__7656;
    wire N__7653;
    wire N__7648;
    wire N__7645;
    wire N__7640;
    wire N__7633;
    wire N__7630;
    wire N__7599;
    wire N__7598;
    wire N__7597;
    wire N__7596;
    wire N__7595;
    wire N__7594;
    wire N__7593;
    wire N__7592;
    wire N__7591;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7583;
    wire N__7582;
    wire N__7581;
    wire N__7580;
    wire N__7579;
    wire N__7578;
    wire N__7575;
    wire N__7572;
    wire N__7569;
    wire N__7562;
    wire N__7557;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7549;
    wire N__7548;
    wire N__7547;
    wire N__7546;
    wire N__7545;
    wire N__7542;
    wire N__7541;
    wire N__7540;
    wire N__7537;
    wire N__7534;
    wire N__7527;
    wire N__7524;
    wire N__7517;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7505;
    wire N__7500;
    wire N__7495;
    wire N__7490;
    wire N__7483;
    wire N__7478;
    wire N__7471;
    wire N__7452;
    wire N__7451;
    wire N__7450;
    wire N__7447;
    wire N__7444;
    wire N__7443;
    wire N__7440;
    wire N__7439;
    wire N__7438;
    wire N__7435;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7425;
    wire N__7420;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7397;
    wire N__7394;
    wire N__7391;
    wire N__7380;
    wire N__7379;
    wire N__7378;
    wire N__7375;
    wire N__7372;
    wire N__7371;
    wire N__7368;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7341;
    wire N__7338;
    wire N__7335;
    wire N__7332;
    wire N__7329;
    wire N__7326;
    wire N__7323;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7298;
    wire N__7295;
    wire N__7290;
    wire N__7287;
    wire N__7284;
    wire N__7281;
    wire N__7278;
    wire N__7277;
    wire N__7276;
    wire N__7271;
    wire N__7270;
    wire N__7267;
    wire N__7264;
    wire N__7261;
    wire N__7254;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7242;
    wire N__7241;
    wire N__7238;
    wire N__7237;
    wire N__7236;
    wire N__7233;
    wire N__7230;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7216;
    wire N__7215;
    wire N__7212;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7194;
    wire N__7191;
    wire N__7188;
    wire N__7187;
    wire N__7184;
    wire N__7183;
    wire N__7182;
    wire N__7179;
    wire N__7176;
    wire N__7171;
    wire N__7164;
    wire N__7161;
    wire N__7158;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7146;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7134;
    wire N__7131;
    wire N__7128;
    wire N__7125;
    wire N__7122;
    wire N__7119;
    wire N__7116;
    wire N__7113;
    wire N__7110;
    wire N__7107;
    wire N__7104;
    wire N__7101;
    wire N__7098;
    wire N__7095;
    wire N__7092;
    wire N__7089;
    wire N__7086;
    wire N__7083;
    wire N__7080;
    wire N__7077;
    wire N__7074;
    wire N__7073;
    wire N__7070;
    wire N__7067;
    wire N__7064;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7047;
    wire N__7044;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7029;
    wire N__7026;
    wire N__7023;
    wire N__7020;
    wire N__7017;
    wire N__7014;
    wire N__7011;
    wire N__7008;
    wire N__7007;
    wire N__7006;
    wire N__7005;
    wire N__7004;
    wire N__7003;
    wire N__7002;
    wire N__7001;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6987;
    wire N__6984;
    wire N__6977;
    wire N__6974;
    wire N__6963;
    wire N__6960;
    wire N__6957;
    wire N__6954;
    wire N__6951;
    wire N__6948;
    wire N__6945;
    wire N__6942;
    wire N__6939;
    wire N__6936;
    wire N__6933;
    wire N__6930;
    wire N__6927;
    wire N__6924;
    wire N__6921;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6900;
    wire N__6899;
    wire N__6898;
    wire N__6895;
    wire N__6894;
    wire N__6893;
    wire N__6892;
    wire N__6889;
    wire N__6886;
    wire N__6883;
    wire N__6880;
    wire N__6879;
    wire N__6870;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6846;
    wire N__6843;
    wire N__6840;
    wire N__6837;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6819;
    wire N__6816;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6804;
    wire N__6803;
    wire N__6800;
    wire N__6797;
    wire N__6792;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6777;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6765;
    wire N__6762;
    wire N__6759;
    wire N__6756;
    wire N__6753;
    wire N__6750;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6732;
    wire N__6729;
    wire N__6726;
    wire N__6723;
    wire N__6720;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6710;
    wire N__6707;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6684;
    wire N__6681;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6663;
    wire N__6660;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6648;
    wire N__6645;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6633;
    wire N__6630;
    wire N__6627;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6611;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6594;
    wire N__6593;
    wire N__6588;
    wire N__6585;
    wire N__6582;
    wire N__6579;
    wire N__6576;
    wire N__6573;
    wire N__6572;
    wire N__6571;
    wire N__6568;
    wire N__6563;
    wire N__6558;
    wire N__6557;
    wire N__6554;
    wire N__6553;
    wire N__6548;
    wire N__6545;
    wire N__6540;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6528;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6516;
    wire N__6515;
    wire N__6514;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6502;
    wire N__6495;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6483;
    wire N__6480;
    wire N__6477;
    wire N__6474;
    wire N__6471;
    wire N__6468;
    wire N__6465;
    wire N__6462;
    wire N__6459;
    wire N__6456;
    wire N__6453;
    wire N__6450;
    wire N__6449;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6441;
    wire N__6438;
    wire N__6435;
    wire N__6432;
    wire N__6429;
    wire N__6420;
    wire N__6419;
    wire N__6418;
    wire N__6415;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6405;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6390;
    wire N__6389;
    wire N__6386;
    wire N__6385;
    wire N__6384;
    wire N__6383;
    wire N__6380;
    wire N__6379;
    wire N__6378;
    wire N__6377;
    wire N__6376;
    wire N__6375;
    wire N__6372;
    wire N__6369;
    wire N__6364;
    wire N__6359;
    wire N__6352;
    wire N__6349;
    wire N__6346;
    wire N__6343;
    wire N__6338;
    wire N__6333;
    wire N__6312;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6300;
    wire N__6297;
    wire N__6296;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6284;
    wire N__6279;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6255;
    wire N__6252;
    wire N__6249;
    wire N__6246;
    wire N__6243;
    wire N__6242;
    wire N__6241;
    wire N__6238;
    wire N__6233;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6216;
    wire N__6215;
    wire N__6212;
    wire N__6209;
    wire N__6204;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6186;
    wire N__6183;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6171;
    wire N__6168;
    wire N__6165;
    wire N__6162;
    wire N__6161;
    wire N__6158;
    wire N__6155;
    wire N__6154;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6137;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6122;
    wire N__6119;
    wire N__6114;
    wire N__6113;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6099;
    wire N__6096;
    wire N__6093;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6081;
    wire N__6080;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6067;
    wire N__6062;
    wire N__6059;
    wire N__6054;
    wire N__6051;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6038;
    wire N__6035;
    wire N__6032;
    wire N__6027;
    wire N__6024;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5987;
    wire N__5982;
    wire N__5979;
    wire N__5978;
    wire N__5975;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5943;
    wire N__5940;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5907;
    wire N__5904;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5871;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5829;
    wire N__5826;
    wire N__5823;
    wire N__5820;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5769;
    wire N__5766;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5754;
    wire N__5751;
    wire N__5748;
    wire N__5745;
    wire N__5742;
    wire N__5739;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5729;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5709;
    wire N__5706;
    wire N__5703;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5682;
    wire N__5679;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5667;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5640;
    wire N__5639;
    wire N__5638;
    wire N__5637;
    wire N__5636;
    wire N__5635;
    wire N__5634;
    wire N__5631;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5613;
    wire N__5606;
    wire N__5605;
    wire N__5604;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5596;
    wire N__5595;
    wire N__5594;
    wire N__5593;
    wire N__5592;
    wire N__5591;
    wire N__5588;
    wire N__5583;
    wire N__5578;
    wire N__5575;
    wire N__5566;
    wire N__5563;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5540;
    wire N__5537;
    wire N__5536;
    wire N__5535;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5520;
    wire N__5517;
    wire N__5508;
    wire N__5505;
    wire N__5502;
    wire N__5499;
    wire N__5498;
    wire N__5497;
    wire N__5494;
    wire N__5493;
    wire N__5490;
    wire N__5487;
    wire N__5482;
    wire N__5481;
    wire N__5474;
    wire N__5471;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5427;
    wire N__5424;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5409;
    wire N__5406;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5391;
    wire N__5388;
    wire N__5385;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5370;
    wire N__5367;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5352;
    wire N__5349;
    wire N__5346;
    wire N__5343;
    wire N__5340;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5325;
    wire N__5322;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5304;
    wire N__5301;
    wire N__5298;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5286;
    wire N__5283;
    wire N__5280;
    wire N__5279;
    wire N__5278;
    wire N__5277;
    wire N__5276;
    wire N__5273;
    wire N__5272;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5250;
    wire N__5247;
    wire N__5242;
    wire N__5239;
    wire N__5234;
    wire N__5233;
    wire N__5232;
    wire N__5231;
    wire N__5230;
    wire N__5229;
    wire N__5226;
    wire N__5225;
    wire N__5224;
    wire N__5219;
    wire N__5216;
    wire N__5209;
    wire N__5206;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5186;
    wire N__5169;
    wire N__5166;
    wire N__5163;
    wire N__5160;
    wire N__5159;
    wire N__5158;
    wire N__5157;
    wire N__5156;
    wire N__5155;
    wire N__5154;
    wire N__5153;
    wire N__5146;
    wire N__5141;
    wire N__5134;
    wire N__5127;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5115;
    wire N__5112;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5097;
    wire N__5094;
    wire N__5091;
    wire N__5090;
    wire N__5089;
    wire N__5084;
    wire N__5081;
    wire N__5076;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5064;
    wire N__5063;
    wire N__5062;
    wire N__5059;
    wire N__5054;
    wire N__5049;
    wire N__5046;
    wire N__5043;
    wire N__5042;
    wire N__5041;
    wire N__5040;
    wire N__5039;
    wire N__5038;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5017;
    wire N__5014;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4983;
    wire N__4980;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4911;
    wire N__4910;
    wire N__4909;
    wire N__4906;
    wire N__4903;
    wire N__4902;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4890;
    wire N__4881;
    wire N__4878;
    wire N__4875;
    wire N__4874;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4854;
    wire N__4845;
    wire N__4842;
    wire N__4839;
    wire N__4836;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4764;
    wire N__4761;
    wire N__4758;
    wire N__4755;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4743;
    wire N__4740;
    wire N__4737;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4727;
    wire N__4724;
    wire N__4723;
    wire N__4722;
    wire N__4719;
    wire N__4716;
    wire N__4711;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4695;
    wire N__4692;
    wire N__4691;
    wire N__4690;
    wire N__4687;
    wire N__4686;
    wire N__4683;
    wire N__4680;
    wire N__4677;
    wire N__4672;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4650;
    wire N__4647;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4607;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4593;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4575;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4562;
    wire N__4561;
    wire N__4560;
    wire N__4559;
    wire N__4558;
    wire N__4557;
    wire N__4556;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4494;
    wire N__4491;
    wire N__4488;
    wire N__4485;
    wire N__4482;
    wire N__4479;
    wire N__4478;
    wire N__4473;
    wire N__4470;
    wire N__4467;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4406;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire DBRn_c_i_0;
    wire CLK80_PLL_i_i;
    wire DBRn_c_i;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_5 ;
    wire \U712_CHIP_RAM.N_458_cascade_ ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_4 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a2_0_cascade_ ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1_cascade_ ;
    wire \U712_CHIP_RAM.N_442_cascade_ ;
    wire \U712_CHIP_RAM.CLK_EN_5_0 ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_7_13_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire DBRn_c;
    wire DBR_SYNCZ0Z_0;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_1_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_1_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_1_5_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_1_4 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_2_2_cascade_ ;
    wire \U712_CHIP_RAM.N_433 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_4_i_2_cascade_ ;
    wire \U712_CHIP_RAM.N_65 ;
    wire \U712_CHIP_RAM.N_173_cascade_ ;
    wire VBENn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_2_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_2_3 ;
    wire \U712_CHIP_RAM.N_301_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_0_1_cascade_ ;
    wire bfn_8_12_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.LATCH_CLK_6 ;
    wire \U712_CHIP_RAM.N_396_cascade_ ;
    wire LATCH_CLK_c;
    wire \U712_CHIP_RAM.N_315 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.N_336 ;
    wire \U712_CHIP_RAM.N_372 ;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.CMA_5_i_0_9 ;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_3_cascade_ ;
    wire \U712_CHIP_RAM.N_191_cascade_ ;
    wire \U712_CHIP_RAM.N_191_0 ;
    wire A_c_18;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_0_4 ;
    wire \U712_CHIP_RAM.N_191 ;
    wire \U712_CHIP_RAM.N_327 ;
    wire \U712_CHIP_RAM.N_300 ;
    wire \U712_CHIP_RAM.N_370 ;
    wire \U712_CHIP_RAM.N_301 ;
    wire \U712_CHIP_RAM.N_466_cascade_ ;
    wire \U712_CHIP_RAM.N_299_cascade_ ;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ;
    wire A_c_16;
    wire \U712_CHIP_RAM.N_399_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_0_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_310 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_385 ;
    wire \U712_CHIP_RAM.N_182 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_0 ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_382 ;
    wire \U712_CHIP_RAM.N_534 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_cascade_ ;
    wire \U712_REG_SM.N_411_cascade_ ;
    wire \U712_BYTE_ENABLE.N_446_cascade_ ;
    wire N_52_i;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire bfn_9_15_0_;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_1 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_2 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_3 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_4 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_5 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_6 ;
    wire \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ;
    wire CONSTANT_ONE_NET;
    wire CMA_c_5;
    wire A_c_11;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ;
    wire A_c_17;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ;
    wire A_c_14;
    wire \U712_CHIP_RAM.N_353 ;
    wire A_c_20;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.DBENn_7_0_0 ;
    wire DBDIR_c;
    wire \U712_CHIP_RAM.un1_CMA25_0_i ;
    wire A_c_12;
    wire A_c_5;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.N_471 ;
    wire A_c_3;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ;
    wire A_c_4;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ;
    wire A_c_6;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.N_429 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.N_319 ;
    wire \U712_CHIP_RAM.N_359 ;
    wire AWEn_c;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0_a2_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.N_419_cascade_ ;
    wire RAMSPACEn_c;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.N_299 ;
    wire \U712_CHIP_RAM.N_307 ;
    wire \U712_CHIP_RAM.N_434 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH5lto7_0 ;
    wire \U712_CHIP_RAM.REFRESH5lt7 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_REG_SM.N_322_cascade_ ;
    wire \U712_REG_SM.N_367_cascade_ ;
    wire \U712_REG_SM.N_408_cascade_ ;
    wire \U712_REG_SM.N_367 ;
    wire \U712_REG_SM.N_410 ;
    wire \U712_REG_SM.WRITE_CYCLEZ0 ;
    wire \U712_REG_SM.REGENn_e_1 ;
    wire REGENn_c;
    wire \U712_REG_SM.N_322 ;
    wire \U712_REG_SM.N_131 ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_1 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_6 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_2 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_0 ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLE_5_i_a2_4_cascade_ ;
    wire \U712_CHIP_RAM.N_456 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_5 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_4 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_3 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_7 ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLE_5_i_a2_5 ;
    wire DMA_LATCH_EN_c;
    wire CMA_c_10;
    wire A_c_9;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_ ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CMA_c_2;
    wire A_c_7;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ;
    wire A_c_2;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ;
    wire A_c_8;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ;
    wire CMA_c_4;
    wire CMA_c_3;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_466 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0 ;
    wire REGSPACEn_c;
    wire TSn_c;
    wire \U712_REG_SM.N_401_cascade_ ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_0 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_REG_SM.N_324_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_2 ;
    wire \U712_REG_SM.STATE_COUNTc_0_0 ;
    wire \U712_BYTE_ENABLE.N_424 ;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0 ;
    wire N_170_i;
    wire \U712_REG_SM.N_325_cascade_ ;
    wire \U712_REG_SM.N_302 ;
    wire \U712_REG_SM.N_302_cascade_ ;
    wire REG_CYCLEm;
    wire N_160_i;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.N_404 ;
    wire TACK_OUTn;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ1Z_2 ;
    wire ASn_c;
    wire \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0 ;
    wire RASn_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire \U712_CHIP_RAM.N_309_cascade_ ;
    wire \U712_CHIP_RAM.N_309 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1_cascade_ ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.un1_CMA25_0_i_0 ;
    wire A_c_15;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire A_c_10;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire A_c_13;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_3 ;
    wire CLK40_PLL_i_i;
    wire TACK_EN;
    wire C3_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ;
    wire \U712_REG_SM.START_RSTZ0 ;
    wire \U712_BYTE_ENABLE.N_443_cascade_ ;
    wire N_54_i;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_1 ;
    wire \U712_CYCLE_TERM.N_452_cascade_ ;
    wire CLK40_PLL_i;
    wire CPU_CYCLEm;
    wire \U712_BYTE_ENABLE.N_421_cascade_ ;
    wire N_168_i;
    wire \U712_CYCLE_TERM.N_326 ;
    wire REG_TACK;
    wire CPU_TACKm;
    wire DBENn_c;
    wire DMA_CYCLEm;
    wire \U712_BYTE_ENABLE.N_425 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_REG_SM.N_402 ;
    wire LDSn_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.un1_REGENn_0_sqmuxa_0 ;
    wire UDSn_c;
    wire RESETn_c_i;
    wire N_166;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ;
    wire \U712_BYTE_ENABLE.N_298_i ;
    wire \U712_REG_SM.N_459 ;
    wire N_390_i;
    wire N_389_i;
    wire A_c_0;
    wire A_c_1;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire N_189;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_6;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire WEn_c;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire DRA_c_7;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire DRA_c_3;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ;
    wire AGNUS_REV_c;
    wire DRA_c_1;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire RAS1n_c;
    wire RAS0n_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire RESETn_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_2 ;
    wire CLK80_PLL;
    wire DMA_WRITE_CYCLE;
    wire RnW_c;
    wire CASUn_c;
    wire CASLn_c;
    wire DRDDIR_c;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__4347),
            .RESETB(N__5871),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__12817),
            .DIN(N__12816),
            .DOUT(N__12815),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__12817),
            .PADOUT(N__12816),
            .PADIN(N__12815),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8787),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__12808),
            .DIN(N__12807),
            .DOUT(N__12806),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__12808),
            .PADOUT(N__12807),
            .PADIN(N__12806),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__12799),
            .DIN(N__12798),
            .DOUT(N__12797),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__12799),
            .PADOUT(N__12798),
            .PADIN(N__12797),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9288),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__12790),
            .DIN(N__12789),
            .DOUT(N__12788),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__12790),
            .PADOUT(N__12789),
            .PADIN(N__12788),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11808),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__12781),
            .DIN(N__12780),
            .DOUT(N__12779),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__12781),
            .PADOUT(N__12780),
            .PADIN(N__12779),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__12772),
            .DIN(N__12771),
            .DOUT(N__12770),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__12772),
            .PADOUT(N__12771),
            .PADIN(N__12770),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__12763),
            .DIN(N__12762),
            .DOUT(N__12761),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__12763),
            .PADOUT(N__12762),
            .PADIN(N__12761),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__12754),
            .DIN(N__12753),
            .DOUT(N__12752),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__12754),
            .PADOUT(N__12753),
            .PADIN(N__12752),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__12745),
            .DIN(N__12744),
            .DOUT(N__12743),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__12745),
            .PADOUT(N__12744),
            .PADIN(N__12743),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__12736),
            .DIN(N__12735),
            .DOUT(N__12734),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__12736),
            .PADOUT(N__12735),
            .PADIN(N__12734),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__12727),
            .DIN(N__12726),
            .DOUT(N__12725),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__12727),
            .PADOUT(N__12726),
            .PADIN(N__12725),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__12718),
            .DIN(N__12717),
            .DOUT(N__12716),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__12718),
            .PADOUT(N__12717),
            .PADIN(N__12716),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6840),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__12709),
            .DIN(N__12708),
            .DOUT(N__12707),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__12709),
            .PADOUT(N__12708),
            .PADIN(N__12707),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9903),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__12700),
            .DIN(N__12699),
            .DOUT(N__12698),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__12700),
            .PADOUT(N__12699),
            .PADIN(N__12698),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__12691),
            .DIN(N__12690),
            .DOUT(N__12689),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__12691),
            .PADOUT(N__12690),
            .PADIN(N__12689),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__12682),
            .DIN(N__12681),
            .DOUT(N__12680),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__12682),
            .PADOUT(N__12681),
            .PADIN(N__12680),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__12673),
            .DIN(N__12672),
            .DOUT(N__12671),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__12673),
            .PADOUT(N__12672),
            .PADIN(N__12671),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4584),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__12664),
            .DIN(N__12663),
            .DOUT(N__12662),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__12664),
            .PADOUT(N__12663),
            .PADIN(N__12662),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__12655),
            .DIN(N__12654),
            .DOUT(N__12653),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__12655),
            .PADOUT(N__12654),
            .PADIN(N__12653),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__12646),
            .DIN(N__12645),
            .DOUT(N__12644),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__12646),
            .PADOUT(N__12645),
            .PADIN(N__12644),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6678),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__12637),
            .DIN(N__12636),
            .DOUT(N__12635),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__12637),
            .PADOUT(N__12636),
            .PADIN(N__12635),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__12628),
            .DIN(N__12627),
            .DOUT(N__12626),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__12628),
            .PADOUT(N__12627),
            .PADIN(N__12626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10050),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__12619),
            .DIN(N__12618),
            .DOUT(N__12617),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__12619),
            .PADOUT(N__12618),
            .PADIN(N__12617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__12610),
            .DIN(N__12609),
            .DOUT(N__12608),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__12610),
            .PADOUT(N__12609),
            .PADIN(N__12608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10326),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__12601),
            .DIN(N__12600),
            .DOUT(N__12599),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__12601),
            .PADOUT(N__12600),
            .PADIN(N__12599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8561),
            .DIN0(),
            .DOUT0(N__7869),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__12592),
            .DIN(N__12591),
            .DOUT(N__12590),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__12592),
            .PADOUT(N__12591),
            .PADIN(N__12590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__12583),
            .DIN(N__12582),
            .DOUT(N__12581),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__12583),
            .PADOUT(N__12582),
            .PADIN(N__12581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__12574),
            .DIN(N__12573),
            .DOUT(N__12572),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__12574),
            .PADOUT(N__12573),
            .PADIN(N__12572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__12565),
            .DIN(N__12564),
            .DOUT(N__12563),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__12565),
            .PADOUT(N__12564),
            .PADIN(N__12563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__12556),
            .DIN(N__12555),
            .DOUT(N__12554),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__12556),
            .PADOUT(N__12555),
            .PADIN(N__12554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__12547),
            .DIN(N__12546),
            .DOUT(N__12545),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__12547),
            .PADOUT(N__12546),
            .PADIN(N__12545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6759),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__12538),
            .DIN(N__12537),
            .DOUT(N__12536),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__12538),
            .PADOUT(N__12537),
            .PADIN(N__12536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__12529),
            .DIN(N__12528),
            .DOUT(N__12527),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__12529),
            .PADOUT(N__12528),
            .PADIN(N__12527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__12520),
            .DIN(N__12519),
            .DOUT(N__12518),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__12520),
            .PADOUT(N__12519),
            .PADIN(N__12518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__12511),
            .DIN(N__12510),
            .DOUT(N__12509),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__12511),
            .PADOUT(N__12510),
            .PADIN(N__12509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__12502),
            .DIN(N__12501),
            .DOUT(N__12500),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__12502),
            .PADOUT(N__12501),
            .PADIN(N__12500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__12493),
            .DIN(N__12492),
            .DOUT(N__12491),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__12493),
            .PADOUT(N__12492),
            .PADIN(N__12491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8055),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__12484),
            .DIN(N__12483),
            .DOUT(N__12482),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__12484),
            .PADOUT(N__12483),
            .PADIN(N__12482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__12475),
            .DIN(N__12474),
            .DOUT(N__12473),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__12475),
            .PADOUT(N__12474),
            .PADIN(N__12473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__12466),
            .DIN(N__12465),
            .DOUT(N__12464),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__12466),
            .PADOUT(N__12465),
            .PADIN(N__12464),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8091),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_0_iopad (
            .OE(N__12457),
            .DIN(N__12456),
            .DOUT(N__12455),
            .PACKAGEPIN(DA[0]));
    defparam DA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_0_preio (
            .PADOEN(N__12457),
            .PADOUT(N__12456),
            .PADIN(N__12455),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6720),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__12448),
            .DIN(N__12447),
            .DOUT(N__12446),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__12448),
            .PADOUT(N__12447),
            .PADIN(N__12446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__12439),
            .DIN(N__12438),
            .DOUT(N__12437),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__12439),
            .PADOUT(N__12438),
            .PADIN(N__12437),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6741),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__12430),
            .DIN(N__12429),
            .DOUT(N__12428),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__12430),
            .PADOUT(N__12429),
            .PADIN(N__12428),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6963),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__12421),
            .DIN(N__12420),
            .DOUT(N__12419),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__12421),
            .PADOUT(N__12420),
            .PADIN(N__12419),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6627),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__12412),
            .DIN(N__12411),
            .DOUT(N__12410),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__12412),
            .PADOUT(N__12411),
            .PADIN(N__12410),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__12403),
            .DIN(N__12402),
            .DOUT(N__12401),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__12403),
            .PADOUT(N__12402),
            .PADIN(N__12401),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8415),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__12394),
            .DIN(N__12393),
            .DOUT(N__12392),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__12394),
            .PADOUT(N__12393),
            .PADIN(N__12392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8562),
            .DIN0(),
            .DOUT0(N__7868),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__12385),
            .DIN(N__12384),
            .DOUT(N__12383),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__12385),
            .PADOUT(N__12384),
            .PADIN(N__12383),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9996),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__12376),
            .DIN(N__12375),
            .DOUT(N__12374),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__12376),
            .PADOUT(N__12375),
            .PADIN(N__12374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6054),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__12367),
            .DIN(N__12366),
            .DOUT(N__12365),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__12367),
            .PADOUT(N__12366),
            .PADIN(N__12365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7134),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__12358),
            .DIN(N__12357),
            .DOUT(N__12356),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__12358),
            .PADOUT(N__12357),
            .PADIN(N__12356),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__12349),
            .DIN(N__12348),
            .DOUT(N__12347),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__12349),
            .PADOUT(N__12348),
            .PADIN(N__12347),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_2_iopad (
            .OE(N__12340),
            .DIN(N__12339),
            .DOUT(N__12338),
            .PACKAGEPIN(DA[2]));
    defparam DA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_2_preio (
            .PADOEN(N__12340),
            .PADOUT(N__12339),
            .PADIN(N__12338),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5814),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__12331),
            .DIN(N__12330),
            .DOUT(N__12329),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__12331),
            .PADOUT(N__12330),
            .PADIN(N__12329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__12322),
            .DIN(N__12321),
            .DOUT(N__12320),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__12322),
            .PADOUT(N__12321),
            .PADIN(N__12320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__12313),
            .DIN(N__12312),
            .DOUT(N__12311),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__12313),
            .PADOUT(N__12312),
            .PADIN(N__12311),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8313),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__12304),
            .DIN(N__12303),
            .DOUT(N__12302),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__12304),
            .PADOUT(N__12303),
            .PADIN(N__12302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9888),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__12295),
            .DIN(N__12294),
            .DOUT(N__12293),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__12295),
            .PADOUT(N__12294),
            .PADIN(N__12293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__12286),
            .DIN(N__12285),
            .DOUT(N__12284),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__12286),
            .PADOUT(N__12285),
            .PADIN(N__12284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8880),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__12277),
            .DIN(N__12276),
            .DOUT(N__12275),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__12277),
            .PADOUT(N__12276),
            .PADIN(N__12275),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8560),
            .DIN0(),
            .DOUT0(N__7861),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__12268),
            .DIN(N__12267),
            .DOUT(N__12266),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__12268),
            .PADOUT(N__12267),
            .PADIN(N__12266),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7104),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__12259),
            .DIN(N__12258),
            .DOUT(N__12257),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__12259),
            .PADOUT(N__12258),
            .PADIN(N__12257),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__12250),
            .DIN(N__12249),
            .DOUT(N__12248),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__12250),
            .PADOUT(N__12249),
            .PADIN(N__12248),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__12241),
            .DIN(N__12240),
            .DOUT(N__12239),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__12241),
            .PADOUT(N__12240),
            .PADIN(N__12239),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4764),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__12232),
            .DIN(N__12231),
            .DOUT(N__12230),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__12232),
            .PADOUT(N__12231),
            .PADIN(N__12230),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__12223),
            .DIN(N__12222),
            .DOUT(N__12221),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__12223),
            .PADOUT(N__12222),
            .PADIN(N__12221),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_1_iopad (
            .OE(N__12214),
            .DIN(N__12213),
            .DOUT(N__12212),
            .PACKAGEPIN(DA[1]));
    defparam DA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_1_preio (
            .PADOEN(N__12214),
            .PADOUT(N__12213),
            .PADIN(N__12212),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8205),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__12205),
            .DIN(N__12204),
            .DOUT(N__12203),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__12205),
            .PADOUT(N__12204),
            .PADIN(N__12203),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__12196),
            .DIN(N__12195),
            .DOUT(N__12194),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__12196),
            .PADOUT(N__12195),
            .PADIN(N__12194),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__12187),
            .DIN(N__12186),
            .DOUT(N__12185),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__12187),
            .PADOUT(N__12186),
            .PADIN(N__12185),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5838),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__12178),
            .DIN(N__12177),
            .DOUT(N__12176),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__12178),
            .PADOUT(N__12177),
            .PADIN(N__12176),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9510),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__12169),
            .DIN(N__12168),
            .DOUT(N__12167),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__12169),
            .PADOUT(N__12168),
            .PADIN(N__12167),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9468),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__12160),
            .DIN(N__12159),
            .DOUT(N__12158),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__12160),
            .PADOUT(N__12159),
            .PADIN(N__12158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4395),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__12151),
            .DIN(N__12150),
            .DOUT(N__12149),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__12151),
            .PADOUT(N__12150),
            .PADIN(N__12149),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__12142),
            .DIN(N__12141),
            .DOUT(N__12140),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__12142),
            .PADOUT(N__12141),
            .PADIN(N__12140),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__12133),
            .DIN(N__12132),
            .DOUT(N__12131),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__12133),
            .PADOUT(N__12132),
            .PADIN(N__12131),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6915),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__12124),
            .DIN(N__12123),
            .DOUT(N__12122),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__12124),
            .PADOUT(N__12123),
            .PADIN(N__12122),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__12115),
            .DIN(N__12114),
            .DOUT(N__12113),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__12115),
            .PADOUT(N__12114),
            .PADIN(N__12113),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__12106),
            .DIN(N__12105),
            .DOUT(N__12104),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__12106),
            .PADOUT(N__12105),
            .PADIN(N__12104),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4656),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__12097),
            .DIN(N__12096),
            .DOUT(N__12095),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__12097),
            .PADOUT(N__12096),
            .PADIN(N__12095),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9645),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__12088),
            .DIN(N__12087),
            .DOUT(N__12086),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__12088),
            .PADOUT(N__12087),
            .PADIN(N__12086),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8616),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__12079),
            .DIN(N__12078),
            .DOUT(N__12077),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__12079),
            .PADOUT(N__12078),
            .PADIN(N__12077),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__12070),
            .DIN(N__12069),
            .DOUT(N__12068),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__12070),
            .PADOUT(N__12069),
            .PADIN(N__12068),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8615),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__12061),
            .DIN(N__12060),
            .DOUT(N__12059),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__12061),
            .PADOUT(N__12060),
            .PADIN(N__12059),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4362),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__12052),
            .DIN(N__12051),
            .DOUT(N__12050),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__12052),
            .PADOUT(N__12051),
            .PADIN(N__12050),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6939),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__12043),
            .DIN(N__12042),
            .DOUT(N__12041),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__12043),
            .PADOUT(N__12042),
            .PADIN(N__12041),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__12034),
            .DIN(N__12033),
            .DOUT(N__12032),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__12034),
            .PADOUT(N__12033),
            .PADIN(N__12032),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__12025),
            .DIN(N__12024),
            .DOUT(N__12023),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__12025),
            .PADOUT(N__12024),
            .PADIN(N__12023),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__12016),
            .DIN(N__12015),
            .DOUT(N__12014),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__12016),
            .PADOUT(N__12015),
            .PADIN(N__12014),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__12007),
            .DIN(N__12006),
            .DOUT(N__12005),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__12007),
            .PADOUT(N__12006),
            .PADIN(N__12005),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8614),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11998),
            .DIN(N__11997),
            .DOUT(N__11996),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11998),
            .PADOUT(N__11997),
            .PADIN(N__11996),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7932),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11989),
            .DIN(N__11988),
            .DOUT(N__11987),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11989),
            .PADOUT(N__11988),
            .PADIN(N__11987),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5457),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11980),
            .DIN(N__11979),
            .DOUT(N__11978),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11980),
            .PADOUT(N__11979),
            .PADIN(N__11978),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4944),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11971),
            .DIN(N__11970),
            .DOUT(N__11969),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11971),
            .PADOUT(N__11970),
            .PADIN(N__11969),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2915 (
            .O(N__11952),
            .I(N__11947));
    InMux I__2914 (
            .O(N__11951),
            .I(N__11944));
    InMux I__2913 (
            .O(N__11950),
            .I(N__11941));
    LocalMux I__2912 (
            .O(N__11947),
            .I(N__11938));
    LocalMux I__2911 (
            .O(N__11944),
            .I(N__11933));
    LocalMux I__2910 (
            .O(N__11941),
            .I(N__11933));
    Span4Mux_v I__2909 (
            .O(N__11938),
            .I(N__11928));
    Span4Mux_v I__2908 (
            .O(N__11933),
            .I(N__11928));
    Span4Mux_v I__2907 (
            .O(N__11928),
            .I(N__11924));
    InMux I__2906 (
            .O(N__11927),
            .I(N__11920));
    Span4Mux_h I__2905 (
            .O(N__11924),
            .I(N__11916));
    CascadeMux I__2904 (
            .O(N__11923),
            .I(N__11913));
    LocalMux I__2903 (
            .O(N__11920),
            .I(N__11910));
    InMux I__2902 (
            .O(N__11919),
            .I(N__11907));
    Span4Mux_h I__2901 (
            .O(N__11916),
            .I(N__11904));
    InMux I__2900 (
            .O(N__11913),
            .I(N__11901));
    Sp12to4 I__2899 (
            .O(N__11910),
            .I(N__11896));
    LocalMux I__2898 (
            .O(N__11907),
            .I(N__11896));
    Span4Mux_h I__2897 (
            .O(N__11904),
            .I(N__11891));
    LocalMux I__2896 (
            .O(N__11901),
            .I(N__11891));
    Span12Mux_v I__2895 (
            .O(N__11896),
            .I(N__11888));
    Span4Mux_h I__2894 (
            .O(N__11891),
            .I(N__11885));
    Span12Mux_h I__2893 (
            .O(N__11888),
            .I(N__11882));
    Span4Mux_v I__2892 (
            .O(N__11885),
            .I(N__11879));
    Odrv12 I__2891 (
            .O(N__11882),
            .I(CASUn_c));
    Odrv4 I__2890 (
            .O(N__11879),
            .I(CASUn_c));
    InMux I__2889 (
            .O(N__11874),
            .I(N__11869));
    InMux I__2888 (
            .O(N__11873),
            .I(N__11865));
    InMux I__2887 (
            .O(N__11872),
            .I(N__11862));
    LocalMux I__2886 (
            .O(N__11869),
            .I(N__11859));
    InMux I__2885 (
            .O(N__11868),
            .I(N__11856));
    LocalMux I__2884 (
            .O(N__11865),
            .I(N__11851));
    LocalMux I__2883 (
            .O(N__11862),
            .I(N__11851));
    Span4Mux_v I__2882 (
            .O(N__11859),
            .I(N__11845));
    LocalMux I__2881 (
            .O(N__11856),
            .I(N__11845));
    Span4Mux_h I__2880 (
            .O(N__11851),
            .I(N__11842));
    InMux I__2879 (
            .O(N__11850),
            .I(N__11839));
    Span4Mux_v I__2878 (
            .O(N__11845),
            .I(N__11836));
    Sp12to4 I__2877 (
            .O(N__11842),
            .I(N__11830));
    LocalMux I__2876 (
            .O(N__11839),
            .I(N__11830));
    Span4Mux_v I__2875 (
            .O(N__11836),
            .I(N__11827));
    InMux I__2874 (
            .O(N__11835),
            .I(N__11824));
    Span12Mux_v I__2873 (
            .O(N__11830),
            .I(N__11819));
    Sp12to4 I__2872 (
            .O(N__11827),
            .I(N__11819));
    LocalMux I__2871 (
            .O(N__11824),
            .I(N__11816));
    Span12Mux_h I__2870 (
            .O(N__11819),
            .I(N__11811));
    Span12Mux_v I__2869 (
            .O(N__11816),
            .I(N__11811));
    Odrv12 I__2868 (
            .O(N__11811),
            .I(CASLn_c));
    IoInMux I__2867 (
            .O(N__11808),
            .I(N__11805));
    LocalMux I__2866 (
            .O(N__11805),
            .I(N__11802));
    Span4Mux_s3_h I__2865 (
            .O(N__11802),
            .I(N__11799));
    Span4Mux_v I__2864 (
            .O(N__11799),
            .I(N__11796));
    Odrv4 I__2863 (
            .O(N__11796),
            .I(DRDDIR_c));
    InMux I__2862 (
            .O(N__11793),
            .I(N__11787));
    InMux I__2861 (
            .O(N__11792),
            .I(N__11787));
    LocalMux I__2860 (
            .O(N__11787),
            .I(N__11784));
    Span4Mux_h I__2859 (
            .O(N__11784),
            .I(N__11781));
    Odrv4 I__2858 (
            .O(N__11781),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__2857 (
            .O(N__11778),
            .I(N__11774));
    InMux I__2856 (
            .O(N__11777),
            .I(N__11771));
    LocalMux I__2855 (
            .O(N__11774),
            .I(N__11768));
    LocalMux I__2854 (
            .O(N__11771),
            .I(N__11763));
    Span4Mux_v I__2853 (
            .O(N__11768),
            .I(N__11760));
    InMux I__2852 (
            .O(N__11767),
            .I(N__11755));
    InMux I__2851 (
            .O(N__11766),
            .I(N__11755));
    Span4Mux_v I__2850 (
            .O(N__11763),
            .I(N__11752));
    Sp12to4 I__2849 (
            .O(N__11760),
            .I(N__11747));
    LocalMux I__2848 (
            .O(N__11755),
            .I(N__11747));
    Sp12to4 I__2847 (
            .O(N__11752),
            .I(N__11744));
    Span12Mux_h I__2846 (
            .O(N__11747),
            .I(N__11741));
    Span12Mux_h I__2845 (
            .O(N__11744),
            .I(N__11738));
    Odrv12 I__2844 (
            .O(N__11741),
            .I(DRA_c_7));
    Odrv12 I__2843 (
            .O(N__11738),
            .I(DRA_c_7));
    InMux I__2842 (
            .O(N__11733),
            .I(N__11727));
    InMux I__2841 (
            .O(N__11732),
            .I(N__11724));
    InMux I__2840 (
            .O(N__11731),
            .I(N__11721));
    InMux I__2839 (
            .O(N__11730),
            .I(N__11718));
    LocalMux I__2838 (
            .O(N__11727),
            .I(N__11715));
    LocalMux I__2837 (
            .O(N__11724),
            .I(N__11712));
    LocalMux I__2836 (
            .O(N__11721),
            .I(N__11707));
    LocalMux I__2835 (
            .O(N__11718),
            .I(N__11707));
    Span4Mux_v I__2834 (
            .O(N__11715),
            .I(N__11702));
    Span4Mux_v I__2833 (
            .O(N__11712),
            .I(N__11702));
    Span4Mux_v I__2832 (
            .O(N__11707),
            .I(N__11699));
    Span4Mux_h I__2831 (
            .O(N__11702),
            .I(N__11696));
    Span4Mux_h I__2830 (
            .O(N__11699),
            .I(N__11693));
    Sp12to4 I__2829 (
            .O(N__11696),
            .I(N__11688));
    Sp12to4 I__2828 (
            .O(N__11693),
            .I(N__11688));
    Odrv12 I__2827 (
            .O(N__11688),
            .I(DRA_c_8));
    InMux I__2826 (
            .O(N__11685),
            .I(N__11682));
    LocalMux I__2825 (
            .O(N__11682),
            .I(N__11679));
    Span4Mux_v I__2824 (
            .O(N__11679),
            .I(N__11676));
    Odrv4 I__2823 (
            .O(N__11676),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2822 (
            .O(N__11673),
            .I(N__11670));
    LocalMux I__2821 (
            .O(N__11670),
            .I(N__11664));
    InMux I__2820 (
            .O(N__11669),
            .I(N__11661));
    InMux I__2819 (
            .O(N__11668),
            .I(N__11658));
    InMux I__2818 (
            .O(N__11667),
            .I(N__11655));
    Span4Mux_h I__2817 (
            .O(N__11664),
            .I(N__11650));
    LocalMux I__2816 (
            .O(N__11661),
            .I(N__11650));
    LocalMux I__2815 (
            .O(N__11658),
            .I(N__11647));
    LocalMux I__2814 (
            .O(N__11655),
            .I(N__11642));
    Sp12to4 I__2813 (
            .O(N__11650),
            .I(N__11642));
    Span4Mux_h I__2812 (
            .O(N__11647),
            .I(N__11639));
    Span12Mux_v I__2811 (
            .O(N__11642),
            .I(N__11636));
    Span4Mux_v I__2810 (
            .O(N__11639),
            .I(N__11633));
    Span12Mux_h I__2809 (
            .O(N__11636),
            .I(N__11630));
    Sp12to4 I__2808 (
            .O(N__11633),
            .I(N__11627));
    Odrv12 I__2807 (
            .O(N__11630),
            .I(DRA_c_3));
    Odrv12 I__2806 (
            .O(N__11627),
            .I(DRA_c_3));
    InMux I__2805 (
            .O(N__11622),
            .I(N__11619));
    LocalMux I__2804 (
            .O(N__11619),
            .I(N__11615));
    InMux I__2803 (
            .O(N__11618),
            .I(N__11612));
    Span4Mux_v I__2802 (
            .O(N__11615),
            .I(N__11605));
    LocalMux I__2801 (
            .O(N__11612),
            .I(N__11605));
    InMux I__2800 (
            .O(N__11611),
            .I(N__11602));
    InMux I__2799 (
            .O(N__11610),
            .I(N__11599));
    Span4Mux_v I__2798 (
            .O(N__11605),
            .I(N__11596));
    LocalMux I__2797 (
            .O(N__11602),
            .I(N__11593));
    LocalMux I__2796 (
            .O(N__11599),
            .I(N__11590));
    Span4Mux_v I__2795 (
            .O(N__11596),
            .I(N__11587));
    Span4Mux_h I__2794 (
            .O(N__11593),
            .I(N__11584));
    Span12Mux_v I__2793 (
            .O(N__11590),
            .I(N__11579));
    Sp12to4 I__2792 (
            .O(N__11587),
            .I(N__11579));
    Sp12to4 I__2791 (
            .O(N__11584),
            .I(N__11576));
    Span12Mux_h I__2790 (
            .O(N__11579),
            .I(N__11573));
    Span12Mux_v I__2789 (
            .O(N__11576),
            .I(N__11570));
    Odrv12 I__2788 (
            .O(N__11573),
            .I(DRA_c_2));
    Odrv12 I__2787 (
            .O(N__11570),
            .I(DRA_c_2));
    InMux I__2786 (
            .O(N__11565),
            .I(N__11562));
    LocalMux I__2785 (
            .O(N__11562),
            .I(N__11559));
    Span4Mux_h I__2784 (
            .O(N__11559),
            .I(N__11556));
    Odrv4 I__2783 (
            .O(N__11556),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    CascadeMux I__2782 (
            .O(N__11553),
            .I(N__11549));
    InMux I__2781 (
            .O(N__11552),
            .I(N__11545));
    InMux I__2780 (
            .O(N__11549),
            .I(N__11540));
    InMux I__2779 (
            .O(N__11548),
            .I(N__11540));
    LocalMux I__2778 (
            .O(N__11545),
            .I(N__11536));
    LocalMux I__2777 (
            .O(N__11540),
            .I(N__11525));
    InMux I__2776 (
            .O(N__11539),
            .I(N__11522));
    Span4Mux_v I__2775 (
            .O(N__11536),
            .I(N__11519));
    InMux I__2774 (
            .O(N__11535),
            .I(N__11516));
    InMux I__2773 (
            .O(N__11534),
            .I(N__11513));
    InMux I__2772 (
            .O(N__11533),
            .I(N__11510));
    InMux I__2771 (
            .O(N__11532),
            .I(N__11507));
    InMux I__2770 (
            .O(N__11531),
            .I(N__11504));
    InMux I__2769 (
            .O(N__11530),
            .I(N__11501));
    CascadeMux I__2768 (
            .O(N__11529),
            .I(N__11497));
    CascadeMux I__2767 (
            .O(N__11528),
            .I(N__11491));
    Span4Mux_v I__2766 (
            .O(N__11525),
            .I(N__11487));
    LocalMux I__2765 (
            .O(N__11522),
            .I(N__11484));
    Span4Mux_h I__2764 (
            .O(N__11519),
            .I(N__11481));
    LocalMux I__2763 (
            .O(N__11516),
            .I(N__11472));
    LocalMux I__2762 (
            .O(N__11513),
            .I(N__11472));
    LocalMux I__2761 (
            .O(N__11510),
            .I(N__11472));
    LocalMux I__2760 (
            .O(N__11507),
            .I(N__11472));
    LocalMux I__2759 (
            .O(N__11504),
            .I(N__11467));
    LocalMux I__2758 (
            .O(N__11501),
            .I(N__11464));
    InMux I__2757 (
            .O(N__11500),
            .I(N__11455));
    InMux I__2756 (
            .O(N__11497),
            .I(N__11455));
    InMux I__2755 (
            .O(N__11496),
            .I(N__11455));
    InMux I__2754 (
            .O(N__11495),
            .I(N__11455));
    InMux I__2753 (
            .O(N__11494),
            .I(N__11452));
    InMux I__2752 (
            .O(N__11491),
            .I(N__11447));
    InMux I__2751 (
            .O(N__11490),
            .I(N__11447));
    Span4Mux_h I__2750 (
            .O(N__11487),
            .I(N__11440));
    Span4Mux_v I__2749 (
            .O(N__11484),
            .I(N__11440));
    Span4Mux_h I__2748 (
            .O(N__11481),
            .I(N__11435));
    Span4Mux_v I__2747 (
            .O(N__11472),
            .I(N__11435));
    InMux I__2746 (
            .O(N__11471),
            .I(N__11430));
    InMux I__2745 (
            .O(N__11470),
            .I(N__11430));
    Span4Mux_h I__2744 (
            .O(N__11467),
            .I(N__11419));
    Span4Mux_h I__2743 (
            .O(N__11464),
            .I(N__11419));
    LocalMux I__2742 (
            .O(N__11455),
            .I(N__11419));
    LocalMux I__2741 (
            .O(N__11452),
            .I(N__11419));
    LocalMux I__2740 (
            .O(N__11447),
            .I(N__11419));
    InMux I__2739 (
            .O(N__11446),
            .I(N__11414));
    InMux I__2738 (
            .O(N__11445),
            .I(N__11414));
    Sp12to4 I__2737 (
            .O(N__11440),
            .I(N__11409));
    Sp12to4 I__2736 (
            .O(N__11435),
            .I(N__11409));
    LocalMux I__2735 (
            .O(N__11430),
            .I(N__11406));
    Sp12to4 I__2734 (
            .O(N__11419),
            .I(N__11403));
    LocalMux I__2733 (
            .O(N__11414),
            .I(N__11400));
    Span12Mux_h I__2732 (
            .O(N__11409),
            .I(N__11397));
    Span12Mux_v I__2731 (
            .O(N__11406),
            .I(N__11394));
    Span12Mux_v I__2730 (
            .O(N__11403),
            .I(N__11391));
    Span12Mux_h I__2729 (
            .O(N__11400),
            .I(N__11388));
    Span12Mux_v I__2728 (
            .O(N__11397),
            .I(N__11383));
    Span12Mux_h I__2727 (
            .O(N__11394),
            .I(N__11383));
    Span12Mux_h I__2726 (
            .O(N__11391),
            .I(N__11378));
    Span12Mux_v I__2725 (
            .O(N__11388),
            .I(N__11378));
    Odrv12 I__2724 (
            .O(N__11383),
            .I(AGNUS_REV_c));
    Odrv12 I__2723 (
            .O(N__11378),
            .I(AGNUS_REV_c));
    InMux I__2722 (
            .O(N__11373),
            .I(N__11368));
    InMux I__2721 (
            .O(N__11372),
            .I(N__11365));
    InMux I__2720 (
            .O(N__11371),
            .I(N__11361));
    LocalMux I__2719 (
            .O(N__11368),
            .I(N__11358));
    LocalMux I__2718 (
            .O(N__11365),
            .I(N__11355));
    InMux I__2717 (
            .O(N__11364),
            .I(N__11352));
    LocalMux I__2716 (
            .O(N__11361),
            .I(N__11349));
    Span4Mux_v I__2715 (
            .O(N__11358),
            .I(N__11346));
    Span4Mux_v I__2714 (
            .O(N__11355),
            .I(N__11339));
    LocalMux I__2713 (
            .O(N__11352),
            .I(N__11339));
    Span4Mux_v I__2712 (
            .O(N__11349),
            .I(N__11339));
    Sp12to4 I__2711 (
            .O(N__11346),
            .I(N__11334));
    Sp12to4 I__2710 (
            .O(N__11339),
            .I(N__11334));
    Span12Mux_h I__2709 (
            .O(N__11334),
            .I(N__11331));
    Span12Mux_v I__2708 (
            .O(N__11331),
            .I(N__11328));
    Odrv12 I__2707 (
            .O(N__11328),
            .I(DRA_c_1));
    InMux I__2706 (
            .O(N__11325),
            .I(N__11322));
    LocalMux I__2705 (
            .O(N__11322),
            .I(N__11318));
    InMux I__2704 (
            .O(N__11321),
            .I(N__11315));
    Span4Mux_h I__2703 (
            .O(N__11318),
            .I(N__11310));
    LocalMux I__2702 (
            .O(N__11315),
            .I(N__11310));
    Sp12to4 I__2701 (
            .O(N__11310),
            .I(N__11307));
    Span12Mux_v I__2700 (
            .O(N__11307),
            .I(N__11304));
    Span12Mux_h I__2699 (
            .O(N__11304),
            .I(N__11301));
    Odrv12 I__2698 (
            .O(N__11301),
            .I(DRA_c_0));
    InMux I__2697 (
            .O(N__11298),
            .I(N__11295));
    LocalMux I__2696 (
            .O(N__11295),
            .I(N__11292));
    Span4Mux_h I__2695 (
            .O(N__11292),
            .I(N__11289));
    Odrv4 I__2694 (
            .O(N__11289),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    ClkMux I__2693 (
            .O(N__11286),
            .I(N__11268));
    ClkMux I__2692 (
            .O(N__11285),
            .I(N__11268));
    ClkMux I__2691 (
            .O(N__11284),
            .I(N__11268));
    ClkMux I__2690 (
            .O(N__11283),
            .I(N__11268));
    ClkMux I__2689 (
            .O(N__11282),
            .I(N__11268));
    ClkMux I__2688 (
            .O(N__11281),
            .I(N__11268));
    GlobalMux I__2687 (
            .O(N__11268),
            .I(N__11265));
    gio2CtrlBuf I__2686 (
            .O(N__11265),
            .I(C3_c_g));
    CEMux I__2685 (
            .O(N__11262),
            .I(N__11226));
    CEMux I__2684 (
            .O(N__11261),
            .I(N__11226));
    CEMux I__2683 (
            .O(N__11260),
            .I(N__11226));
    CEMux I__2682 (
            .O(N__11259),
            .I(N__11226));
    CEMux I__2681 (
            .O(N__11258),
            .I(N__11226));
    CEMux I__2680 (
            .O(N__11257),
            .I(N__11226));
    CEMux I__2679 (
            .O(N__11256),
            .I(N__11226));
    CEMux I__2678 (
            .O(N__11255),
            .I(N__11226));
    CEMux I__2677 (
            .O(N__11254),
            .I(N__11226));
    CEMux I__2676 (
            .O(N__11253),
            .I(N__11226));
    CEMux I__2675 (
            .O(N__11252),
            .I(N__11226));
    CEMux I__2674 (
            .O(N__11251),
            .I(N__11226));
    GlobalMux I__2673 (
            .O(N__11226),
            .I(N__11223));
    gio2CtrlBuf I__2672 (
            .O(N__11223),
            .I(DBRn_c_i_0_g));
    InMux I__2671 (
            .O(N__11220),
            .I(N__11213));
    InMux I__2670 (
            .O(N__11219),
            .I(N__11210));
    InMux I__2669 (
            .O(N__11218),
            .I(N__11207));
    InMux I__2668 (
            .O(N__11217),
            .I(N__11204));
    InMux I__2667 (
            .O(N__11216),
            .I(N__11201));
    LocalMux I__2666 (
            .O(N__11213),
            .I(N__11198));
    LocalMux I__2665 (
            .O(N__11210),
            .I(N__11181));
    LocalMux I__2664 (
            .O(N__11207),
            .I(N__11178));
    LocalMux I__2663 (
            .O(N__11204),
            .I(N__11164));
    LocalMux I__2662 (
            .O(N__11201),
            .I(N__11151));
    Glb2LocalMux I__2661 (
            .O(N__11198),
            .I(N__11064));
    SRMux I__2660 (
            .O(N__11197),
            .I(N__11064));
    SRMux I__2659 (
            .O(N__11196),
            .I(N__11064));
    SRMux I__2658 (
            .O(N__11195),
            .I(N__11064));
    SRMux I__2657 (
            .O(N__11194),
            .I(N__11064));
    SRMux I__2656 (
            .O(N__11193),
            .I(N__11064));
    SRMux I__2655 (
            .O(N__11192),
            .I(N__11064));
    SRMux I__2654 (
            .O(N__11191),
            .I(N__11064));
    SRMux I__2653 (
            .O(N__11190),
            .I(N__11064));
    SRMux I__2652 (
            .O(N__11189),
            .I(N__11064));
    SRMux I__2651 (
            .O(N__11188),
            .I(N__11064));
    SRMux I__2650 (
            .O(N__11187),
            .I(N__11064));
    SRMux I__2649 (
            .O(N__11186),
            .I(N__11064));
    SRMux I__2648 (
            .O(N__11185),
            .I(N__11064));
    SRMux I__2647 (
            .O(N__11184),
            .I(N__11064));
    Glb2LocalMux I__2646 (
            .O(N__11181),
            .I(N__11064));
    Glb2LocalMux I__2645 (
            .O(N__11178),
            .I(N__11064));
    SRMux I__2644 (
            .O(N__11177),
            .I(N__11064));
    SRMux I__2643 (
            .O(N__11176),
            .I(N__11064));
    SRMux I__2642 (
            .O(N__11175),
            .I(N__11064));
    SRMux I__2641 (
            .O(N__11174),
            .I(N__11064));
    SRMux I__2640 (
            .O(N__11173),
            .I(N__11064));
    SRMux I__2639 (
            .O(N__11172),
            .I(N__11064));
    SRMux I__2638 (
            .O(N__11171),
            .I(N__11064));
    SRMux I__2637 (
            .O(N__11170),
            .I(N__11064));
    SRMux I__2636 (
            .O(N__11169),
            .I(N__11064));
    SRMux I__2635 (
            .O(N__11168),
            .I(N__11064));
    SRMux I__2634 (
            .O(N__11167),
            .I(N__11064));
    Glb2LocalMux I__2633 (
            .O(N__11164),
            .I(N__11064));
    SRMux I__2632 (
            .O(N__11163),
            .I(N__11064));
    SRMux I__2631 (
            .O(N__11162),
            .I(N__11064));
    SRMux I__2630 (
            .O(N__11161),
            .I(N__11064));
    SRMux I__2629 (
            .O(N__11160),
            .I(N__11064));
    SRMux I__2628 (
            .O(N__11159),
            .I(N__11064));
    SRMux I__2627 (
            .O(N__11158),
            .I(N__11064));
    SRMux I__2626 (
            .O(N__11157),
            .I(N__11064));
    SRMux I__2625 (
            .O(N__11156),
            .I(N__11064));
    SRMux I__2624 (
            .O(N__11155),
            .I(N__11064));
    SRMux I__2623 (
            .O(N__11154),
            .I(N__11064));
    Glb2LocalMux I__2622 (
            .O(N__11151),
            .I(N__11064));
    SRMux I__2621 (
            .O(N__11150),
            .I(N__11064));
    SRMux I__2620 (
            .O(N__11149),
            .I(N__11064));
    GlobalMux I__2619 (
            .O(N__11064),
            .I(N__11061));
    gio2CtrlBuf I__2618 (
            .O(N__11061),
            .I(RESETn_c_i_g));
    InMux I__2617 (
            .O(N__11058),
            .I(N__11055));
    LocalMux I__2616 (
            .O(N__11055),
            .I(N__11052));
    Span12Mux_v I__2615 (
            .O(N__11052),
            .I(N__11049));
    Span12Mux_h I__2614 (
            .O(N__11049),
            .I(N__11046));
    Odrv12 I__2613 (
            .O(N__11046),
            .I(RAS1n_c));
    InMux I__2612 (
            .O(N__11043),
            .I(N__11039));
    InMux I__2611 (
            .O(N__11042),
            .I(N__11036));
    LocalMux I__2610 (
            .O(N__11039),
            .I(N__11033));
    LocalMux I__2609 (
            .O(N__11036),
            .I(N__11030));
    Span4Mux_v I__2608 (
            .O(N__11033),
            .I(N__11027));
    Span12Mux_h I__2607 (
            .O(N__11030),
            .I(N__11024));
    Sp12to4 I__2606 (
            .O(N__11027),
            .I(N__11021));
    Odrv12 I__2605 (
            .O(N__11024),
            .I(RAS0n_c));
    Odrv12 I__2604 (
            .O(N__11021),
            .I(RAS0n_c));
    InMux I__2603 (
            .O(N__11016),
            .I(N__11013));
    LocalMux I__2602 (
            .O(N__11013),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2601 (
            .O(N__11010),
            .I(N__10993));
    InMux I__2600 (
            .O(N__11009),
            .I(N__10990));
    InMux I__2599 (
            .O(N__11008),
            .I(N__10987));
    InMux I__2598 (
            .O(N__11007),
            .I(N__10982));
    InMux I__2597 (
            .O(N__11006),
            .I(N__10982));
    InMux I__2596 (
            .O(N__11005),
            .I(N__10977));
    InMux I__2595 (
            .O(N__11004),
            .I(N__10977));
    InMux I__2594 (
            .O(N__11003),
            .I(N__10972));
    InMux I__2593 (
            .O(N__11002),
            .I(N__10972));
    InMux I__2592 (
            .O(N__11001),
            .I(N__10969));
    InMux I__2591 (
            .O(N__11000),
            .I(N__10966));
    InMux I__2590 (
            .O(N__10999),
            .I(N__10963));
    InMux I__2589 (
            .O(N__10998),
            .I(N__10949));
    InMux I__2588 (
            .O(N__10997),
            .I(N__10949));
    CascadeMux I__2587 (
            .O(N__10996),
            .I(N__10944));
    LocalMux I__2586 (
            .O(N__10993),
            .I(N__10938));
    LocalMux I__2585 (
            .O(N__10990),
            .I(N__10923));
    LocalMux I__2584 (
            .O(N__10987),
            .I(N__10923));
    LocalMux I__2583 (
            .O(N__10982),
            .I(N__10923));
    LocalMux I__2582 (
            .O(N__10977),
            .I(N__10923));
    LocalMux I__2581 (
            .O(N__10972),
            .I(N__10923));
    LocalMux I__2580 (
            .O(N__10969),
            .I(N__10923));
    LocalMux I__2579 (
            .O(N__10966),
            .I(N__10923));
    LocalMux I__2578 (
            .O(N__10963),
            .I(N__10920));
    InMux I__2577 (
            .O(N__10962),
            .I(N__10917));
    InMux I__2576 (
            .O(N__10961),
            .I(N__10914));
    InMux I__2575 (
            .O(N__10960),
            .I(N__10909));
    InMux I__2574 (
            .O(N__10959),
            .I(N__10909));
    InMux I__2573 (
            .O(N__10958),
            .I(N__10902));
    InMux I__2572 (
            .O(N__10957),
            .I(N__10902));
    InMux I__2571 (
            .O(N__10956),
            .I(N__10902));
    InMux I__2570 (
            .O(N__10955),
            .I(N__10897));
    InMux I__2569 (
            .O(N__10954),
            .I(N__10897));
    LocalMux I__2568 (
            .O(N__10949),
            .I(N__10894));
    InMux I__2567 (
            .O(N__10948),
            .I(N__10891));
    InMux I__2566 (
            .O(N__10947),
            .I(N__10888));
    InMux I__2565 (
            .O(N__10944),
            .I(N__10881));
    InMux I__2564 (
            .O(N__10943),
            .I(N__10881));
    InMux I__2563 (
            .O(N__10942),
            .I(N__10881));
    InMux I__2562 (
            .O(N__10941),
            .I(N__10878));
    Span4Mux_v I__2561 (
            .O(N__10938),
            .I(N__10870));
    Span4Mux_v I__2560 (
            .O(N__10923),
            .I(N__10870));
    Span4Mux_v I__2559 (
            .O(N__10920),
            .I(N__10863));
    LocalMux I__2558 (
            .O(N__10917),
            .I(N__10863));
    LocalMux I__2557 (
            .O(N__10914),
            .I(N__10863));
    LocalMux I__2556 (
            .O(N__10909),
            .I(N__10860));
    LocalMux I__2555 (
            .O(N__10902),
            .I(N__10855));
    LocalMux I__2554 (
            .O(N__10897),
            .I(N__10855));
    Span4Mux_v I__2553 (
            .O(N__10894),
            .I(N__10844));
    LocalMux I__2552 (
            .O(N__10891),
            .I(N__10844));
    LocalMux I__2551 (
            .O(N__10888),
            .I(N__10844));
    LocalMux I__2550 (
            .O(N__10881),
            .I(N__10844));
    LocalMux I__2549 (
            .O(N__10878),
            .I(N__10844));
    CascadeMux I__2548 (
            .O(N__10877),
            .I(N__10841));
    InMux I__2547 (
            .O(N__10876),
            .I(N__10835));
    InMux I__2546 (
            .O(N__10875),
            .I(N__10835));
    Span4Mux_h I__2545 (
            .O(N__10870),
            .I(N__10829));
    Span4Mux_v I__2544 (
            .O(N__10863),
            .I(N__10829));
    Span4Mux_v I__2543 (
            .O(N__10860),
            .I(N__10822));
    Span4Mux_h I__2542 (
            .O(N__10855),
            .I(N__10822));
    Span4Mux_v I__2541 (
            .O(N__10844),
            .I(N__10822));
    InMux I__2540 (
            .O(N__10841),
            .I(N__10819));
    InMux I__2539 (
            .O(N__10840),
            .I(N__10816));
    LocalMux I__2538 (
            .O(N__10835),
            .I(N__10813));
    InMux I__2537 (
            .O(N__10834),
            .I(N__10810));
    Sp12to4 I__2536 (
            .O(N__10829),
            .I(N__10801));
    Sp12to4 I__2535 (
            .O(N__10822),
            .I(N__10801));
    LocalMux I__2534 (
            .O(N__10819),
            .I(N__10801));
    LocalMux I__2533 (
            .O(N__10816),
            .I(N__10801));
    Span12Mux_v I__2532 (
            .O(N__10813),
            .I(N__10796));
    LocalMux I__2531 (
            .O(N__10810),
            .I(N__10796));
    Span12Mux_h I__2530 (
            .O(N__10801),
            .I(N__10793));
    Span12Mux_h I__2529 (
            .O(N__10796),
            .I(N__10790));
    Odrv12 I__2528 (
            .O(N__10793),
            .I(RESETn_c));
    Odrv12 I__2527 (
            .O(N__10790),
            .I(RESETn_c));
    InMux I__2526 (
            .O(N__10785),
            .I(N__10782));
    LocalMux I__2525 (
            .O(N__10782),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    InMux I__2524 (
            .O(N__10779),
            .I(N__10776));
    LocalMux I__2523 (
            .O(N__10776),
            .I(N__10773));
    Odrv12 I__2522 (
            .O(N__10773),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ));
    InMux I__2521 (
            .O(N__10770),
            .I(N__10767));
    LocalMux I__2520 (
            .O(N__10767),
            .I(N__10725));
    ClkMux I__2519 (
            .O(N__10766),
            .I(N__10623));
    ClkMux I__2518 (
            .O(N__10765),
            .I(N__10623));
    ClkMux I__2517 (
            .O(N__10764),
            .I(N__10623));
    ClkMux I__2516 (
            .O(N__10763),
            .I(N__10623));
    ClkMux I__2515 (
            .O(N__10762),
            .I(N__10623));
    ClkMux I__2514 (
            .O(N__10761),
            .I(N__10623));
    ClkMux I__2513 (
            .O(N__10760),
            .I(N__10623));
    ClkMux I__2512 (
            .O(N__10759),
            .I(N__10623));
    ClkMux I__2511 (
            .O(N__10758),
            .I(N__10623));
    ClkMux I__2510 (
            .O(N__10757),
            .I(N__10623));
    ClkMux I__2509 (
            .O(N__10756),
            .I(N__10623));
    ClkMux I__2508 (
            .O(N__10755),
            .I(N__10623));
    ClkMux I__2507 (
            .O(N__10754),
            .I(N__10623));
    ClkMux I__2506 (
            .O(N__10753),
            .I(N__10623));
    ClkMux I__2505 (
            .O(N__10752),
            .I(N__10623));
    ClkMux I__2504 (
            .O(N__10751),
            .I(N__10623));
    ClkMux I__2503 (
            .O(N__10750),
            .I(N__10623));
    ClkMux I__2502 (
            .O(N__10749),
            .I(N__10623));
    ClkMux I__2501 (
            .O(N__10748),
            .I(N__10623));
    ClkMux I__2500 (
            .O(N__10747),
            .I(N__10623));
    ClkMux I__2499 (
            .O(N__10746),
            .I(N__10623));
    ClkMux I__2498 (
            .O(N__10745),
            .I(N__10623));
    ClkMux I__2497 (
            .O(N__10744),
            .I(N__10623));
    ClkMux I__2496 (
            .O(N__10743),
            .I(N__10623));
    ClkMux I__2495 (
            .O(N__10742),
            .I(N__10623));
    ClkMux I__2494 (
            .O(N__10741),
            .I(N__10623));
    ClkMux I__2493 (
            .O(N__10740),
            .I(N__10623));
    ClkMux I__2492 (
            .O(N__10739),
            .I(N__10623));
    ClkMux I__2491 (
            .O(N__10738),
            .I(N__10623));
    ClkMux I__2490 (
            .O(N__10737),
            .I(N__10623));
    ClkMux I__2489 (
            .O(N__10736),
            .I(N__10623));
    ClkMux I__2488 (
            .O(N__10735),
            .I(N__10623));
    ClkMux I__2487 (
            .O(N__10734),
            .I(N__10623));
    ClkMux I__2486 (
            .O(N__10733),
            .I(N__10623));
    ClkMux I__2485 (
            .O(N__10732),
            .I(N__10623));
    ClkMux I__2484 (
            .O(N__10731),
            .I(N__10623));
    ClkMux I__2483 (
            .O(N__10730),
            .I(N__10623));
    ClkMux I__2482 (
            .O(N__10729),
            .I(N__10623));
    ClkMux I__2481 (
            .O(N__10728),
            .I(N__10623));
    Glb2LocalMux I__2480 (
            .O(N__10725),
            .I(N__10623));
    ClkMux I__2479 (
            .O(N__10724),
            .I(N__10623));
    ClkMux I__2478 (
            .O(N__10723),
            .I(N__10623));
    ClkMux I__2477 (
            .O(N__10722),
            .I(N__10623));
    ClkMux I__2476 (
            .O(N__10721),
            .I(N__10623));
    ClkMux I__2475 (
            .O(N__10720),
            .I(N__10623));
    ClkMux I__2474 (
            .O(N__10719),
            .I(N__10623));
    ClkMux I__2473 (
            .O(N__10718),
            .I(N__10623));
    GlobalMux I__2472 (
            .O(N__10623),
            .I(CLK80_PLL));
    InMux I__2471 (
            .O(N__10620),
            .I(N__10616));
    InMux I__2470 (
            .O(N__10619),
            .I(N__10613));
    LocalMux I__2469 (
            .O(N__10616),
            .I(N__10610));
    LocalMux I__2468 (
            .O(N__10613),
            .I(N__10607));
    Span12Mux_v I__2467 (
            .O(N__10610),
            .I(N__10604));
    Span4Mux_v I__2466 (
            .O(N__10607),
            .I(N__10601));
    Span12Mux_h I__2465 (
            .O(N__10604),
            .I(N__10597));
    Span4Mux_v I__2464 (
            .O(N__10601),
            .I(N__10594));
    InMux I__2463 (
            .O(N__10600),
            .I(N__10591));
    Odrv12 I__2462 (
            .O(N__10597),
            .I(DMA_WRITE_CYCLE));
    Odrv4 I__2461 (
            .O(N__10594),
            .I(DMA_WRITE_CYCLE));
    LocalMux I__2460 (
            .O(N__10591),
            .I(DMA_WRITE_CYCLE));
    InMux I__2459 (
            .O(N__10584),
            .I(N__10580));
    InMux I__2458 (
            .O(N__10583),
            .I(N__10576));
    LocalMux I__2457 (
            .O(N__10580),
            .I(N__10572));
    InMux I__2456 (
            .O(N__10579),
            .I(N__10569));
    LocalMux I__2455 (
            .O(N__10576),
            .I(N__10566));
    CascadeMux I__2454 (
            .O(N__10575),
            .I(N__10563));
    Span4Mux_v I__2453 (
            .O(N__10572),
            .I(N__10560));
    LocalMux I__2452 (
            .O(N__10569),
            .I(N__10557));
    Span4Mux_v I__2451 (
            .O(N__10566),
            .I(N__10553));
    InMux I__2450 (
            .O(N__10563),
            .I(N__10550));
    Span4Mux_h I__2449 (
            .O(N__10560),
            .I(N__10545));
    Span4Mux_v I__2448 (
            .O(N__10557),
            .I(N__10545));
    InMux I__2447 (
            .O(N__10556),
            .I(N__10542));
    Span4Mux_v I__2446 (
            .O(N__10553),
            .I(N__10539));
    LocalMux I__2445 (
            .O(N__10550),
            .I(N__10536));
    Sp12to4 I__2444 (
            .O(N__10545),
            .I(N__10531));
    LocalMux I__2443 (
            .O(N__10542),
            .I(N__10531));
    Sp12to4 I__2442 (
            .O(N__10539),
            .I(N__10528));
    Sp12to4 I__2441 (
            .O(N__10536),
            .I(N__10525));
    Span12Mux_h I__2440 (
            .O(N__10531),
            .I(N__10522));
    Span12Mux_h I__2439 (
            .O(N__10528),
            .I(N__10517));
    Span12Mux_v I__2438 (
            .O(N__10525),
            .I(N__10517));
    Span12Mux_v I__2437 (
            .O(N__10522),
            .I(N__10512));
    Span12Mux_h I__2436 (
            .O(N__10517),
            .I(N__10512));
    Odrv12 I__2435 (
            .O(N__10512),
            .I(RnW_c));
    InMux I__2434 (
            .O(N__10509),
            .I(N__10504));
    InMux I__2433 (
            .O(N__10508),
            .I(N__10501));
    CascadeMux I__2432 (
            .O(N__10507),
            .I(N__10495));
    LocalMux I__2431 (
            .O(N__10504),
            .I(N__10492));
    LocalMux I__2430 (
            .O(N__10501),
            .I(N__10489));
    InMux I__2429 (
            .O(N__10500),
            .I(N__10486));
    InMux I__2428 (
            .O(N__10499),
            .I(N__10479));
    InMux I__2427 (
            .O(N__10498),
            .I(N__10479));
    InMux I__2426 (
            .O(N__10495),
            .I(N__10479));
    Span4Mux_v I__2425 (
            .O(N__10492),
            .I(N__10471));
    Span4Mux_h I__2424 (
            .O(N__10489),
            .I(N__10471));
    LocalMux I__2423 (
            .O(N__10486),
            .I(N__10471));
    LocalMux I__2422 (
            .O(N__10479),
            .I(N__10468));
    InMux I__2421 (
            .O(N__10478),
            .I(N__10465));
    Span4Mux_h I__2420 (
            .O(N__10471),
            .I(N__10460));
    Span4Mux_h I__2419 (
            .O(N__10468),
            .I(N__10455));
    LocalMux I__2418 (
            .O(N__10465),
            .I(N__10455));
    InMux I__2417 (
            .O(N__10464),
            .I(N__10450));
    InMux I__2416 (
            .O(N__10463),
            .I(N__10450));
    Span4Mux_v I__2415 (
            .O(N__10460),
            .I(N__10445));
    Span4Mux_h I__2414 (
            .O(N__10455),
            .I(N__10445));
    LocalMux I__2413 (
            .O(N__10450),
            .I(N__10442));
    Span4Mux_v I__2412 (
            .O(N__10445),
            .I(N__10439));
    Span12Mux_v I__2411 (
            .O(N__10442),
            .I(N__10436));
    Span4Mux_h I__2410 (
            .O(N__10439),
            .I(N__10433));
    Span12Mux_h I__2409 (
            .O(N__10436),
            .I(N__10430));
    Sp12to4 I__2408 (
            .O(N__10433),
            .I(N__10427));
    Odrv12 I__2407 (
            .O(N__10430),
            .I(SIZ_c_1));
    Odrv12 I__2406 (
            .O(N__10427),
            .I(SIZ_c_1));
    CascadeMux I__2405 (
            .O(N__10422),
            .I(N__10417));
    InMux I__2404 (
            .O(N__10421),
            .I(N__10412));
    InMux I__2403 (
            .O(N__10420),
            .I(N__10409));
    InMux I__2402 (
            .O(N__10417),
            .I(N__10406));
    CascadeMux I__2401 (
            .O(N__10416),
            .I(N__10402));
    CascadeMux I__2400 (
            .O(N__10415),
            .I(N__10399));
    LocalMux I__2399 (
            .O(N__10412),
            .I(N__10394));
    LocalMux I__2398 (
            .O(N__10409),
            .I(N__10391));
    LocalMux I__2397 (
            .O(N__10406),
            .I(N__10388));
    InMux I__2396 (
            .O(N__10405),
            .I(N__10385));
    InMux I__2395 (
            .O(N__10402),
            .I(N__10378));
    InMux I__2394 (
            .O(N__10399),
            .I(N__10378));
    InMux I__2393 (
            .O(N__10398),
            .I(N__10378));
    CascadeMux I__2392 (
            .O(N__10397),
            .I(N__10375));
    Span4Mux_v I__2391 (
            .O(N__10394),
            .I(N__10372));
    Span4Mux_v I__2390 (
            .O(N__10391),
            .I(N__10365));
    Span4Mux_h I__2389 (
            .O(N__10388),
            .I(N__10365));
    LocalMux I__2388 (
            .O(N__10385),
            .I(N__10365));
    LocalMux I__2387 (
            .O(N__10378),
            .I(N__10362));
    InMux I__2386 (
            .O(N__10375),
            .I(N__10359));
    Span4Mux_v I__2385 (
            .O(N__10372),
            .I(N__10356));
    Span4Mux_h I__2384 (
            .O(N__10365),
            .I(N__10353));
    Span4Mux_h I__2383 (
            .O(N__10362),
            .I(N__10348));
    LocalMux I__2382 (
            .O(N__10359),
            .I(N__10348));
    Span4Mux_v I__2381 (
            .O(N__10356),
            .I(N__10345));
    Span4Mux_v I__2380 (
            .O(N__10353),
            .I(N__10340));
    Span4Mux_h I__2379 (
            .O(N__10348),
            .I(N__10340));
    Span4Mux_h I__2378 (
            .O(N__10345),
            .I(N__10337));
    Span4Mux_v I__2377 (
            .O(N__10340),
            .I(N__10334));
    Sp12to4 I__2376 (
            .O(N__10337),
            .I(N__10329));
    Sp12to4 I__2375 (
            .O(N__10334),
            .I(N__10329));
    Odrv12 I__2374 (
            .O(N__10329),
            .I(SIZ_c_0));
    IoInMux I__2373 (
            .O(N__10326),
            .I(N__10323));
    LocalMux I__2372 (
            .O(N__10323),
            .I(N__10320));
    Span12Mux_s6_v I__2371 (
            .O(N__10320),
            .I(N__10317));
    Odrv12 I__2370 (
            .O(N__10317),
            .I(N_189));
    InMux I__2369 (
            .O(N__10314),
            .I(N__10311));
    LocalMux I__2368 (
            .O(N__10311),
            .I(N__10308));
    Odrv4 I__2367 (
            .O(N__10308),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__2366 (
            .O(N__10305),
            .I(N__10300));
    InMux I__2365 (
            .O(N__10304),
            .I(N__10297));
    InMux I__2364 (
            .O(N__10303),
            .I(N__10293));
    LocalMux I__2363 (
            .O(N__10300),
            .I(N__10288));
    LocalMux I__2362 (
            .O(N__10297),
            .I(N__10288));
    InMux I__2361 (
            .O(N__10296),
            .I(N__10285));
    LocalMux I__2360 (
            .O(N__10293),
            .I(N__10282));
    Span4Mux_v I__2359 (
            .O(N__10288),
            .I(N__10277));
    LocalMux I__2358 (
            .O(N__10285),
            .I(N__10277));
    Span4Mux_v I__2357 (
            .O(N__10282),
            .I(N__10274));
    Span4Mux_h I__2356 (
            .O(N__10277),
            .I(N__10271));
    Span4Mux_v I__2355 (
            .O(N__10274),
            .I(N__10268));
    Span4Mux_v I__2354 (
            .O(N__10271),
            .I(N__10265));
    Sp12to4 I__2353 (
            .O(N__10268),
            .I(N__10260));
    Sp12to4 I__2352 (
            .O(N__10265),
            .I(N__10260));
    Span12Mux_h I__2351 (
            .O(N__10260),
            .I(N__10257));
    Odrv12 I__2350 (
            .O(N__10257),
            .I(DRA_c_4));
    CascadeMux I__2349 (
            .O(N__10254),
            .I(N__10251));
    InMux I__2348 (
            .O(N__10251),
            .I(N__10248));
    LocalMux I__2347 (
            .O(N__10248),
            .I(N__10245));
    Odrv12 I__2346 (
            .O(N__10245),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2345 (
            .O(N__10242),
            .I(N__10235));
    InMux I__2344 (
            .O(N__10241),
            .I(N__10235));
    InMux I__2343 (
            .O(N__10240),
            .I(N__10232));
    LocalMux I__2342 (
            .O(N__10235),
            .I(N__10226));
    LocalMux I__2341 (
            .O(N__10232),
            .I(N__10226));
    InMux I__2340 (
            .O(N__10231),
            .I(N__10223));
    Span4Mux_v I__2339 (
            .O(N__10226),
            .I(N__10220));
    LocalMux I__2338 (
            .O(N__10223),
            .I(N__10217));
    Sp12to4 I__2337 (
            .O(N__10220),
            .I(N__10212));
    Span12Mux_v I__2336 (
            .O(N__10217),
            .I(N__10212));
    Span12Mux_h I__2335 (
            .O(N__10212),
            .I(N__10209));
    Odrv12 I__2334 (
            .O(N__10209),
            .I(DRA_c_6));
    InMux I__2333 (
            .O(N__10206),
            .I(N__10203));
    LocalMux I__2332 (
            .O(N__10203),
            .I(N__10199));
    InMux I__2331 (
            .O(N__10202),
            .I(N__10196));
    Span4Mux_h I__2330 (
            .O(N__10199),
            .I(N__10189));
    LocalMux I__2329 (
            .O(N__10196),
            .I(N__10189));
    InMux I__2328 (
            .O(N__10195),
            .I(N__10186));
    InMux I__2327 (
            .O(N__10194),
            .I(N__10183));
    Span4Mux_v I__2326 (
            .O(N__10189),
            .I(N__10180));
    LocalMux I__2325 (
            .O(N__10186),
            .I(N__10175));
    LocalMux I__2324 (
            .O(N__10183),
            .I(N__10175));
    Sp12to4 I__2323 (
            .O(N__10180),
            .I(N__10170));
    Span12Mux_v I__2322 (
            .O(N__10175),
            .I(N__10170));
    Span12Mux_h I__2321 (
            .O(N__10170),
            .I(N__10167));
    Odrv12 I__2320 (
            .O(N__10167),
            .I(DRA_c_5));
    InMux I__2319 (
            .O(N__10164),
            .I(N__10161));
    LocalMux I__2318 (
            .O(N__10161),
            .I(N__10158));
    Span4Mux_v I__2317 (
            .O(N__10158),
            .I(N__10155));
    Odrv4 I__2316 (
            .O(N__10155),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2315 (
            .O(N__10152),
            .I(N__10149));
    LocalMux I__2314 (
            .O(N__10149),
            .I(N__10144));
    InMux I__2313 (
            .O(N__10148),
            .I(N__10139));
    InMux I__2312 (
            .O(N__10147),
            .I(N__10139));
    Span4Mux_h I__2311 (
            .O(N__10144),
            .I(N__10134));
    LocalMux I__2310 (
            .O(N__10139),
            .I(N__10134));
    Span4Mux_h I__2309 (
            .O(N__10134),
            .I(N__10130));
    InMux I__2308 (
            .O(N__10133),
            .I(N__10127));
    Span4Mux_v I__2307 (
            .O(N__10130),
            .I(N__10124));
    LocalMux I__2306 (
            .O(N__10127),
            .I(N__10121));
    Sp12to4 I__2305 (
            .O(N__10124),
            .I(N__10118));
    Sp12to4 I__2304 (
            .O(N__10121),
            .I(N__10115));
    Span12Mux_h I__2303 (
            .O(N__10118),
            .I(N__10112));
    Span12Mux_v I__2302 (
            .O(N__10115),
            .I(N__10109));
    Span12Mux_v I__2301 (
            .O(N__10112),
            .I(N__10104));
    Span12Mux_h I__2300 (
            .O(N__10109),
            .I(N__10104));
    Odrv12 I__2299 (
            .O(N__10104),
            .I(DRA_c_9));
    InMux I__2298 (
            .O(N__10101),
            .I(N__10098));
    LocalMux I__2297 (
            .O(N__10098),
            .I(N__10095));
    Odrv12 I__2296 (
            .O(N__10095),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__2295 (
            .O(N__10092),
            .I(N__10088));
    InMux I__2294 (
            .O(N__10091),
            .I(N__10085));
    LocalMux I__2293 (
            .O(N__10088),
            .I(N__10082));
    LocalMux I__2292 (
            .O(N__10085),
            .I(N__10079));
    Span4Mux_v I__2291 (
            .O(N__10082),
            .I(N__10073));
    Span4Mux_h I__2290 (
            .O(N__10079),
            .I(N__10073));
    InMux I__2289 (
            .O(N__10078),
            .I(N__10068));
    Span4Mux_h I__2288 (
            .O(N__10073),
            .I(N__10065));
    InMux I__2287 (
            .O(N__10072),
            .I(N__10062));
    InMux I__2286 (
            .O(N__10071),
            .I(N__10059));
    LocalMux I__2285 (
            .O(N__10068),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__2284 (
            .O(N__10065),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__2283 (
            .O(N__10062),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__2282 (
            .O(N__10059),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__2281 (
            .O(N__10050),
            .I(N__10047));
    LocalMux I__2280 (
            .O(N__10047),
            .I(N__10044));
    Span4Mux_s3_v I__2279 (
            .O(N__10044),
            .I(N__10041));
    Span4Mux_v I__2278 (
            .O(N__10041),
            .I(N__10038));
    Span4Mux_h I__2277 (
            .O(N__10038),
            .I(N__10035));
    Odrv4 I__2276 (
            .O(N__10035),
            .I(CRCSn_c));
    InMux I__2275 (
            .O(N__10032),
            .I(N__10029));
    LocalMux I__2274 (
            .O(N__10029),
            .I(N__10024));
    InMux I__2273 (
            .O(N__10028),
            .I(N__10021));
    InMux I__2272 (
            .O(N__10027),
            .I(N__10018));
    Span12Mux_h I__2271 (
            .O(N__10024),
            .I(N__10014));
    LocalMux I__2270 (
            .O(N__10021),
            .I(N__10011));
    LocalMux I__2269 (
            .O(N__10018),
            .I(N__10008));
    InMux I__2268 (
            .O(N__10017),
            .I(N__10005));
    Odrv12 I__2267 (
            .O(N__10014),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__2266 (
            .O(N__10011),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__2265 (
            .O(N__10008),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__2264 (
            .O(N__10005),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__2263 (
            .O(N__9996),
            .I(N__9993));
    LocalMux I__2262 (
            .O(N__9993),
            .I(N__9990));
    Span12Mux_s5_h I__2261 (
            .O(N__9990),
            .I(N__9987));
    Span12Mux_v I__2260 (
            .O(N__9987),
            .I(N__9984));
    Odrv12 I__2259 (
            .O(N__9984),
            .I(WEn_c));
    InMux I__2258 (
            .O(N__9981),
            .I(N__9978));
    LocalMux I__2257 (
            .O(N__9978),
            .I(N__9975));
    Span4Mux_h I__2256 (
            .O(N__9975),
            .I(N__9972));
    Odrv4 I__2255 (
            .O(N__9972),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__2254 (
            .O(N__9969),
            .I(N__9966));
    LocalMux I__2253 (
            .O(N__9966),
            .I(N__9963));
    Odrv12 I__2252 (
            .O(N__9963),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__2251 (
            .O(N__9960),
            .I(N__9957));
    LocalMux I__2250 (
            .O(N__9957),
            .I(N__9954));
    Span4Mux_h I__2249 (
            .O(N__9954),
            .I(N__9951));
    Odrv4 I__2248 (
            .O(N__9951),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    CascadeMux I__2247 (
            .O(N__9948),
            .I(N__9945));
    InMux I__2246 (
            .O(N__9945),
            .I(N__9942));
    LocalMux I__2245 (
            .O(N__9942),
            .I(N__9939));
    Odrv4 I__2244 (
            .O(N__9939),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2243 (
            .O(N__9936),
            .I(N__9933));
    LocalMux I__2242 (
            .O(N__9933),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__2241 (
            .O(N__9930),
            .I(N__9927));
    LocalMux I__2240 (
            .O(N__9927),
            .I(N__9924));
    Odrv4 I__2239 (
            .O(N__9924),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    CascadeMux I__2238 (
            .O(N__9921),
            .I(N__9917));
    InMux I__2237 (
            .O(N__9920),
            .I(N__9912));
    InMux I__2236 (
            .O(N__9917),
            .I(N__9912));
    LocalMux I__2235 (
            .O(N__9912),
            .I(\U712_BYTE_ENABLE.N_298_i ));
    InMux I__2234 (
            .O(N__9909),
            .I(N__9906));
    LocalMux I__2233 (
            .O(N__9906),
            .I(\U712_REG_SM.N_459 ));
    IoInMux I__2232 (
            .O(N__9903),
            .I(N__9900));
    LocalMux I__2231 (
            .O(N__9900),
            .I(N__9897));
    Span4Mux_s2_v I__2230 (
            .O(N__9897),
            .I(N__9894));
    Span4Mux_v I__2229 (
            .O(N__9894),
            .I(N__9891));
    Odrv4 I__2228 (
            .O(N__9891),
            .I(N_390_i));
    IoInMux I__2227 (
            .O(N__9888),
            .I(N__9885));
    LocalMux I__2226 (
            .O(N__9885),
            .I(N__9882));
    Span4Mux_s2_v I__2225 (
            .O(N__9882),
            .I(N__9879));
    Span4Mux_v I__2224 (
            .O(N__9879),
            .I(N__9876));
    Odrv4 I__2223 (
            .O(N__9876),
            .I(N_389_i));
    InMux I__2222 (
            .O(N__9873),
            .I(N__9860));
    InMux I__2221 (
            .O(N__9872),
            .I(N__9860));
    InMux I__2220 (
            .O(N__9871),
            .I(N__9860));
    InMux I__2219 (
            .O(N__9870),
            .I(N__9855));
    InMux I__2218 (
            .O(N__9869),
            .I(N__9855));
    InMux I__2217 (
            .O(N__9868),
            .I(N__9851));
    InMux I__2216 (
            .O(N__9867),
            .I(N__9848));
    LocalMux I__2215 (
            .O(N__9860),
            .I(N__9845));
    LocalMux I__2214 (
            .O(N__9855),
            .I(N__9842));
    InMux I__2213 (
            .O(N__9854),
            .I(N__9839));
    LocalMux I__2212 (
            .O(N__9851),
            .I(N__9836));
    LocalMux I__2211 (
            .O(N__9848),
            .I(N__9832));
    Span4Mux_v I__2210 (
            .O(N__9845),
            .I(N__9827));
    Span4Mux_v I__2209 (
            .O(N__9842),
            .I(N__9827));
    LocalMux I__2208 (
            .O(N__9839),
            .I(N__9824));
    Span4Mux_v I__2207 (
            .O(N__9836),
            .I(N__9821));
    InMux I__2206 (
            .O(N__9835),
            .I(N__9818));
    Span12Mux_s10_v I__2205 (
            .O(N__9832),
            .I(N__9807));
    Sp12to4 I__2204 (
            .O(N__9827),
            .I(N__9807));
    Span12Mux_h I__2203 (
            .O(N__9824),
            .I(N__9807));
    Sp12to4 I__2202 (
            .O(N__9821),
            .I(N__9807));
    LocalMux I__2201 (
            .O(N__9818),
            .I(N__9807));
    Span12Mux_h I__2200 (
            .O(N__9807),
            .I(N__9804));
    Odrv12 I__2199 (
            .O(N__9804),
            .I(A_c_0));
    InMux I__2198 (
            .O(N__9801),
            .I(N__9797));
    InMux I__2197 (
            .O(N__9800),
            .I(N__9794));
    LocalMux I__2196 (
            .O(N__9797),
            .I(N__9786));
    LocalMux I__2195 (
            .O(N__9794),
            .I(N__9783));
    InMux I__2194 (
            .O(N__9793),
            .I(N__9776));
    InMux I__2193 (
            .O(N__9792),
            .I(N__9776));
    InMux I__2192 (
            .O(N__9791),
            .I(N__9776));
    InMux I__2191 (
            .O(N__9790),
            .I(N__9770));
    InMux I__2190 (
            .O(N__9789),
            .I(N__9770));
    Span4Mux_v I__2189 (
            .O(N__9786),
            .I(N__9767));
    Span4Mux_v I__2188 (
            .O(N__9783),
            .I(N__9764));
    LocalMux I__2187 (
            .O(N__9776),
            .I(N__9761));
    InMux I__2186 (
            .O(N__9775),
            .I(N__9758));
    LocalMux I__2185 (
            .O(N__9770),
            .I(N__9755));
    Span4Mux_v I__2184 (
            .O(N__9767),
            .I(N__9752));
    Span4Mux_v I__2183 (
            .O(N__9764),
            .I(N__9747));
    Span4Mux_v I__2182 (
            .O(N__9761),
            .I(N__9747));
    LocalMux I__2181 (
            .O(N__9758),
            .I(N__9744));
    Span12Mux_v I__2180 (
            .O(N__9755),
            .I(N__9735));
    Sp12to4 I__2179 (
            .O(N__9752),
            .I(N__9735));
    Sp12to4 I__2178 (
            .O(N__9747),
            .I(N__9735));
    Span12Mux_s7_v I__2177 (
            .O(N__9744),
            .I(N__9735));
    Span12Mux_h I__2176 (
            .O(N__9735),
            .I(N__9732));
    Odrv12 I__2175 (
            .O(N__9732),
            .I(A_c_1));
    InMux I__2174 (
            .O(N__9729),
            .I(N__9725));
    InMux I__2173 (
            .O(N__9728),
            .I(N__9721));
    LocalMux I__2172 (
            .O(N__9725),
            .I(N__9717));
    InMux I__2171 (
            .O(N__9724),
            .I(N__9714));
    LocalMux I__2170 (
            .O(N__9721),
            .I(N__9711));
    InMux I__2169 (
            .O(N__9720),
            .I(N__9708));
    Odrv4 I__2168 (
            .O(N__9717),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__2167 (
            .O(N__9714),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    Odrv4 I__2166 (
            .O(N__9711),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__2165 (
            .O(N__9708),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__2164 (
            .O(N__9699),
            .I(N__9696));
    LocalMux I__2163 (
            .O(N__9696),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ));
    CascadeMux I__2162 (
            .O(N__9693),
            .I(N__9690));
    InMux I__2161 (
            .O(N__9690),
            .I(N__9687));
    LocalMux I__2160 (
            .O(N__9687),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    InMux I__2159 (
            .O(N__9684),
            .I(N__9681));
    LocalMux I__2158 (
            .O(N__9681),
            .I(N__9677));
    InMux I__2157 (
            .O(N__9680),
            .I(N__9674));
    Odrv4 I__2156 (
            .O(N__9677),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__2155 (
            .O(N__9674),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    InMux I__2154 (
            .O(N__9669),
            .I(N__9660));
    InMux I__2153 (
            .O(N__9668),
            .I(N__9660));
    InMux I__2152 (
            .O(N__9667),
            .I(N__9660));
    LocalMux I__2151 (
            .O(N__9660),
            .I(N__9657));
    Odrv4 I__2150 (
            .O(N__9657),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__2149 (
            .O(N__9654),
            .I(N__9651));
    LocalMux I__2148 (
            .O(N__9651),
            .I(N__9648));
    Odrv4 I__2147 (
            .O(N__9648),
            .I(\U712_REG_SM.N_402 ));
    IoInMux I__2146 (
            .O(N__9645),
            .I(N__9642));
    LocalMux I__2145 (
            .O(N__9642),
            .I(N__9639));
    Span12Mux_s0_v I__2144 (
            .O(N__9639),
            .I(N__9635));
    CascadeMux I__2143 (
            .O(N__9638),
            .I(N__9632));
    Span12Mux_h I__2142 (
            .O(N__9635),
            .I(N__9629));
    InMux I__2141 (
            .O(N__9632),
            .I(N__9626));
    Odrv12 I__2140 (
            .O(N__9629),
            .I(LDSn_c));
    LocalMux I__2139 (
            .O(N__9626),
            .I(LDSn_c));
    InMux I__2138 (
            .O(N__9621),
            .I(N__9614));
    CascadeMux I__2137 (
            .O(N__9620),
            .I(N__9610));
    CascadeMux I__2136 (
            .O(N__9619),
            .I(N__9607));
    CascadeMux I__2135 (
            .O(N__9618),
            .I(N__9602));
    InMux I__2134 (
            .O(N__9617),
            .I(N__9597));
    LocalMux I__2133 (
            .O(N__9614),
            .I(N__9594));
    InMux I__2132 (
            .O(N__9613),
            .I(N__9588));
    InMux I__2131 (
            .O(N__9610),
            .I(N__9583));
    InMux I__2130 (
            .O(N__9607),
            .I(N__9583));
    InMux I__2129 (
            .O(N__9606),
            .I(N__9578));
    InMux I__2128 (
            .O(N__9605),
            .I(N__9578));
    InMux I__2127 (
            .O(N__9602),
            .I(N__9574));
    InMux I__2126 (
            .O(N__9601),
            .I(N__9569));
    InMux I__2125 (
            .O(N__9600),
            .I(N__9569));
    LocalMux I__2124 (
            .O(N__9597),
            .I(N__9564));
    Span4Mux_h I__2123 (
            .O(N__9594),
            .I(N__9564));
    InMux I__2122 (
            .O(N__9593),
            .I(N__9557));
    InMux I__2121 (
            .O(N__9592),
            .I(N__9557));
    InMux I__2120 (
            .O(N__9591),
            .I(N__9557));
    LocalMux I__2119 (
            .O(N__9588),
            .I(N__9550));
    LocalMux I__2118 (
            .O(N__9583),
            .I(N__9550));
    LocalMux I__2117 (
            .O(N__9578),
            .I(N__9550));
    InMux I__2116 (
            .O(N__9577),
            .I(N__9547));
    LocalMux I__2115 (
            .O(N__9574),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__2114 (
            .O(N__9569),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__2113 (
            .O(N__9564),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__2112 (
            .O(N__9557),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__2111 (
            .O(N__9550),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__2110 (
            .O(N__9547),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    CascadeMux I__2109 (
            .O(N__9534),
            .I(N__9530));
    InMux I__2108 (
            .O(N__9533),
            .I(N__9524));
    InMux I__2107 (
            .O(N__9530),
            .I(N__9524));
    InMux I__2106 (
            .O(N__9529),
            .I(N__9521));
    LocalMux I__2105 (
            .O(N__9524),
            .I(N__9518));
    LocalMux I__2104 (
            .O(N__9521),
            .I(N__9515));
    Odrv4 I__2103 (
            .O(N__9518),
            .I(\U712_REG_SM.un1_REGENn_0_sqmuxa_0 ));
    Odrv4 I__2102 (
            .O(N__9515),
            .I(\U712_REG_SM.un1_REGENn_0_sqmuxa_0 ));
    IoInMux I__2101 (
            .O(N__9510),
            .I(N__9507));
    LocalMux I__2100 (
            .O(N__9507),
            .I(N__9504));
    Span4Mux_s2_v I__2099 (
            .O(N__9504),
            .I(N__9501));
    Span4Mux_v I__2098 (
            .O(N__9501),
            .I(N__9498));
    Span4Mux_v I__2097 (
            .O(N__9498),
            .I(N__9495));
    Sp12to4 I__2096 (
            .O(N__9495),
            .I(N__9491));
    InMux I__2095 (
            .O(N__9494),
            .I(N__9488));
    Odrv12 I__2094 (
            .O(N__9491),
            .I(UDSn_c));
    LocalMux I__2093 (
            .O(N__9488),
            .I(UDSn_c));
    IoInMux I__2092 (
            .O(N__9483),
            .I(N__9480));
    LocalMux I__2091 (
            .O(N__9480),
            .I(N__9477));
    Span4Mux_s0_v I__2090 (
            .O(N__9477),
            .I(N__9474));
    Span4Mux_v I__2089 (
            .O(N__9474),
            .I(N__9471));
    Odrv4 I__2088 (
            .O(N__9471),
            .I(RESETn_c_i));
    IoInMux I__2087 (
            .O(N__9468),
            .I(N__9465));
    LocalMux I__2086 (
            .O(N__9465),
            .I(N__9462));
    Span12Mux_s6_v I__2085 (
            .O(N__9462),
            .I(N__9459));
    Odrv12 I__2084 (
            .O(N__9459),
            .I(N_166));
    InMux I__2083 (
            .O(N__9456),
            .I(N__9443));
    InMux I__2082 (
            .O(N__9455),
            .I(N__9425));
    InMux I__2081 (
            .O(N__9454),
            .I(N__9425));
    InMux I__2080 (
            .O(N__9453),
            .I(N__9425));
    InMux I__2079 (
            .O(N__9452),
            .I(N__9425));
    InMux I__2078 (
            .O(N__9451),
            .I(N__9425));
    InMux I__2077 (
            .O(N__9450),
            .I(N__9425));
    InMux I__2076 (
            .O(N__9449),
            .I(N__9420));
    InMux I__2075 (
            .O(N__9448),
            .I(N__9420));
    CascadeMux I__2074 (
            .O(N__9447),
            .I(N__9414));
    CascadeMux I__2073 (
            .O(N__9446),
            .I(N__9411));
    LocalMux I__2072 (
            .O(N__9443),
            .I(N__9403));
    InMux I__2071 (
            .O(N__9442),
            .I(N__9400));
    InMux I__2070 (
            .O(N__9441),
            .I(N__9391));
    InMux I__2069 (
            .O(N__9440),
            .I(N__9391));
    InMux I__2068 (
            .O(N__9439),
            .I(N__9391));
    InMux I__2067 (
            .O(N__9438),
            .I(N__9391));
    LocalMux I__2066 (
            .O(N__9425),
            .I(N__9386));
    LocalMux I__2065 (
            .O(N__9420),
            .I(N__9386));
    InMux I__2064 (
            .O(N__9419),
            .I(N__9381));
    InMux I__2063 (
            .O(N__9418),
            .I(N__9381));
    InMux I__2062 (
            .O(N__9417),
            .I(N__9378));
    InMux I__2061 (
            .O(N__9414),
            .I(N__9375));
    InMux I__2060 (
            .O(N__9411),
            .I(N__9372));
    CascadeMux I__2059 (
            .O(N__9410),
            .I(N__9369));
    CascadeMux I__2058 (
            .O(N__9409),
            .I(N__9366));
    CascadeMux I__2057 (
            .O(N__9408),
            .I(N__9363));
    CascadeMux I__2056 (
            .O(N__9407),
            .I(N__9360));
    InMux I__2055 (
            .O(N__9406),
            .I(N__9357));
    Span4Mux_v I__2054 (
            .O(N__9403),
            .I(N__9345));
    LocalMux I__2053 (
            .O(N__9400),
            .I(N__9345));
    LocalMux I__2052 (
            .O(N__9391),
            .I(N__9345));
    Span4Mux_v I__2051 (
            .O(N__9386),
            .I(N__9345));
    LocalMux I__2050 (
            .O(N__9381),
            .I(N__9345));
    LocalMux I__2049 (
            .O(N__9378),
            .I(N__9339));
    LocalMux I__2048 (
            .O(N__9375),
            .I(N__9339));
    LocalMux I__2047 (
            .O(N__9372),
            .I(N__9336));
    InMux I__2046 (
            .O(N__9369),
            .I(N__9333));
    InMux I__2045 (
            .O(N__9366),
            .I(N__9330));
    InMux I__2044 (
            .O(N__9363),
            .I(N__9327));
    InMux I__2043 (
            .O(N__9360),
            .I(N__9324));
    LocalMux I__2042 (
            .O(N__9357),
            .I(N__9321));
    InMux I__2041 (
            .O(N__9356),
            .I(N__9318));
    Span4Mux_h I__2040 (
            .O(N__9345),
            .I(N__9315));
    InMux I__2039 (
            .O(N__9344),
            .I(N__9312));
    Span4Mux_h I__2038 (
            .O(N__9339),
            .I(N__9303));
    Span4Mux_h I__2037 (
            .O(N__9336),
            .I(N__9303));
    LocalMux I__2036 (
            .O(N__9333),
            .I(N__9303));
    LocalMux I__2035 (
            .O(N__9330),
            .I(N__9303));
    LocalMux I__2034 (
            .O(N__9327),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2033 (
            .O(N__9324),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__2032 (
            .O(N__9321),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2031 (
            .O(N__9318),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2030 (
            .O(N__9315),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2029 (
            .O(N__9312),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2028 (
            .O(N__9303),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    IoInMux I__2027 (
            .O(N__9288),
            .I(N__9285));
    LocalMux I__2026 (
            .O(N__9285),
            .I(N__9282));
    Span4Mux_s2_v I__2025 (
            .O(N__9282),
            .I(N__9279));
    Span4Mux_h I__2024 (
            .O(N__9279),
            .I(N__9276));
    Sp12to4 I__2023 (
            .O(N__9276),
            .I(N__9273));
    Span12Mux_s11_v I__2022 (
            .O(N__9273),
            .I(N__9270));
    Odrv12 I__2021 (
            .O(N__9270),
            .I(CASn_c));
    InMux I__2020 (
            .O(N__9267),
            .I(N__9264));
    LocalMux I__2019 (
            .O(N__9264),
            .I(N__9261));
    Span4Mux_v I__2018 (
            .O(N__9261),
            .I(N__9258));
    Odrv4 I__2017 (
            .O(N__9258),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2016 (
            .O(N__9255),
            .I(N__9252));
    LocalMux I__2015 (
            .O(N__9252),
            .I(N__9249));
    Odrv4 I__2014 (
            .O(N__9249),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2013 (
            .O(N__9246),
            .I(N__9243));
    LocalMux I__2012 (
            .O(N__9243),
            .I(N__9240));
    Odrv4 I__2011 (
            .O(N__9240),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2010 (
            .O(N__9237),
            .I(N__9229));
    InMux I__2009 (
            .O(N__9236),
            .I(N__9229));
    InMux I__2008 (
            .O(N__9235),
            .I(N__9223));
    InMux I__2007 (
            .O(N__9234),
            .I(N__9223));
    LocalMux I__2006 (
            .O(N__9229),
            .I(N__9220));
    InMux I__2005 (
            .O(N__9228),
            .I(N__9217));
    LocalMux I__2004 (
            .O(N__9223),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    Odrv4 I__2003 (
            .O(N__9220),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__2002 (
            .O(N__9217),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    CascadeMux I__2001 (
            .O(N__9210),
            .I(N__9206));
    InMux I__2000 (
            .O(N__9209),
            .I(N__9201));
    InMux I__1999 (
            .O(N__9206),
            .I(N__9201));
    LocalMux I__1998 (
            .O(N__9201),
            .I(N__9189));
    InMux I__1997 (
            .O(N__9200),
            .I(N__9182));
    InMux I__1996 (
            .O(N__9199),
            .I(N__9182));
    InMux I__1995 (
            .O(N__9198),
            .I(N__9182));
    InMux I__1994 (
            .O(N__9197),
            .I(N__9174));
    InMux I__1993 (
            .O(N__9196),
            .I(N__9174));
    InMux I__1992 (
            .O(N__9195),
            .I(N__9174));
    InMux I__1991 (
            .O(N__9194),
            .I(N__9167));
    InMux I__1990 (
            .O(N__9193),
            .I(N__9167));
    InMux I__1989 (
            .O(N__9192),
            .I(N__9167));
    Span4Mux_v I__1988 (
            .O(N__9189),
            .I(N__9164));
    LocalMux I__1987 (
            .O(N__9182),
            .I(N__9161));
    InMux I__1986 (
            .O(N__9181),
            .I(N__9158));
    LocalMux I__1985 (
            .O(N__9174),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1984 (
            .O(N__9167),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1983 (
            .O(N__9164),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1982 (
            .O(N__9161),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1981 (
            .O(N__9158),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    CascadeMux I__1980 (
            .O(N__9147),
            .I(N__9140));
    CascadeMux I__1979 (
            .O(N__9146),
            .I(N__9136));
    InMux I__1978 (
            .O(N__9145),
            .I(N__9133));
    InMux I__1977 (
            .O(N__9144),
            .I(N__9130));
    InMux I__1976 (
            .O(N__9143),
            .I(N__9127));
    InMux I__1975 (
            .O(N__9140),
            .I(N__9122));
    InMux I__1974 (
            .O(N__9139),
            .I(N__9122));
    InMux I__1973 (
            .O(N__9136),
            .I(N__9119));
    LocalMux I__1972 (
            .O(N__9133),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__1971 (
            .O(N__9130),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__1970 (
            .O(N__9127),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__1969 (
            .O(N__9122),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__1968 (
            .O(N__9119),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    CascadeMux I__1967 (
            .O(N__9108),
            .I(\U712_CYCLE_TERM.N_452_cascade_ ));
    CascadeMux I__1966 (
            .O(N__9105),
            .I(N__9102));
    InMux I__1965 (
            .O(N__9102),
            .I(N__9098));
    InMux I__1964 (
            .O(N__9101),
            .I(N__9093));
    LocalMux I__1963 (
            .O(N__9098),
            .I(N__9090));
    InMux I__1962 (
            .O(N__9097),
            .I(N__9087));
    InMux I__1961 (
            .O(N__9096),
            .I(N__9084));
    LocalMux I__1960 (
            .O(N__9093),
            .I(N__9081));
    Span4Mux_v I__1959 (
            .O(N__9090),
            .I(N__9078));
    LocalMux I__1958 (
            .O(N__9087),
            .I(N__9071));
    LocalMux I__1957 (
            .O(N__9084),
            .I(N__9071));
    Span4Mux_h I__1956 (
            .O(N__9081),
            .I(N__9071));
    Sp12to4 I__1955 (
            .O(N__9078),
            .I(N__9068));
    Sp12to4 I__1954 (
            .O(N__9071),
            .I(N__9063));
    Span12Mux_h I__1953 (
            .O(N__9068),
            .I(N__9063));
    Span12Mux_v I__1952 (
            .O(N__9063),
            .I(N__9060));
    Odrv12 I__1951 (
            .O(N__9060),
            .I(CLK40_PLL_i));
    CascadeMux I__1950 (
            .O(N__9057),
            .I(N__9052));
    CascadeMux I__1949 (
            .O(N__9056),
            .I(N__9048));
    CascadeMux I__1948 (
            .O(N__9055),
            .I(N__9040));
    InMux I__1947 (
            .O(N__9052),
            .I(N__9029));
    InMux I__1946 (
            .O(N__9051),
            .I(N__9029));
    InMux I__1945 (
            .O(N__9048),
            .I(N__9026));
    InMux I__1944 (
            .O(N__9047),
            .I(N__9018));
    InMux I__1943 (
            .O(N__9046),
            .I(N__9018));
    InMux I__1942 (
            .O(N__9045),
            .I(N__9018));
    InMux I__1941 (
            .O(N__9044),
            .I(N__9013));
    InMux I__1940 (
            .O(N__9043),
            .I(N__9013));
    InMux I__1939 (
            .O(N__9040),
            .I(N__9008));
    InMux I__1938 (
            .O(N__9039),
            .I(N__9005));
    InMux I__1937 (
            .O(N__9038),
            .I(N__8996));
    InMux I__1936 (
            .O(N__9037),
            .I(N__8996));
    InMux I__1935 (
            .O(N__9036),
            .I(N__8996));
    InMux I__1934 (
            .O(N__9035),
            .I(N__8991));
    InMux I__1933 (
            .O(N__9034),
            .I(N__8991));
    LocalMux I__1932 (
            .O(N__9029),
            .I(N__8987));
    LocalMux I__1931 (
            .O(N__9026),
            .I(N__8984));
    InMux I__1930 (
            .O(N__9025),
            .I(N__8981));
    LocalMux I__1929 (
            .O(N__9018),
            .I(N__8978));
    LocalMux I__1928 (
            .O(N__9013),
            .I(N__8975));
    InMux I__1927 (
            .O(N__9012),
            .I(N__8970));
    InMux I__1926 (
            .O(N__9011),
            .I(N__8970));
    LocalMux I__1925 (
            .O(N__9008),
            .I(N__8967));
    LocalMux I__1924 (
            .O(N__9005),
            .I(N__8964));
    InMux I__1923 (
            .O(N__9004),
            .I(N__8959));
    InMux I__1922 (
            .O(N__9003),
            .I(N__8959));
    LocalMux I__1921 (
            .O(N__8996),
            .I(N__8954));
    LocalMux I__1920 (
            .O(N__8991),
            .I(N__8954));
    InMux I__1919 (
            .O(N__8990),
            .I(N__8951));
    Span4Mux_v I__1918 (
            .O(N__8987),
            .I(N__8948));
    Span4Mux_h I__1917 (
            .O(N__8984),
            .I(N__8945));
    LocalMux I__1916 (
            .O(N__8981),
            .I(N__8940));
    Span4Mux_h I__1915 (
            .O(N__8978),
            .I(N__8940));
    Span4Mux_h I__1914 (
            .O(N__8975),
            .I(N__8937));
    LocalMux I__1913 (
            .O(N__8970),
            .I(N__8931));
    Span4Mux_v I__1912 (
            .O(N__8967),
            .I(N__8922));
    Span4Mux_h I__1911 (
            .O(N__8964),
            .I(N__8922));
    LocalMux I__1910 (
            .O(N__8959),
            .I(N__8922));
    Span4Mux_v I__1909 (
            .O(N__8954),
            .I(N__8922));
    LocalMux I__1908 (
            .O(N__8951),
            .I(N__8919));
    Span4Mux_h I__1907 (
            .O(N__8948),
            .I(N__8914));
    Span4Mux_v I__1906 (
            .O(N__8945),
            .I(N__8914));
    Span4Mux_h I__1905 (
            .O(N__8940),
            .I(N__8911));
    Span4Mux_h I__1904 (
            .O(N__8937),
            .I(N__8908));
    InMux I__1903 (
            .O(N__8936),
            .I(N__8901));
    InMux I__1902 (
            .O(N__8935),
            .I(N__8901));
    InMux I__1901 (
            .O(N__8934),
            .I(N__8901));
    Span4Mux_h I__1900 (
            .O(N__8931),
            .I(N__8896));
    Span4Mux_h I__1899 (
            .O(N__8922),
            .I(N__8896));
    Odrv12 I__1898 (
            .O(N__8919),
            .I(CPU_CYCLEm));
    Odrv4 I__1897 (
            .O(N__8914),
            .I(CPU_CYCLEm));
    Odrv4 I__1896 (
            .O(N__8911),
            .I(CPU_CYCLEm));
    Odrv4 I__1895 (
            .O(N__8908),
            .I(CPU_CYCLEm));
    LocalMux I__1894 (
            .O(N__8901),
            .I(CPU_CYCLEm));
    Odrv4 I__1893 (
            .O(N__8896),
            .I(CPU_CYCLEm));
    CascadeMux I__1892 (
            .O(N__8883),
            .I(\U712_BYTE_ENABLE.N_421_cascade_ ));
    IoInMux I__1891 (
            .O(N__8880),
            .I(N__8877));
    LocalMux I__1890 (
            .O(N__8877),
            .I(N__8874));
    Span4Mux_s3_h I__1889 (
            .O(N__8874),
            .I(N__8871));
    Span4Mux_v I__1888 (
            .O(N__8871),
            .I(N__8868));
    Sp12to4 I__1887 (
            .O(N__8868),
            .I(N__8865));
    Span12Mux_h I__1886 (
            .O(N__8865),
            .I(N__8862));
    Odrv12 I__1885 (
            .O(N__8862),
            .I(N_168_i));
    InMux I__1884 (
            .O(N__8859),
            .I(N__8856));
    LocalMux I__1883 (
            .O(N__8856),
            .I(\U712_CYCLE_TERM.N_326 ));
    CascadeMux I__1882 (
            .O(N__8853),
            .I(N__8850));
    InMux I__1881 (
            .O(N__8850),
            .I(N__8844));
    InMux I__1880 (
            .O(N__8849),
            .I(N__8841));
    InMux I__1879 (
            .O(N__8848),
            .I(N__8838));
    CascadeMux I__1878 (
            .O(N__8847),
            .I(N__8835));
    LocalMux I__1877 (
            .O(N__8844),
            .I(N__8830));
    LocalMux I__1876 (
            .O(N__8841),
            .I(N__8830));
    LocalMux I__1875 (
            .O(N__8838),
            .I(N__8827));
    InMux I__1874 (
            .O(N__8835),
            .I(N__8824));
    Span4Mux_h I__1873 (
            .O(N__8830),
            .I(N__8819));
    Span4Mux_v I__1872 (
            .O(N__8827),
            .I(N__8819));
    LocalMux I__1871 (
            .O(N__8824),
            .I(REG_TACK));
    Odrv4 I__1870 (
            .O(N__8819),
            .I(REG_TACK));
    InMux I__1869 (
            .O(N__8814),
            .I(N__8807));
    InMux I__1868 (
            .O(N__8813),
            .I(N__8807));
    InMux I__1867 (
            .O(N__8812),
            .I(N__8804));
    LocalMux I__1866 (
            .O(N__8807),
            .I(N__8798));
    LocalMux I__1865 (
            .O(N__8804),
            .I(N__8798));
    InMux I__1864 (
            .O(N__8803),
            .I(N__8795));
    Span12Mux_v I__1863 (
            .O(N__8798),
            .I(N__8792));
    LocalMux I__1862 (
            .O(N__8795),
            .I(CPU_TACKm));
    Odrv12 I__1861 (
            .O(N__8792),
            .I(CPU_TACKm));
    IoInMux I__1860 (
            .O(N__8787),
            .I(N__8784));
    LocalMux I__1859 (
            .O(N__8784),
            .I(N__8781));
    Span4Mux_s1_v I__1858 (
            .O(N__8781),
            .I(N__8775));
    InMux I__1857 (
            .O(N__8780),
            .I(N__8772));
    InMux I__1856 (
            .O(N__8779),
            .I(N__8767));
    InMux I__1855 (
            .O(N__8778),
            .I(N__8767));
    Sp12to4 I__1854 (
            .O(N__8775),
            .I(N__8763));
    LocalMux I__1853 (
            .O(N__8772),
            .I(N__8758));
    LocalMux I__1852 (
            .O(N__8767),
            .I(N__8758));
    InMux I__1851 (
            .O(N__8766),
            .I(N__8755));
    Span12Mux_h I__1850 (
            .O(N__8763),
            .I(N__8752));
    Span4Mux_v I__1849 (
            .O(N__8758),
            .I(N__8749));
    LocalMux I__1848 (
            .O(N__8755),
            .I(N__8746));
    Span12Mux_v I__1847 (
            .O(N__8752),
            .I(N__8742));
    Span4Mux_v I__1846 (
            .O(N__8749),
            .I(N__8739));
    Span4Mux_v I__1845 (
            .O(N__8746),
            .I(N__8736));
    InMux I__1844 (
            .O(N__8745),
            .I(N__8733));
    Odrv12 I__1843 (
            .O(N__8742),
            .I(DBENn_c));
    Odrv4 I__1842 (
            .O(N__8739),
            .I(DBENn_c));
    Odrv4 I__1841 (
            .O(N__8736),
            .I(DBENn_c));
    LocalMux I__1840 (
            .O(N__8733),
            .I(DBENn_c));
    InMux I__1839 (
            .O(N__8724),
            .I(N__8717));
    InMux I__1838 (
            .O(N__8723),
            .I(N__8714));
    InMux I__1837 (
            .O(N__8722),
            .I(N__8709));
    InMux I__1836 (
            .O(N__8721),
            .I(N__8709));
    InMux I__1835 (
            .O(N__8720),
            .I(N__8705));
    LocalMux I__1834 (
            .O(N__8717),
            .I(N__8702));
    LocalMux I__1833 (
            .O(N__8714),
            .I(N__8697));
    LocalMux I__1832 (
            .O(N__8709),
            .I(N__8697));
    InMux I__1831 (
            .O(N__8708),
            .I(N__8694));
    LocalMux I__1830 (
            .O(N__8705),
            .I(N__8691));
    Span4Mux_v I__1829 (
            .O(N__8702),
            .I(N__8686));
    Span4Mux_v I__1828 (
            .O(N__8697),
            .I(N__8686));
    LocalMux I__1827 (
            .O(N__8694),
            .I(N__8683));
    Span4Mux_h I__1826 (
            .O(N__8691),
            .I(N__8680));
    Odrv4 I__1825 (
            .O(N__8686),
            .I(DMA_CYCLEm));
    Odrv12 I__1824 (
            .O(N__8683),
            .I(DMA_CYCLEm));
    Odrv4 I__1823 (
            .O(N__8680),
            .I(DMA_CYCLEm));
    CascadeMux I__1822 (
            .O(N__8673),
            .I(N__8670));
    InMux I__1821 (
            .O(N__8670),
            .I(N__8667));
    LocalMux I__1820 (
            .O(N__8667),
            .I(\U712_BYTE_ENABLE.N_425 ));
    CascadeMux I__1819 (
            .O(N__8664),
            .I(N__8660));
    InMux I__1818 (
            .O(N__8663),
            .I(N__8656));
    InMux I__1817 (
            .O(N__8660),
            .I(N__8653));
    InMux I__1816 (
            .O(N__8659),
            .I(N__8650));
    LocalMux I__1815 (
            .O(N__8656),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__1814 (
            .O(N__8653),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__1813 (
            .O(N__8650),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__1812 (
            .O(N__8643),
            .I(N__8640));
    LocalMux I__1811 (
            .O(N__8640),
            .I(N__8637));
    Span4Mux_h I__1810 (
            .O(N__8637),
            .I(N__8634));
    Odrv4 I__1809 (
            .O(N__8634),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    InMux I__1808 (
            .O(N__8631),
            .I(N__8628));
    LocalMux I__1807 (
            .O(N__8628),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    InMux I__1806 (
            .O(N__8625),
            .I(N__8622));
    LocalMux I__1805 (
            .O(N__8622),
            .I(N__8619));
    Odrv12 I__1804 (
            .O(N__8619),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ));
    IoInMux I__1803 (
            .O(N__8616),
            .I(N__8611));
    IoInMux I__1802 (
            .O(N__8615),
            .I(N__8608));
    IoInMux I__1801 (
            .O(N__8614),
            .I(N__8605));
    LocalMux I__1800 (
            .O(N__8611),
            .I(N__8602));
    LocalMux I__1799 (
            .O(N__8608),
            .I(N__8599));
    LocalMux I__1798 (
            .O(N__8605),
            .I(N__8596));
    Span4Mux_s2_v I__1797 (
            .O(N__8602),
            .I(N__8593));
    Span4Mux_s2_v I__1796 (
            .O(N__8599),
            .I(N__8590));
    Span4Mux_s3_h I__1795 (
            .O(N__8596),
            .I(N__8587));
    Sp12to4 I__1794 (
            .O(N__8593),
            .I(N__8582));
    Sp12to4 I__1793 (
            .O(N__8590),
            .I(N__8582));
    Sp12to4 I__1792 (
            .O(N__8587),
            .I(N__8579));
    Span12Mux_h I__1791 (
            .O(N__8582),
            .I(N__8576));
    Span12Mux_v I__1790 (
            .O(N__8579),
            .I(N__8573));
    Span12Mux_v I__1789 (
            .O(N__8576),
            .I(N__8570));
    Span12Mux_h I__1788 (
            .O(N__8573),
            .I(N__8567));
    Odrv12 I__1787 (
            .O(N__8570),
            .I(CLK40_PLL_i_i));
    Odrv12 I__1786 (
            .O(N__8567),
            .I(CLK40_PLL_i_i));
    IoInMux I__1785 (
            .O(N__8562),
            .I(N__8557));
    IoInMux I__1784 (
            .O(N__8561),
            .I(N__8554));
    IoInMux I__1783 (
            .O(N__8560),
            .I(N__8551));
    LocalMux I__1782 (
            .O(N__8557),
            .I(N__8548));
    LocalMux I__1781 (
            .O(N__8554),
            .I(N__8545));
    LocalMux I__1780 (
            .O(N__8551),
            .I(N__8542));
    IoSpan4Mux I__1779 (
            .O(N__8548),
            .I(N__8539));
    Span4Mux_s3_v I__1778 (
            .O(N__8545),
            .I(N__8536));
    Span4Mux_s3_h I__1777 (
            .O(N__8542),
            .I(N__8533));
    Sp12to4 I__1776 (
            .O(N__8539),
            .I(N__8530));
    Sp12to4 I__1775 (
            .O(N__8536),
            .I(N__8527));
    Sp12to4 I__1774 (
            .O(N__8533),
            .I(N__8524));
    Span12Mux_s7_v I__1773 (
            .O(N__8530),
            .I(N__8521));
    Span12Mux_h I__1772 (
            .O(N__8527),
            .I(N__8518));
    Span12Mux_v I__1771 (
            .O(N__8524),
            .I(N__8515));
    Span12Mux_h I__1770 (
            .O(N__8521),
            .I(N__8511));
    Span12Mux_v I__1769 (
            .O(N__8518),
            .I(N__8506));
    Span12Mux_h I__1768 (
            .O(N__8515),
            .I(N__8506));
    InMux I__1767 (
            .O(N__8514),
            .I(N__8503));
    Odrv12 I__1766 (
            .O(N__8511),
            .I(TACK_EN));
    Odrv12 I__1765 (
            .O(N__8506),
            .I(TACK_EN));
    LocalMux I__1764 (
            .O(N__8503),
            .I(TACK_EN));
    IoInMux I__1763 (
            .O(N__8496),
            .I(N__8493));
    LocalMux I__1762 (
            .O(N__8493),
            .I(N__8490));
    IoSpan4Mux I__1761 (
            .O(N__8490),
            .I(N__8487));
    IoSpan4Mux I__1760 (
            .O(N__8487),
            .I(N__8484));
    Span4Mux_s3_h I__1759 (
            .O(N__8484),
            .I(N__8481));
    Span4Mux_v I__1758 (
            .O(N__8481),
            .I(N__8478));
    Span4Mux_v I__1757 (
            .O(N__8478),
            .I(N__8474));
    InMux I__1756 (
            .O(N__8477),
            .I(N__8471));
    Sp12to4 I__1755 (
            .O(N__8474),
            .I(N__8468));
    LocalMux I__1754 (
            .O(N__8471),
            .I(N__8465));
    Span12Mux_h I__1753 (
            .O(N__8468),
            .I(N__8460));
    Span12Mux_v I__1752 (
            .O(N__8465),
            .I(N__8460));
    Span12Mux_h I__1751 (
            .O(N__8460),
            .I(N__8457));
    Odrv12 I__1750 (
            .O(N__8457),
            .I(C3_c));
    InMux I__1749 (
            .O(N__8454),
            .I(N__8451));
    LocalMux I__1748 (
            .O(N__8451),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__1747 (
            .O(N__8448),
            .I(N__8443));
    InMux I__1746 (
            .O(N__8447),
            .I(N__8440));
    InMux I__1745 (
            .O(N__8446),
            .I(N__8437));
    LocalMux I__1744 (
            .O(N__8443),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    LocalMux I__1743 (
            .O(N__8440),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    LocalMux I__1742 (
            .O(N__8437),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    InMux I__1741 (
            .O(N__8430),
            .I(N__8426));
    InMux I__1740 (
            .O(N__8429),
            .I(N__8423));
    LocalMux I__1739 (
            .O(N__8426),
            .I(\U712_REG_SM.START_RSTZ0 ));
    LocalMux I__1738 (
            .O(N__8423),
            .I(\U712_REG_SM.START_RSTZ0 ));
    CascadeMux I__1737 (
            .O(N__8418),
            .I(\U712_BYTE_ENABLE.N_443_cascade_ ));
    IoInMux I__1736 (
            .O(N__8415),
            .I(N__8412));
    LocalMux I__1735 (
            .O(N__8412),
            .I(N__8409));
    IoSpan4Mux I__1734 (
            .O(N__8409),
            .I(N__8406));
    Span4Mux_s2_h I__1733 (
            .O(N__8406),
            .I(N__8403));
    Sp12to4 I__1732 (
            .O(N__8403),
            .I(N__8400));
    Span12Mux_h I__1731 (
            .O(N__8400),
            .I(N__8397));
    Span12Mux_v I__1730 (
            .O(N__8397),
            .I(N__8394));
    Odrv12 I__1729 (
            .O(N__8394),
            .I(N_54_i));
    InMux I__1728 (
            .O(N__8391),
            .I(N__8385));
    InMux I__1727 (
            .O(N__8390),
            .I(N__8382));
    InMux I__1726 (
            .O(N__8389),
            .I(N__8379));
    CascadeMux I__1725 (
            .O(N__8388),
            .I(N__8370));
    LocalMux I__1724 (
            .O(N__8385),
            .I(N__8365));
    LocalMux I__1723 (
            .O(N__8382),
            .I(N__8365));
    LocalMux I__1722 (
            .O(N__8379),
            .I(N__8362));
    InMux I__1721 (
            .O(N__8378),
            .I(N__8359));
    InMux I__1720 (
            .O(N__8377),
            .I(N__8356));
    InMux I__1719 (
            .O(N__8376),
            .I(N__8351));
    InMux I__1718 (
            .O(N__8375),
            .I(N__8351));
    InMux I__1717 (
            .O(N__8374),
            .I(N__8346));
    InMux I__1716 (
            .O(N__8373),
            .I(N__8346));
    InMux I__1715 (
            .O(N__8370),
            .I(N__8343));
    Span4Mux_v I__1714 (
            .O(N__8365),
            .I(N__8340));
    Span4Mux_h I__1713 (
            .O(N__8362),
            .I(N__8337));
    LocalMux I__1712 (
            .O(N__8359),
            .I(\U712_CHIP_RAM.N_309 ));
    LocalMux I__1711 (
            .O(N__8356),
            .I(\U712_CHIP_RAM.N_309 ));
    LocalMux I__1710 (
            .O(N__8351),
            .I(\U712_CHIP_RAM.N_309 ));
    LocalMux I__1709 (
            .O(N__8346),
            .I(\U712_CHIP_RAM.N_309 ));
    LocalMux I__1708 (
            .O(N__8343),
            .I(\U712_CHIP_RAM.N_309 ));
    Odrv4 I__1707 (
            .O(N__8340),
            .I(\U712_CHIP_RAM.N_309 ));
    Odrv4 I__1706 (
            .O(N__8337),
            .I(\U712_CHIP_RAM.N_309 ));
    InMux I__1705 (
            .O(N__8322),
            .I(N__8319));
    LocalMux I__1704 (
            .O(N__8319),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    CascadeMux I__1703 (
            .O(N__8316),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1_cascade_ ));
    IoInMux I__1702 (
            .O(N__8313),
            .I(N__8310));
    LocalMux I__1701 (
            .O(N__8310),
            .I(N__8307));
    Span12Mux_s9_v I__1700 (
            .O(N__8307),
            .I(N__8304));
    Odrv12 I__1699 (
            .O(N__8304),
            .I(CMA_c_1));
    CEMux I__1698 (
            .O(N__8301),
            .I(N__8297));
    CEMux I__1697 (
            .O(N__8300),
            .I(N__8294));
    LocalMux I__1696 (
            .O(N__8297),
            .I(N__8287));
    LocalMux I__1695 (
            .O(N__8294),
            .I(N__8284));
    CEMux I__1694 (
            .O(N__8293),
            .I(N__8281));
    CEMux I__1693 (
            .O(N__8292),
            .I(N__8278));
    CEMux I__1692 (
            .O(N__8291),
            .I(N__8275));
    CEMux I__1691 (
            .O(N__8290),
            .I(N__8272));
    Span4Mux_v I__1690 (
            .O(N__8287),
            .I(N__8265));
    Span4Mux_h I__1689 (
            .O(N__8284),
            .I(N__8265));
    LocalMux I__1688 (
            .O(N__8281),
            .I(N__8265));
    LocalMux I__1687 (
            .O(N__8278),
            .I(N__8260));
    LocalMux I__1686 (
            .O(N__8275),
            .I(N__8260));
    LocalMux I__1685 (
            .O(N__8272),
            .I(N__8257));
    Span4Mux_h I__1684 (
            .O(N__8265),
            .I(N__8254));
    Span4Mux_v I__1683 (
            .O(N__8260),
            .I(N__8251));
    Span4Mux_v I__1682 (
            .O(N__8257),
            .I(N__8248));
    Odrv4 I__1681 (
            .O(N__8254),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv4 I__1680 (
            .O(N__8251),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv4 I__1679 (
            .O(N__8248),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    InMux I__1678 (
            .O(N__8241),
            .I(N__8238));
    LocalMux I__1677 (
            .O(N__8238),
            .I(N__8235));
    Span12Mux_v I__1676 (
            .O(N__8235),
            .I(N__8232));
    Span12Mux_h I__1675 (
            .O(N__8232),
            .I(N__8229));
    Odrv12 I__1674 (
            .O(N__8229),
            .I(A_c_15));
    InMux I__1673 (
            .O(N__8226),
            .I(N__8222));
    InMux I__1672 (
            .O(N__8225),
            .I(N__8219));
    LocalMux I__1671 (
            .O(N__8222),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ));
    LocalMux I__1670 (
            .O(N__8219),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ));
    CascadeMux I__1669 (
            .O(N__8214),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ));
    InMux I__1668 (
            .O(N__8211),
            .I(N__8208));
    LocalMux I__1667 (
            .O(N__8208),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__1666 (
            .O(N__8205),
            .I(N__8202));
    LocalMux I__1665 (
            .O(N__8202),
            .I(N__8199));
    IoSpan4Mux I__1664 (
            .O(N__8199),
            .I(N__8196));
    IoSpan4Mux I__1663 (
            .O(N__8196),
            .I(N__8192));
    InMux I__1662 (
            .O(N__8195),
            .I(N__8189));
    Span4Mux_s2_v I__1661 (
            .O(N__8192),
            .I(N__8186));
    LocalMux I__1660 (
            .O(N__8189),
            .I(N__8183));
    Sp12to4 I__1659 (
            .O(N__8186),
            .I(N__8180));
    Span4Mux_v I__1658 (
            .O(N__8183),
            .I(N__8177));
    Span12Mux_s8_v I__1657 (
            .O(N__8180),
            .I(N__8174));
    Sp12to4 I__1656 (
            .O(N__8177),
            .I(N__8171));
    Span12Mux_v I__1655 (
            .O(N__8174),
            .I(N__8166));
    Span12Mux_h I__1654 (
            .O(N__8171),
            .I(N__8166));
    Odrv12 I__1653 (
            .O(N__8166),
            .I(A_c_10));
    InMux I__1652 (
            .O(N__8163),
            .I(N__8159));
    InMux I__1651 (
            .O(N__8162),
            .I(N__8156));
    LocalMux I__1650 (
            .O(N__8159),
            .I(N__8153));
    LocalMux I__1649 (
            .O(N__8156),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ));
    Odrv4 I__1648 (
            .O(N__8153),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ));
    CascadeMux I__1647 (
            .O(N__8148),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ));
    InMux I__1646 (
            .O(N__8145),
            .I(N__8142));
    LocalMux I__1645 (
            .O(N__8142),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    InMux I__1644 (
            .O(N__8139),
            .I(N__8136));
    LocalMux I__1643 (
            .O(N__8136),
            .I(N__8133));
    Span12Mux_v I__1642 (
            .O(N__8133),
            .I(N__8130));
    Span12Mux_h I__1641 (
            .O(N__8130),
            .I(N__8127));
    Odrv12 I__1640 (
            .O(N__8127),
            .I(A_c_13));
    InMux I__1639 (
            .O(N__8124),
            .I(N__8120));
    InMux I__1638 (
            .O(N__8123),
            .I(N__8117));
    LocalMux I__1637 (
            .O(N__8120),
            .I(N__8114));
    LocalMux I__1636 (
            .O(N__8117),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ));
    Odrv4 I__1635 (
            .O(N__8114),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ));
    CascadeMux I__1634 (
            .O(N__8109),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ));
    InMux I__1633 (
            .O(N__8106),
            .I(N__8103));
    LocalMux I__1632 (
            .O(N__8103),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    InMux I__1631 (
            .O(N__8100),
            .I(N__8094));
    InMux I__1630 (
            .O(N__8099),
            .I(N__8094));
    LocalMux I__1629 (
            .O(N__8094),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    IoInMux I__1628 (
            .O(N__8091),
            .I(N__8088));
    LocalMux I__1627 (
            .O(N__8088),
            .I(N__8085));
    IoSpan4Mux I__1626 (
            .O(N__8085),
            .I(N__8082));
    IoSpan4Mux I__1625 (
            .O(N__8082),
            .I(N__8079));
    Span4Mux_s1_v I__1624 (
            .O(N__8079),
            .I(N__8076));
    Sp12to4 I__1623 (
            .O(N__8076),
            .I(N__8073));
    Span12Mux_s9_v I__1622 (
            .O(N__8073),
            .I(N__8070));
    Odrv12 I__1621 (
            .O(N__8070),
            .I(ASn_c));
    CEMux I__1620 (
            .O(N__8067),
            .I(N__8064));
    LocalMux I__1619 (
            .O(N__8064),
            .I(N__8061));
    Span4Mux_h I__1618 (
            .O(N__8061),
            .I(N__8058));
    Odrv4 I__1617 (
            .O(N__8058),
            .I(\U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0 ));
    IoInMux I__1616 (
            .O(N__8055),
            .I(N__8052));
    LocalMux I__1615 (
            .O(N__8052),
            .I(N__8049));
    Span4Mux_s3_v I__1614 (
            .O(N__8049),
            .I(N__8046));
    Span4Mux_h I__1613 (
            .O(N__8046),
            .I(N__8043));
    Span4Mux_h I__1612 (
            .O(N__8043),
            .I(N__8040));
    Odrv4 I__1611 (
            .O(N__8040),
            .I(RASn_c));
    InMux I__1610 (
            .O(N__8037),
            .I(N__8034));
    LocalMux I__1609 (
            .O(N__8034),
            .I(N__8031));
    Odrv12 I__1608 (
            .O(N__8031),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__1607 (
            .O(N__8028),
            .I(N__8025));
    LocalMux I__1606 (
            .O(N__8025),
            .I(N__8022));
    Odrv12 I__1605 (
            .O(N__8022),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    InMux I__1604 (
            .O(N__8019),
            .I(N__8016));
    LocalMux I__1603 (
            .O(N__8016),
            .I(N__8013));
    Span4Mux_h I__1602 (
            .O(N__8013),
            .I(N__8007));
    InMux I__1601 (
            .O(N__8012),
            .I(N__8004));
    InMux I__1600 (
            .O(N__8011),
            .I(N__8001));
    InMux I__1599 (
            .O(N__8010),
            .I(N__7998));
    Span4Mux_v I__1598 (
            .O(N__8007),
            .I(N__7991));
    LocalMux I__1597 (
            .O(N__8004),
            .I(N__7991));
    LocalMux I__1596 (
            .O(N__8001),
            .I(N__7986));
    LocalMux I__1595 (
            .O(N__7998),
            .I(N__7986));
    InMux I__1594 (
            .O(N__7997),
            .I(N__7983));
    InMux I__1593 (
            .O(N__7996),
            .I(N__7980));
    Odrv4 I__1592 (
            .O(N__7991),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv12 I__1591 (
            .O(N__7986),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1590 (
            .O(N__7983),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1589 (
            .O(N__7980),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    CascadeMux I__1588 (
            .O(N__7971),
            .I(\U712_CHIP_RAM.N_309_cascade_ ));
    CascadeMux I__1587 (
            .O(N__7968),
            .I(\U712_REG_SM.N_325_cascade_ ));
    InMux I__1586 (
            .O(N__7965),
            .I(N__7962));
    LocalMux I__1585 (
            .O(N__7962),
            .I(\U712_REG_SM.N_302 ));
    CascadeMux I__1584 (
            .O(N__7959),
            .I(\U712_REG_SM.N_302_cascade_ ));
    InMux I__1583 (
            .O(N__7956),
            .I(N__7953));
    LocalMux I__1582 (
            .O(N__7953),
            .I(N__7950));
    Span4Mux_v I__1581 (
            .O(N__7950),
            .I(N__7945));
    InMux I__1580 (
            .O(N__7949),
            .I(N__7942));
    InMux I__1579 (
            .O(N__7948),
            .I(N__7939));
    Odrv4 I__1578 (
            .O(N__7945),
            .I(REG_CYCLEm));
    LocalMux I__1577 (
            .O(N__7942),
            .I(REG_CYCLEm));
    LocalMux I__1576 (
            .O(N__7939),
            .I(REG_CYCLEm));
    IoInMux I__1575 (
            .O(N__7932),
            .I(N__7929));
    LocalMux I__1574 (
            .O(N__7929),
            .I(N__7926));
    IoSpan4Mux I__1573 (
            .O(N__7926),
            .I(N__7923));
    IoSpan4Mux I__1572 (
            .O(N__7923),
            .I(N__7920));
    Sp12to4 I__1571 (
            .O(N__7920),
            .I(N__7917));
    Span12Mux_v I__1570 (
            .O(N__7917),
            .I(N__7914));
    Odrv12 I__1569 (
            .O(N__7914),
            .I(N_160_i));
    CascadeMux I__1568 (
            .O(N__7911),
            .I(N__7906));
    InMux I__1567 (
            .O(N__7910),
            .I(N__7898));
    InMux I__1566 (
            .O(N__7909),
            .I(N__7898));
    InMux I__1565 (
            .O(N__7906),
            .I(N__7895));
    InMux I__1564 (
            .O(N__7905),
            .I(N__7892));
    InMux I__1563 (
            .O(N__7904),
            .I(N__7887));
    InMux I__1562 (
            .O(N__7903),
            .I(N__7887));
    LocalMux I__1561 (
            .O(N__7898),
            .I(N__7884));
    LocalMux I__1560 (
            .O(N__7895),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1559 (
            .O(N__7892),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1558 (
            .O(N__7887),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv12 I__1557 (
            .O(N__7884),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    InMux I__1556 (
            .O(N__7875),
            .I(N__7872));
    LocalMux I__1555 (
            .O(N__7872),
            .I(\U712_REG_SM.N_404 ));
    IoInMux I__1554 (
            .O(N__7869),
            .I(N__7865));
    IoInMux I__1553 (
            .O(N__7868),
            .I(N__7862));
    LocalMux I__1552 (
            .O(N__7865),
            .I(N__7858));
    LocalMux I__1551 (
            .O(N__7862),
            .I(N__7855));
    IoInMux I__1550 (
            .O(N__7861),
            .I(N__7852));
    Span4Mux_s3_v I__1549 (
            .O(N__7858),
            .I(N__7849));
    Span4Mux_s1_v I__1548 (
            .O(N__7855),
            .I(N__7846));
    LocalMux I__1547 (
            .O(N__7852),
            .I(N__7843));
    Span4Mux_v I__1546 (
            .O(N__7849),
            .I(N__7840));
    Span4Mux_v I__1545 (
            .O(N__7846),
            .I(N__7837));
    Span4Mux_s2_h I__1544 (
            .O(N__7843),
            .I(N__7834));
    Span4Mux_h I__1543 (
            .O(N__7840),
            .I(N__7831));
    Sp12to4 I__1542 (
            .O(N__7837),
            .I(N__7828));
    Sp12to4 I__1541 (
            .O(N__7834),
            .I(N__7825));
    Sp12to4 I__1540 (
            .O(N__7831),
            .I(N__7822));
    Span12Mux_h I__1539 (
            .O(N__7828),
            .I(N__7819));
    Span12Mux_v I__1538 (
            .O(N__7825),
            .I(N__7816));
    Span12Mux_v I__1537 (
            .O(N__7822),
            .I(N__7812));
    Span12Mux_v I__1536 (
            .O(N__7819),
            .I(N__7807));
    Span12Mux_h I__1535 (
            .O(N__7816),
            .I(N__7807));
    InMux I__1534 (
            .O(N__7815),
            .I(N__7804));
    Odrv12 I__1533 (
            .O(N__7812),
            .I(TACK_OUTn));
    Odrv12 I__1532 (
            .O(N__7807),
            .I(TACK_OUTn));
    LocalMux I__1531 (
            .O(N__7804),
            .I(TACK_OUTn));
    InMux I__1530 (
            .O(N__7797),
            .I(N__7793));
    IoInMux I__1529 (
            .O(N__7796),
            .I(N__7790));
    LocalMux I__1528 (
            .O(N__7793),
            .I(N__7787));
    LocalMux I__1527 (
            .O(N__7790),
            .I(N__7784));
    Sp12to4 I__1526 (
            .O(N__7787),
            .I(N__7781));
    IoSpan4Mux I__1525 (
            .O(N__7784),
            .I(N__7778));
    Span12Mux_v I__1524 (
            .O(N__7781),
            .I(N__7775));
    IoSpan4Mux I__1523 (
            .O(N__7778),
            .I(N__7772));
    Span12Mux_h I__1522 (
            .O(N__7775),
            .I(N__7769));
    IoSpan4Mux I__1521 (
            .O(N__7772),
            .I(N__7766));
    Odrv12 I__1520 (
            .O(N__7769),
            .I(C1_c));
    Odrv4 I__1519 (
            .O(N__7766),
            .I(C1_c));
    InMux I__1518 (
            .O(N__7761),
            .I(N__7758));
    LocalMux I__1517 (
            .O(N__7758),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__1516 (
            .O(N__7755),
            .I(N__7750));
    InMux I__1515 (
            .O(N__7754),
            .I(N__7747));
    InMux I__1514 (
            .O(N__7753),
            .I(N__7734));
    LocalMux I__1513 (
            .O(N__7750),
            .I(N__7731));
    LocalMux I__1512 (
            .O(N__7747),
            .I(N__7727));
    InMux I__1511 (
            .O(N__7746),
            .I(N__7720));
    InMux I__1510 (
            .O(N__7745),
            .I(N__7720));
    InMux I__1509 (
            .O(N__7744),
            .I(N__7720));
    InMux I__1508 (
            .O(N__7743),
            .I(N__7714));
    InMux I__1507 (
            .O(N__7742),
            .I(N__7714));
    InMux I__1506 (
            .O(N__7741),
            .I(N__7711));
    InMux I__1505 (
            .O(N__7740),
            .I(N__7702));
    InMux I__1504 (
            .O(N__7739),
            .I(N__7702));
    CascadeMux I__1503 (
            .O(N__7738),
            .I(N__7699));
    InMux I__1502 (
            .O(N__7737),
            .I(N__7688));
    LocalMux I__1501 (
            .O(N__7734),
            .I(N__7685));
    Span4Mux_h I__1500 (
            .O(N__7731),
            .I(N__7682));
    InMux I__1499 (
            .O(N__7730),
            .I(N__7679));
    Span4Mux_h I__1498 (
            .O(N__7727),
            .I(N__7674));
    LocalMux I__1497 (
            .O(N__7720),
            .I(N__7674));
    InMux I__1496 (
            .O(N__7719),
            .I(N__7671));
    LocalMux I__1495 (
            .O(N__7714),
            .I(N__7666));
    LocalMux I__1494 (
            .O(N__7711),
            .I(N__7666));
    InMux I__1493 (
            .O(N__7710),
            .I(N__7661));
    InMux I__1492 (
            .O(N__7709),
            .I(N__7661));
    InMux I__1491 (
            .O(N__7708),
            .I(N__7656));
    InMux I__1490 (
            .O(N__7707),
            .I(N__7656));
    LocalMux I__1489 (
            .O(N__7702),
            .I(N__7653));
    InMux I__1488 (
            .O(N__7699),
            .I(N__7648));
    InMux I__1487 (
            .O(N__7698),
            .I(N__7648));
    InMux I__1486 (
            .O(N__7697),
            .I(N__7645));
    InMux I__1485 (
            .O(N__7696),
            .I(N__7640));
    InMux I__1484 (
            .O(N__7695),
            .I(N__7640));
    InMux I__1483 (
            .O(N__7694),
            .I(N__7633));
    InMux I__1482 (
            .O(N__7693),
            .I(N__7633));
    InMux I__1481 (
            .O(N__7692),
            .I(N__7633));
    InMux I__1480 (
            .O(N__7691),
            .I(N__7630));
    LocalMux I__1479 (
            .O(N__7688),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1478 (
            .O(N__7685),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1477 (
            .O(N__7682),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1476 (
            .O(N__7679),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1475 (
            .O(N__7674),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1474 (
            .O(N__7671),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv12 I__1473 (
            .O(N__7666),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1472 (
            .O(N__7661),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1471 (
            .O(N__7656),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1470 (
            .O(N__7653),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1469 (
            .O(N__7648),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1468 (
            .O(N__7645),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1467 (
            .O(N__7640),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1466 (
            .O(N__7633),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1465 (
            .O(N__7630),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1464 (
            .O(N__7599),
            .I(N__7587));
    InMux I__1463 (
            .O(N__7598),
            .I(N__7584));
    InMux I__1462 (
            .O(N__7597),
            .I(N__7575));
    InMux I__1461 (
            .O(N__7596),
            .I(N__7572));
    InMux I__1460 (
            .O(N__7595),
            .I(N__7569));
    InMux I__1459 (
            .O(N__7594),
            .I(N__7562));
    InMux I__1458 (
            .O(N__7593),
            .I(N__7562));
    InMux I__1457 (
            .O(N__7592),
            .I(N__7562));
    InMux I__1456 (
            .O(N__7591),
            .I(N__7557));
    InMux I__1455 (
            .O(N__7590),
            .I(N__7557));
    LocalMux I__1454 (
            .O(N__7587),
            .I(N__7553));
    LocalMux I__1453 (
            .O(N__7584),
            .I(N__7550));
    CascadeMux I__1452 (
            .O(N__7583),
            .I(N__7542));
    CascadeMux I__1451 (
            .O(N__7582),
            .I(N__7537));
    InMux I__1450 (
            .O(N__7581),
            .I(N__7534));
    InMux I__1449 (
            .O(N__7580),
            .I(N__7527));
    InMux I__1448 (
            .O(N__7579),
            .I(N__7527));
    InMux I__1447 (
            .O(N__7578),
            .I(N__7527));
    LocalMux I__1446 (
            .O(N__7575),
            .I(N__7524));
    LocalMux I__1445 (
            .O(N__7572),
            .I(N__7517));
    LocalMux I__1444 (
            .O(N__7569),
            .I(N__7517));
    LocalMux I__1443 (
            .O(N__7562),
            .I(N__7517));
    LocalMux I__1442 (
            .O(N__7557),
            .I(N__7514));
    InMux I__1441 (
            .O(N__7556),
            .I(N__7511));
    Span4Mux_h I__1440 (
            .O(N__7553),
            .I(N__7508));
    Span12Mux_v I__1439 (
            .O(N__7550),
            .I(N__7505));
    InMux I__1438 (
            .O(N__7549),
            .I(N__7500));
    InMux I__1437 (
            .O(N__7548),
            .I(N__7500));
    InMux I__1436 (
            .O(N__7547),
            .I(N__7495));
    InMux I__1435 (
            .O(N__7546),
            .I(N__7495));
    InMux I__1434 (
            .O(N__7545),
            .I(N__7490));
    InMux I__1433 (
            .O(N__7542),
            .I(N__7490));
    InMux I__1432 (
            .O(N__7541),
            .I(N__7483));
    InMux I__1431 (
            .O(N__7540),
            .I(N__7483));
    InMux I__1430 (
            .O(N__7537),
            .I(N__7483));
    LocalMux I__1429 (
            .O(N__7534),
            .I(N__7478));
    LocalMux I__1428 (
            .O(N__7527),
            .I(N__7478));
    Span4Mux_h I__1427 (
            .O(N__7524),
            .I(N__7471));
    Span4Mux_v I__1426 (
            .O(N__7517),
            .I(N__7471));
    Span4Mux_h I__1425 (
            .O(N__7514),
            .I(N__7471));
    LocalMux I__1424 (
            .O(N__7511),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1423 (
            .O(N__7508),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv12 I__1422 (
            .O(N__7505),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1421 (
            .O(N__7500),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1420 (
            .O(N__7495),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1419 (
            .O(N__7490),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1418 (
            .O(N__7483),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1417 (
            .O(N__7478),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1416 (
            .O(N__7471),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__1415 (
            .O(N__7452),
            .I(N__7447));
    CascadeMux I__1414 (
            .O(N__7451),
            .I(N__7444));
    CascadeMux I__1413 (
            .O(N__7450),
            .I(N__7440));
    InMux I__1412 (
            .O(N__7447),
            .I(N__7435));
    InMux I__1411 (
            .O(N__7444),
            .I(N__7432));
    CascadeMux I__1410 (
            .O(N__7443),
            .I(N__7429));
    InMux I__1409 (
            .O(N__7440),
            .I(N__7426));
    InMux I__1408 (
            .O(N__7439),
            .I(N__7420));
    InMux I__1407 (
            .O(N__7438),
            .I(N__7420));
    LocalMux I__1406 (
            .O(N__7435),
            .I(N__7415));
    LocalMux I__1405 (
            .O(N__7432),
            .I(N__7415));
    InMux I__1404 (
            .O(N__7429),
            .I(N__7412));
    LocalMux I__1403 (
            .O(N__7426),
            .I(N__7409));
    InMux I__1402 (
            .O(N__7425),
            .I(N__7405));
    LocalMux I__1401 (
            .O(N__7420),
            .I(N__7402));
    Span4Mux_h I__1400 (
            .O(N__7415),
            .I(N__7397));
    LocalMux I__1399 (
            .O(N__7412),
            .I(N__7397));
    Span4Mux_h I__1398 (
            .O(N__7409),
            .I(N__7394));
    InMux I__1397 (
            .O(N__7408),
            .I(N__7391));
    LocalMux I__1396 (
            .O(N__7405),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1395 (
            .O(N__7402),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1394 (
            .O(N__7397),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1393 (
            .O(N__7394),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1392 (
            .O(N__7391),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1391 (
            .O(N__7380),
            .I(N__7375));
    InMux I__1390 (
            .O(N__7379),
            .I(N__7372));
    InMux I__1389 (
            .O(N__7378),
            .I(N__7368));
    LocalMux I__1388 (
            .O(N__7375),
            .I(N__7364));
    LocalMux I__1387 (
            .O(N__7372),
            .I(N__7361));
    InMux I__1386 (
            .O(N__7371),
            .I(N__7358));
    LocalMux I__1385 (
            .O(N__7368),
            .I(N__7355));
    InMux I__1384 (
            .O(N__7367),
            .I(N__7352));
    Odrv4 I__1383 (
            .O(N__7364),
            .I(\U712_CHIP_RAM.N_466 ));
    Odrv4 I__1382 (
            .O(N__7361),
            .I(\U712_CHIP_RAM.N_466 ));
    LocalMux I__1381 (
            .O(N__7358),
            .I(\U712_CHIP_RAM.N_466 ));
    Odrv4 I__1380 (
            .O(N__7355),
            .I(\U712_CHIP_RAM.N_466 ));
    LocalMux I__1379 (
            .O(N__7352),
            .I(\U712_CHIP_RAM.N_466 ));
    CEMux I__1378 (
            .O(N__7341),
            .I(N__7338));
    LocalMux I__1377 (
            .O(N__7338),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0 ));
    InMux I__1376 (
            .O(N__7335),
            .I(N__7332));
    LocalMux I__1375 (
            .O(N__7332),
            .I(N__7329));
    Span4Mux_v I__1374 (
            .O(N__7329),
            .I(N__7326));
    Sp12to4 I__1373 (
            .O(N__7326),
            .I(N__7323));
    Span12Mux_h I__1372 (
            .O(N__7323),
            .I(N__7320));
    Span12Mux_v I__1371 (
            .O(N__7320),
            .I(N__7317));
    Odrv12 I__1370 (
            .O(N__7317),
            .I(REGSPACEn_c));
    InMux I__1369 (
            .O(N__7314),
            .I(N__7310));
    InMux I__1368 (
            .O(N__7313),
            .I(N__7307));
    LocalMux I__1367 (
            .O(N__7310),
            .I(N__7304));
    LocalMux I__1366 (
            .O(N__7307),
            .I(N__7301));
    Span4Mux_v I__1365 (
            .O(N__7304),
            .I(N__7298));
    Span4Mux_v I__1364 (
            .O(N__7301),
            .I(N__7295));
    Sp12to4 I__1363 (
            .O(N__7298),
            .I(N__7290));
    Sp12to4 I__1362 (
            .O(N__7295),
            .I(N__7290));
    Span12Mux_h I__1361 (
            .O(N__7290),
            .I(N__7287));
    Span12Mux_v I__1360 (
            .O(N__7287),
            .I(N__7284));
    Odrv12 I__1359 (
            .O(N__7284),
            .I(TSn_c));
    CascadeMux I__1358 (
            .O(N__7281),
            .I(\U712_REG_SM.N_401_cascade_ ));
    InMux I__1357 (
            .O(N__7278),
            .I(N__7271));
    InMux I__1356 (
            .O(N__7277),
            .I(N__7271));
    InMux I__1355 (
            .O(N__7276),
            .I(N__7267));
    LocalMux I__1354 (
            .O(N__7271),
            .I(N__7264));
    InMux I__1353 (
            .O(N__7270),
            .I(N__7261));
    LocalMux I__1352 (
            .O(N__7267),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    Odrv4 I__1351 (
            .O(N__7264),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1350 (
            .O(N__7261),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__1349 (
            .O(N__7254),
            .I(N__7250));
    InMux I__1348 (
            .O(N__7253),
            .I(N__7247));
    LocalMux I__1347 (
            .O(N__7250),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    LocalMux I__1346 (
            .O(N__7247),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    CascadeMux I__1345 (
            .O(N__7242),
            .I(N__7238));
    InMux I__1344 (
            .O(N__7241),
            .I(N__7233));
    InMux I__1343 (
            .O(N__7238),
            .I(N__7230));
    InMux I__1342 (
            .O(N__7237),
            .I(N__7227));
    InMux I__1341 (
            .O(N__7236),
            .I(N__7224));
    LocalMux I__1340 (
            .O(N__7233),
            .I(N__7221));
    LocalMux I__1339 (
            .O(N__7230),
            .I(N__7216));
    LocalMux I__1338 (
            .O(N__7227),
            .I(N__7216));
    LocalMux I__1337 (
            .O(N__7224),
            .I(N__7212));
    Span4Mux_h I__1336 (
            .O(N__7221),
            .I(N__7209));
    Span4Mux_h I__1335 (
            .O(N__7216),
            .I(N__7206));
    InMux I__1334 (
            .O(N__7215),
            .I(N__7203));
    Odrv4 I__1333 (
            .O(N__7212),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__1332 (
            .O(N__7209),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__1331 (
            .O(N__7206),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1330 (
            .O(N__7203),
            .I(DBR_SYNCZ0Z_1));
    CascadeMux I__1329 (
            .O(N__7194),
            .I(\U712_REG_SM.N_324_cascade_ ));
    InMux I__1328 (
            .O(N__7191),
            .I(N__7188));
    LocalMux I__1327 (
            .O(N__7188),
            .I(N__7184));
    InMux I__1326 (
            .O(N__7187),
            .I(N__7179));
    Span4Mux_v I__1325 (
            .O(N__7184),
            .I(N__7176));
    InMux I__1324 (
            .O(N__7183),
            .I(N__7171));
    InMux I__1323 (
            .O(N__7182),
            .I(N__7171));
    LocalMux I__1322 (
            .O(N__7179),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    Odrv4 I__1321 (
            .O(N__7176),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    LocalMux I__1320 (
            .O(N__7171),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    InMux I__1319 (
            .O(N__7164),
            .I(N__7161));
    LocalMux I__1318 (
            .O(N__7161),
            .I(\U712_REG_SM.STATE_COUNTc_0_0 ));
    InMux I__1317 (
            .O(N__7158),
            .I(N__7154));
    InMux I__1316 (
            .O(N__7157),
            .I(N__7151));
    LocalMux I__1315 (
            .O(N__7154),
            .I(\U712_BYTE_ENABLE.N_424 ));
    LocalMux I__1314 (
            .O(N__7151),
            .I(\U712_BYTE_ENABLE.N_424 ));
    InMux I__1313 (
            .O(N__7146),
            .I(N__7142));
    InMux I__1312 (
            .O(N__7145),
            .I(N__7139));
    LocalMux I__1311 (
            .O(N__7142),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0 ));
    LocalMux I__1310 (
            .O(N__7139),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0 ));
    IoInMux I__1309 (
            .O(N__7134),
            .I(N__7131));
    LocalMux I__1308 (
            .O(N__7131),
            .I(N__7128));
    IoSpan4Mux I__1307 (
            .O(N__7128),
            .I(N__7125));
    IoSpan4Mux I__1306 (
            .O(N__7125),
            .I(N__7122));
    Sp12to4 I__1305 (
            .O(N__7122),
            .I(N__7119));
    Span12Mux_s7_v I__1304 (
            .O(N__7119),
            .I(N__7116));
    Span12Mux_h I__1303 (
            .O(N__7116),
            .I(N__7113));
    Odrv12 I__1302 (
            .O(N__7113),
            .I(N_170_i));
    InMux I__1301 (
            .O(N__7110),
            .I(N__7107));
    LocalMux I__1300 (
            .O(N__7107),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__1299 (
            .O(N__7104),
            .I(N__7101));
    LocalMux I__1298 (
            .O(N__7101),
            .I(N__7098));
    Span12Mux_s6_v I__1297 (
            .O(N__7098),
            .I(N__7095));
    Odrv12 I__1296 (
            .O(N__7095),
            .I(CMA_c_2));
    InMux I__1295 (
            .O(N__7092),
            .I(N__7089));
    LocalMux I__1294 (
            .O(N__7089),
            .I(N__7086));
    Span4Mux_v I__1293 (
            .O(N__7086),
            .I(N__7083));
    Span4Mux_h I__1292 (
            .O(N__7083),
            .I(N__7080));
    Sp12to4 I__1291 (
            .O(N__7080),
            .I(N__7077));
    Odrv12 I__1290 (
            .O(N__7077),
            .I(A_c_7));
    InMux I__1289 (
            .O(N__7074),
            .I(N__7070));
    InMux I__1288 (
            .O(N__7073),
            .I(N__7067));
    LocalMux I__1287 (
            .O(N__7070),
            .I(N__7064));
    LocalMux I__1286 (
            .O(N__7067),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ));
    Odrv4 I__1285 (
            .O(N__7064),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ));
    InMux I__1284 (
            .O(N__7059),
            .I(N__7056));
    LocalMux I__1283 (
            .O(N__7056),
            .I(N__7053));
    Span12Mux_h I__1282 (
            .O(N__7053),
            .I(N__7050));
    Span12Mux_v I__1281 (
            .O(N__7050),
            .I(N__7047));
    Odrv12 I__1280 (
            .O(N__7047),
            .I(A_c_2));
    InMux I__1279 (
            .O(N__7044),
            .I(N__7040));
    InMux I__1278 (
            .O(N__7043),
            .I(N__7037));
    LocalMux I__1277 (
            .O(N__7040),
            .I(N__7034));
    LocalMux I__1276 (
            .O(N__7037),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ));
    Odrv4 I__1275 (
            .O(N__7034),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ));
    InMux I__1274 (
            .O(N__7029),
            .I(N__7026));
    LocalMux I__1273 (
            .O(N__7026),
            .I(N__7023));
    Span4Mux_v I__1272 (
            .O(N__7023),
            .I(N__7020));
    Sp12to4 I__1271 (
            .O(N__7020),
            .I(N__7017));
    Span12Mux_h I__1270 (
            .O(N__7017),
            .I(N__7014));
    Odrv12 I__1269 (
            .O(N__7014),
            .I(A_c_8));
    InMux I__1268 (
            .O(N__7011),
            .I(N__7008));
    LocalMux I__1267 (
            .O(N__7008),
            .I(N__6997));
    InMux I__1266 (
            .O(N__7007),
            .I(N__6994));
    InMux I__1265 (
            .O(N__7006),
            .I(N__6987));
    InMux I__1264 (
            .O(N__7005),
            .I(N__6987));
    InMux I__1263 (
            .O(N__7004),
            .I(N__6987));
    InMux I__1262 (
            .O(N__7003),
            .I(N__6984));
    InMux I__1261 (
            .O(N__7002),
            .I(N__6977));
    InMux I__1260 (
            .O(N__7001),
            .I(N__6977));
    InMux I__1259 (
            .O(N__7000),
            .I(N__6977));
    Span4Mux_h I__1258 (
            .O(N__6997),
            .I(N__6974));
    LocalMux I__1257 (
            .O(N__6994),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    LocalMux I__1256 (
            .O(N__6987),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    LocalMux I__1255 (
            .O(N__6984),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    LocalMux I__1254 (
            .O(N__6977),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    Odrv4 I__1253 (
            .O(N__6974),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    IoInMux I__1252 (
            .O(N__6963),
            .I(N__6960));
    LocalMux I__1251 (
            .O(N__6960),
            .I(N__6957));
    IoSpan4Mux I__1250 (
            .O(N__6957),
            .I(N__6954));
    Span4Mux_s2_h I__1249 (
            .O(N__6954),
            .I(N__6951));
    Sp12to4 I__1248 (
            .O(N__6951),
            .I(N__6948));
    Span12Mux_s11_h I__1247 (
            .O(N__6948),
            .I(N__6945));
    Span12Mux_v I__1246 (
            .O(N__6945),
            .I(N__6942));
    Odrv12 I__1245 (
            .O(N__6942),
            .I(CMA_c_4));
    IoInMux I__1244 (
            .O(N__6939),
            .I(N__6936));
    LocalMux I__1243 (
            .O(N__6936),
            .I(N__6933));
    IoSpan4Mux I__1242 (
            .O(N__6933),
            .I(N__6930));
    Span4Mux_s3_h I__1241 (
            .O(N__6930),
            .I(N__6927));
    Sp12to4 I__1240 (
            .O(N__6927),
            .I(N__6924));
    Span12Mux_h I__1239 (
            .O(N__6924),
            .I(N__6921));
    Span12Mux_v I__1238 (
            .O(N__6921),
            .I(N__6918));
    Odrv12 I__1237 (
            .O(N__6918),
            .I(CMA_c_3));
    IoInMux I__1236 (
            .O(N__6915),
            .I(N__6912));
    LocalMux I__1235 (
            .O(N__6912),
            .I(N__6909));
    Span12Mux_s7_h I__1234 (
            .O(N__6909),
            .I(N__6906));
    Span12Mux_v I__1233 (
            .O(N__6906),
            .I(N__6903));
    Odrv12 I__1232 (
            .O(N__6903),
            .I(CMA_c_6));
    CascadeMux I__1231 (
            .O(N__6900),
            .I(N__6895));
    CascadeMux I__1230 (
            .O(N__6899),
            .I(N__6889));
    CascadeMux I__1229 (
            .O(N__6898),
            .I(N__6886));
    InMux I__1228 (
            .O(N__6895),
            .I(N__6883));
    CascadeMux I__1227 (
            .O(N__6894),
            .I(N__6880));
    InMux I__1226 (
            .O(N__6893),
            .I(N__6870));
    InMux I__1225 (
            .O(N__6892),
            .I(N__6870));
    InMux I__1224 (
            .O(N__6889),
            .I(N__6870));
    InMux I__1223 (
            .O(N__6886),
            .I(N__6870));
    LocalMux I__1222 (
            .O(N__6883),
            .I(N__6867));
    InMux I__1221 (
            .O(N__6880),
            .I(N__6864));
    InMux I__1220 (
            .O(N__6879),
            .I(N__6861));
    LocalMux I__1219 (
            .O(N__6870),
            .I(N__6858));
    Span4Mux_h I__1218 (
            .O(N__6867),
            .I(N__6855));
    LocalMux I__1217 (
            .O(N__6864),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ));
    LocalMux I__1216 (
            .O(N__6861),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ));
    Odrv4 I__1215 (
            .O(N__6858),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ));
    Odrv4 I__1214 (
            .O(N__6855),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ));
    InMux I__1213 (
            .O(N__6846),
            .I(N__6843));
    LocalMux I__1212 (
            .O(N__6843),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__1211 (
            .O(N__6840),
            .I(N__6837));
    LocalMux I__1210 (
            .O(N__6837),
            .I(N__6834));
    IoSpan4Mux I__1209 (
            .O(N__6834),
            .I(N__6831));
    IoSpan4Mux I__1208 (
            .O(N__6831),
            .I(N__6828));
    Span4Mux_s3_h I__1207 (
            .O(N__6828),
            .I(N__6825));
    Sp12to4 I__1206 (
            .O(N__6825),
            .I(N__6822));
    Span12Mux_h I__1205 (
            .O(N__6822),
            .I(N__6819));
    Odrv12 I__1204 (
            .O(N__6819),
            .I(CMA_c_7));
    InMux I__1203 (
            .O(N__6816),
            .I(N__6812));
    InMux I__1202 (
            .O(N__6815),
            .I(N__6809));
    LocalMux I__1201 (
            .O(N__6812),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_5 ));
    LocalMux I__1200 (
            .O(N__6809),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_5 ));
    InMux I__1199 (
            .O(N__6804),
            .I(N__6800));
    InMux I__1198 (
            .O(N__6803),
            .I(N__6797));
    LocalMux I__1197 (
            .O(N__6800),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_4 ));
    LocalMux I__1196 (
            .O(N__6797),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_4 ));
    CascadeMux I__1195 (
            .O(N__6792),
            .I(N__6788));
    InMux I__1194 (
            .O(N__6791),
            .I(N__6785));
    InMux I__1193 (
            .O(N__6788),
            .I(N__6782));
    LocalMux I__1192 (
            .O(N__6785),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_3 ));
    LocalMux I__1191 (
            .O(N__6782),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_3 ));
    InMux I__1190 (
            .O(N__6777),
            .I(N__6773));
    InMux I__1189 (
            .O(N__6776),
            .I(N__6770));
    LocalMux I__1188 (
            .O(N__6773),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_7 ));
    LocalMux I__1187 (
            .O(N__6770),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_7 ));
    InMux I__1186 (
            .O(N__6765),
            .I(N__6762));
    LocalMux I__1185 (
            .O(N__6762),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLE_5_i_a2_5 ));
    IoInMux I__1184 (
            .O(N__6759),
            .I(N__6756));
    LocalMux I__1183 (
            .O(N__6756),
            .I(N__6753));
    IoSpan4Mux I__1182 (
            .O(N__6753),
            .I(N__6750));
    Span4Mux_s3_v I__1181 (
            .O(N__6750),
            .I(N__6747));
    Span4Mux_v I__1180 (
            .O(N__6747),
            .I(N__6744));
    Odrv4 I__1179 (
            .O(N__6744),
            .I(DMA_LATCH_EN_c));
    IoInMux I__1178 (
            .O(N__6741),
            .I(N__6738));
    LocalMux I__1177 (
            .O(N__6738),
            .I(N__6735));
    Span4Mux_s3_v I__1176 (
            .O(N__6735),
            .I(N__6732));
    Span4Mux_h I__1175 (
            .O(N__6732),
            .I(N__6729));
    Sp12to4 I__1174 (
            .O(N__6729),
            .I(N__6726));
    Span12Mux_v I__1173 (
            .O(N__6726),
            .I(N__6723));
    Odrv12 I__1172 (
            .O(N__6723),
            .I(CMA_c_10));
    IoInMux I__1171 (
            .O(N__6720),
            .I(N__6716));
    InMux I__1170 (
            .O(N__6719),
            .I(N__6713));
    LocalMux I__1169 (
            .O(N__6716),
            .I(N__6710));
    LocalMux I__1168 (
            .O(N__6713),
            .I(N__6707));
    Span12Mux_s4_v I__1167 (
            .O(N__6710),
            .I(N__6704));
    Span4Mux_v I__1166 (
            .O(N__6707),
            .I(N__6701));
    Span12Mux_h I__1165 (
            .O(N__6704),
            .I(N__6698));
    Span4Mux_h I__1164 (
            .O(N__6701),
            .I(N__6695));
    Span12Mux_v I__1163 (
            .O(N__6698),
            .I(N__6692));
    Sp12to4 I__1162 (
            .O(N__6695),
            .I(N__6689));
    Odrv12 I__1161 (
            .O(N__6692),
            .I(A_c_9));
    Odrv12 I__1160 (
            .O(N__6689),
            .I(A_c_9));
    CascadeMux I__1159 (
            .O(N__6684),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ));
    CascadeMux I__1158 (
            .O(N__6681),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_ ));
    IoInMux I__1157 (
            .O(N__6678),
            .I(N__6675));
    LocalMux I__1156 (
            .O(N__6675),
            .I(N__6672));
    Span4Mux_s3_v I__1155 (
            .O(N__6672),
            .I(N__6669));
    Sp12to4 I__1154 (
            .O(N__6669),
            .I(N__6666));
    Span12Mux_h I__1153 (
            .O(N__6666),
            .I(N__6663));
    Odrv12 I__1152 (
            .O(N__6663),
            .I(CMA_c_0));
    CascadeMux I__1151 (
            .O(N__6660),
            .I(\U712_REG_SM.N_408_cascade_ ));
    InMux I__1150 (
            .O(N__6657),
            .I(N__6654));
    LocalMux I__1149 (
            .O(N__6654),
            .I(\U712_REG_SM.N_367 ));
    InMux I__1148 (
            .O(N__6651),
            .I(N__6648));
    LocalMux I__1147 (
            .O(N__6648),
            .I(\U712_REG_SM.N_410 ));
    InMux I__1146 (
            .O(N__6645),
            .I(N__6641));
    InMux I__1145 (
            .O(N__6644),
            .I(N__6638));
    LocalMux I__1144 (
            .O(N__6641),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    LocalMux I__1143 (
            .O(N__6638),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    InMux I__1142 (
            .O(N__6633),
            .I(N__6630));
    LocalMux I__1141 (
            .O(N__6630),
            .I(\U712_REG_SM.REGENn_e_1 ));
    IoInMux I__1140 (
            .O(N__6627),
            .I(N__6624));
    LocalMux I__1139 (
            .O(N__6624),
            .I(N__6621));
    Span4Mux_s0_v I__1138 (
            .O(N__6621),
            .I(N__6618));
    Sp12to4 I__1137 (
            .O(N__6618),
            .I(N__6615));
    Span12Mux_s7_h I__1136 (
            .O(N__6615),
            .I(N__6612));
    Span12Mux_v I__1135 (
            .O(N__6612),
            .I(N__6607));
    InMux I__1134 (
            .O(N__6611),
            .I(N__6604));
    InMux I__1133 (
            .O(N__6610),
            .I(N__6601));
    Odrv12 I__1132 (
            .O(N__6607),
            .I(REGENn_c));
    LocalMux I__1131 (
            .O(N__6604),
            .I(REGENn_c));
    LocalMux I__1130 (
            .O(N__6601),
            .I(REGENn_c));
    InMux I__1129 (
            .O(N__6594),
            .I(N__6588));
    InMux I__1128 (
            .O(N__6593),
            .I(N__6588));
    LocalMux I__1127 (
            .O(N__6588),
            .I(\U712_REG_SM.N_322 ));
    InMux I__1126 (
            .O(N__6585),
            .I(N__6582));
    LocalMux I__1125 (
            .O(N__6582),
            .I(\U712_REG_SM.N_131 ));
    InMux I__1124 (
            .O(N__6579),
            .I(N__6576));
    LocalMux I__1123 (
            .O(N__6576),
            .I(N__6573));
    Span4Mux_v I__1122 (
            .O(N__6573),
            .I(N__6568));
    InMux I__1121 (
            .O(N__6572),
            .I(N__6563));
    InMux I__1120 (
            .O(N__6571),
            .I(N__6563));
    Odrv4 I__1119 (
            .O(N__6568),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    LocalMux I__1118 (
            .O(N__6563),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    CascadeMux I__1117 (
            .O(N__6558),
            .I(N__6554));
    InMux I__1116 (
            .O(N__6557),
            .I(N__6548));
    InMux I__1115 (
            .O(N__6554),
            .I(N__6548));
    InMux I__1114 (
            .O(N__6553),
            .I(N__6545));
    LocalMux I__1113 (
            .O(N__6548),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_1 ));
    LocalMux I__1112 (
            .O(N__6545),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_1 ));
    InMux I__1111 (
            .O(N__6540),
            .I(N__6536));
    InMux I__1110 (
            .O(N__6539),
            .I(N__6533));
    LocalMux I__1109 (
            .O(N__6536),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_6 ));
    LocalMux I__1108 (
            .O(N__6533),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_6 ));
    InMux I__1107 (
            .O(N__6528),
            .I(N__6524));
    InMux I__1106 (
            .O(N__6527),
            .I(N__6521));
    LocalMux I__1105 (
            .O(N__6524),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_2 ));
    LocalMux I__1104 (
            .O(N__6521),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_2 ));
    InMux I__1103 (
            .O(N__6516),
            .I(N__6510));
    InMux I__1102 (
            .O(N__6515),
            .I(N__6507));
    InMux I__1101 (
            .O(N__6514),
            .I(N__6502));
    InMux I__1100 (
            .O(N__6513),
            .I(N__6502));
    LocalMux I__1099 (
            .O(N__6510),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ));
    LocalMux I__1098 (
            .O(N__6507),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ));
    LocalMux I__1097 (
            .O(N__6502),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ));
    CascadeMux I__1096 (
            .O(N__6495),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLE_5_i_a2_4_cascade_ ));
    CascadeMux I__1095 (
            .O(N__6492),
            .I(N__6489));
    InMux I__1094 (
            .O(N__6489),
            .I(N__6486));
    LocalMux I__1093 (
            .O(N__6486),
            .I(N__6483));
    Span4Mux_h I__1092 (
            .O(N__6483),
            .I(N__6480));
    Odrv4 I__1091 (
            .O(N__6480),
            .I(\U712_CHIP_RAM.N_456 ));
    CascadeMux I__1090 (
            .O(N__6477),
            .I(\U712_CHIP_RAM.N_419_cascade_ ));
    InMux I__1089 (
            .O(N__6474),
            .I(N__6471));
    LocalMux I__1088 (
            .O(N__6471),
            .I(N__6468));
    Span4Mux_v I__1087 (
            .O(N__6468),
            .I(N__6465));
    Span4Mux_h I__1086 (
            .O(N__6465),
            .I(N__6462));
    Sp12to4 I__1085 (
            .O(N__6462),
            .I(N__6459));
    Odrv12 I__1084 (
            .O(N__6459),
            .I(RAMSPACEn_c));
    CascadeMux I__1083 (
            .O(N__6456),
            .I(N__6453));
    InMux I__1082 (
            .O(N__6453),
            .I(N__6450));
    LocalMux I__1081 (
            .O(N__6450),
            .I(N__6445));
    InMux I__1080 (
            .O(N__6449),
            .I(N__6442));
    InMux I__1079 (
            .O(N__6448),
            .I(N__6438));
    Span4Mux_v I__1078 (
            .O(N__6445),
            .I(N__6435));
    LocalMux I__1077 (
            .O(N__6442),
            .I(N__6432));
    InMux I__1076 (
            .O(N__6441),
            .I(N__6429));
    LocalMux I__1075 (
            .O(N__6438),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv4 I__1074 (
            .O(N__6435),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv4 I__1073 (
            .O(N__6432),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__1072 (
            .O(N__6429),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__1071 (
            .O(N__6420),
            .I(N__6415));
    InMux I__1070 (
            .O(N__6419),
            .I(N__6411));
    CascadeMux I__1069 (
            .O(N__6418),
            .I(N__6408));
    InMux I__1068 (
            .O(N__6415),
            .I(N__6405));
    CascadeMux I__1067 (
            .O(N__6414),
            .I(N__6401));
    LocalMux I__1066 (
            .O(N__6411),
            .I(N__6398));
    InMux I__1065 (
            .O(N__6408),
            .I(N__6394));
    LocalMux I__1064 (
            .O(N__6405),
            .I(N__6391));
    CascadeMux I__1063 (
            .O(N__6404),
            .I(N__6386));
    InMux I__1062 (
            .O(N__6401),
            .I(N__6380));
    Span4Mux_v I__1061 (
            .O(N__6398),
            .I(N__6372));
    InMux I__1060 (
            .O(N__6397),
            .I(N__6369));
    LocalMux I__1059 (
            .O(N__6394),
            .I(N__6364));
    Span4Mux_v I__1058 (
            .O(N__6391),
            .I(N__6364));
    InMux I__1057 (
            .O(N__6390),
            .I(N__6359));
    InMux I__1056 (
            .O(N__6389),
            .I(N__6359));
    InMux I__1055 (
            .O(N__6386),
            .I(N__6352));
    InMux I__1054 (
            .O(N__6385),
            .I(N__6352));
    InMux I__1053 (
            .O(N__6384),
            .I(N__6352));
    InMux I__1052 (
            .O(N__6383),
            .I(N__6349));
    LocalMux I__1051 (
            .O(N__6380),
            .I(N__6346));
    InMux I__1050 (
            .O(N__6379),
            .I(N__6343));
    InMux I__1049 (
            .O(N__6378),
            .I(N__6338));
    InMux I__1048 (
            .O(N__6377),
            .I(N__6338));
    InMux I__1047 (
            .O(N__6376),
            .I(N__6333));
    InMux I__1046 (
            .O(N__6375),
            .I(N__6333));
    Odrv4 I__1045 (
            .O(N__6372),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1044 (
            .O(N__6369),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1043 (
            .O(N__6364),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1042 (
            .O(N__6359),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1041 (
            .O(N__6352),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1040 (
            .O(N__6349),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1039 (
            .O(N__6346),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1038 (
            .O(N__6343),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1037 (
            .O(N__6338),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1036 (
            .O(N__6333),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1035 (
            .O(N__6312),
            .I(N__6308));
    InMux I__1034 (
            .O(N__6311),
            .I(N__6305));
    LocalMux I__1033 (
            .O(N__6308),
            .I(\U712_CHIP_RAM.N_299 ));
    LocalMux I__1032 (
            .O(N__6305),
            .I(\U712_CHIP_RAM.N_299 ));
    InMux I__1031 (
            .O(N__6300),
            .I(N__6297));
    LocalMux I__1030 (
            .O(N__6297),
            .I(N__6293));
    CascadeMux I__1029 (
            .O(N__6296),
            .I(N__6290));
    Span4Mux_h I__1028 (
            .O(N__6293),
            .I(N__6287));
    InMux I__1027 (
            .O(N__6290),
            .I(N__6284));
    Odrv4 I__1026 (
            .O(N__6287),
            .I(\U712_CHIP_RAM.N_307 ));
    LocalMux I__1025 (
            .O(N__6284),
            .I(\U712_CHIP_RAM.N_307 ));
    InMux I__1024 (
            .O(N__6279),
            .I(N__6276));
    LocalMux I__1023 (
            .O(N__6276),
            .I(\U712_CHIP_RAM.N_434 ));
    InMux I__1022 (
            .O(N__6273),
            .I(N__6270));
    LocalMux I__1021 (
            .O(N__6270),
            .I(N__6266));
    InMux I__1020 (
            .O(N__6269),
            .I(N__6263));
    Span4Mux_h I__1019 (
            .O(N__6266),
            .I(N__6260));
    LocalMux I__1018 (
            .O(N__6263),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv4 I__1017 (
            .O(N__6260),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__1016 (
            .O(N__6255),
            .I(N__6252));
    LocalMux I__1015 (
            .O(N__6252),
            .I(\U712_CHIP_RAM.REFRESH5lto7_0 ));
    InMux I__1014 (
            .O(N__6249),
            .I(N__6246));
    LocalMux I__1013 (
            .O(N__6246),
            .I(\U712_CHIP_RAM.REFRESH5lt7 ));
    InMux I__1012 (
            .O(N__6243),
            .I(N__6238));
    InMux I__1011 (
            .O(N__6242),
            .I(N__6233));
    InMux I__1010 (
            .O(N__6241),
            .I(N__6233));
    LocalMux I__1009 (
            .O(N__6238),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1008 (
            .O(N__6233),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    CascadeMux I__1007 (
            .O(N__6228),
            .I(\U712_REG_SM.N_322_cascade_ ));
    CascadeMux I__1006 (
            .O(N__6225),
            .I(\U712_REG_SM.N_367_cascade_ ));
    CascadeMux I__1005 (
            .O(N__6222),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ));
    InMux I__1004 (
            .O(N__6219),
            .I(N__6216));
    LocalMux I__1003 (
            .O(N__6216),
            .I(N__6212));
    InMux I__1002 (
            .O(N__6215),
            .I(N__6209));
    Span4Mux_v I__1001 (
            .O(N__6212),
            .I(N__6204));
    LocalMux I__1000 (
            .O(N__6209),
            .I(N__6204));
    Odrv4 I__999 (
            .O(N__6204),
            .I(\U712_CHIP_RAM.N_429 ));
    InMux I__998 (
            .O(N__6201),
            .I(N__6198));
    LocalMux I__997 (
            .O(N__6198),
            .I(N__6195));
    Odrv4 I__996 (
            .O(N__6195),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0 ));
    CascadeMux I__995 (
            .O(N__6192),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_cascade_ ));
    InMux I__994 (
            .O(N__6189),
            .I(N__6186));
    LocalMux I__993 (
            .O(N__6186),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__992 (
            .O(N__6183),
            .I(N__6179));
    InMux I__991 (
            .O(N__6182),
            .I(N__6176));
    LocalMux I__990 (
            .O(N__6179),
            .I(\U712_CHIP_RAM.N_319 ));
    LocalMux I__989 (
            .O(N__6176),
            .I(\U712_CHIP_RAM.N_319 ));
    InMux I__988 (
            .O(N__6171),
            .I(N__6168));
    LocalMux I__987 (
            .O(N__6168),
            .I(N__6165));
    Odrv12 I__986 (
            .O(N__6165),
            .I(\U712_CHIP_RAM.N_359 ));
    InMux I__985 (
            .O(N__6162),
            .I(N__6158));
    InMux I__984 (
            .O(N__6161),
            .I(N__6155));
    LocalMux I__983 (
            .O(N__6158),
            .I(N__6151));
    LocalMux I__982 (
            .O(N__6155),
            .I(N__6148));
    InMux I__981 (
            .O(N__6154),
            .I(N__6145));
    Span4Mux_v I__980 (
            .O(N__6151),
            .I(N__6142));
    Span4Mux_h I__979 (
            .O(N__6148),
            .I(N__6137));
    LocalMux I__978 (
            .O(N__6145),
            .I(N__6137));
    Sp12to4 I__977 (
            .O(N__6142),
            .I(N__6134));
    Span4Mux_v I__976 (
            .O(N__6137),
            .I(N__6131));
    Span12Mux_h I__975 (
            .O(N__6134),
            .I(N__6128));
    Span4Mux_h I__974 (
            .O(N__6131),
            .I(N__6125));
    Span12Mux_v I__973 (
            .O(N__6128),
            .I(N__6122));
    Sp12to4 I__972 (
            .O(N__6125),
            .I(N__6119));
    Odrv12 I__971 (
            .O(N__6122),
            .I(AWEn_c));
    Odrv12 I__970 (
            .O(N__6119),
            .I(AWEn_c));
    InMux I__969 (
            .O(N__6114),
            .I(N__6110));
    InMux I__968 (
            .O(N__6113),
            .I(N__6107));
    LocalMux I__967 (
            .O(N__6110),
            .I(N__6104));
    LocalMux I__966 (
            .O(N__6107),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    Odrv4 I__965 (
            .O(N__6104),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    InMux I__964 (
            .O(N__6099),
            .I(N__6096));
    LocalMux I__963 (
            .O(N__6096),
            .I(N__6093));
    Span4Mux_h I__962 (
            .O(N__6093),
            .I(N__6089));
    InMux I__961 (
            .O(N__6092),
            .I(N__6086));
    Odrv4 I__960 (
            .O(N__6089),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0_a2_0 ));
    LocalMux I__959 (
            .O(N__6086),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0_a2_0 ));
    InMux I__958 (
            .O(N__6081),
            .I(N__6077));
    InMux I__957 (
            .O(N__6080),
            .I(N__6074));
    LocalMux I__956 (
            .O(N__6077),
            .I(N__6071));
    LocalMux I__955 (
            .O(N__6074),
            .I(N__6068));
    Span4Mux_v I__954 (
            .O(N__6071),
            .I(N__6062));
    Span4Mux_v I__953 (
            .O(N__6068),
            .I(N__6062));
    InMux I__952 (
            .O(N__6067),
            .I(N__6059));
    Odrv4 I__951 (
            .O(N__6062),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__950 (
            .O(N__6059),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    IoInMux I__949 (
            .O(N__6054),
            .I(N__6051));
    LocalMux I__948 (
            .O(N__6051),
            .I(N__6048));
    IoSpan4Mux I__947 (
            .O(N__6048),
            .I(N__6045));
    Span4Mux_s0_v I__946 (
            .O(N__6045),
            .I(N__6042));
    Sp12to4 I__945 (
            .O(N__6042),
            .I(N__6039));
    Span12Mux_v I__944 (
            .O(N__6039),
            .I(N__6035));
    InMux I__943 (
            .O(N__6038),
            .I(N__6032));
    Odrv12 I__942 (
            .O(N__6035),
            .I(DBDIR_c));
    LocalMux I__941 (
            .O(N__6032),
            .I(DBDIR_c));
    InMux I__940 (
            .O(N__6027),
            .I(N__6024));
    LocalMux I__939 (
            .O(N__6024),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i ));
    InMux I__938 (
            .O(N__6021),
            .I(N__6018));
    LocalMux I__937 (
            .O(N__6018),
            .I(N__6015));
    Span12Mux_v I__936 (
            .O(N__6015),
            .I(N__6012));
    Span12Mux_h I__935 (
            .O(N__6012),
            .I(N__6009));
    Odrv12 I__934 (
            .O(N__6009),
            .I(A_c_12));
    InMux I__933 (
            .O(N__6006),
            .I(N__6003));
    LocalMux I__932 (
            .O(N__6003),
            .I(N__6000));
    Span4Mux_h I__931 (
            .O(N__6000),
            .I(N__5997));
    Span4Mux_v I__930 (
            .O(N__5997),
            .I(N__5994));
    Sp12to4 I__929 (
            .O(N__5994),
            .I(N__5991));
    Odrv12 I__928 (
            .O(N__5991),
            .I(A_c_5));
    InMux I__927 (
            .O(N__5988),
            .I(N__5982));
    InMux I__926 (
            .O(N__5987),
            .I(N__5982));
    LocalMux I__925 (
            .O(N__5982),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ));
    InMux I__924 (
            .O(N__5979),
            .I(N__5975));
    InMux I__923 (
            .O(N__5978),
            .I(N__5971));
    LocalMux I__922 (
            .O(N__5975),
            .I(N__5968));
    InMux I__921 (
            .O(N__5974),
            .I(N__5965));
    LocalMux I__920 (
            .O(N__5971),
            .I(\U712_CHIP_RAM.N_471 ));
    Odrv4 I__919 (
            .O(N__5968),
            .I(\U712_CHIP_RAM.N_471 ));
    LocalMux I__918 (
            .O(N__5965),
            .I(\U712_CHIP_RAM.N_471 ));
    InMux I__917 (
            .O(N__5958),
            .I(N__5955));
    LocalMux I__916 (
            .O(N__5955),
            .I(N__5952));
    Span12Mux_v I__915 (
            .O(N__5952),
            .I(N__5949));
    Span12Mux_h I__914 (
            .O(N__5949),
            .I(N__5946));
    Odrv12 I__913 (
            .O(N__5946),
            .I(A_c_3));
    CascadeMux I__912 (
            .O(N__5943),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ));
    InMux I__911 (
            .O(N__5940),
            .I(N__5937));
    LocalMux I__910 (
            .O(N__5937),
            .I(N__5934));
    Span12Mux_v I__909 (
            .O(N__5934),
            .I(N__5931));
    Span12Mux_h I__908 (
            .O(N__5931),
            .I(N__5928));
    Odrv12 I__907 (
            .O(N__5928),
            .I(A_c_4));
    InMux I__906 (
            .O(N__5925),
            .I(N__5921));
    InMux I__905 (
            .O(N__5924),
            .I(N__5918));
    LocalMux I__904 (
            .O(N__5921),
            .I(N__5915));
    LocalMux I__903 (
            .O(N__5918),
            .I(N__5912));
    Odrv4 I__902 (
            .O(N__5915),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ));
    Odrv4 I__901 (
            .O(N__5912),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ));
    InMux I__900 (
            .O(N__5907),
            .I(N__5904));
    LocalMux I__899 (
            .O(N__5904),
            .I(N__5901));
    Span4Mux_v I__898 (
            .O(N__5901),
            .I(N__5898));
    Sp12to4 I__897 (
            .O(N__5898),
            .I(N__5895));
    Span12Mux_h I__896 (
            .O(N__5895),
            .I(N__5892));
    Odrv12 I__895 (
            .O(N__5892),
            .I(A_c_6));
    SRMux I__894 (
            .O(N__5889),
            .I(N__5885));
    SRMux I__893 (
            .O(N__5888),
            .I(N__5882));
    LocalMux I__892 (
            .O(N__5885),
            .I(N__5879));
    LocalMux I__891 (
            .O(N__5882),
            .I(N__5876));
    Odrv4 I__890 (
            .O(N__5879),
            .I(\U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ));
    Odrv4 I__889 (
            .O(N__5876),
            .I(\U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ));
    IoInMux I__888 (
            .O(N__5871),
            .I(N__5867));
    InMux I__887 (
            .O(N__5870),
            .I(N__5864));
    LocalMux I__886 (
            .O(N__5867),
            .I(N__5861));
    LocalMux I__885 (
            .O(N__5864),
            .I(N__5858));
    IoSpan4Mux I__884 (
            .O(N__5861),
            .I(N__5855));
    Span4Mux_v I__883 (
            .O(N__5858),
            .I(N__5852));
    Span4Mux_s3_v I__882 (
            .O(N__5855),
            .I(N__5849));
    Span4Mux_v I__881 (
            .O(N__5852),
            .I(N__5846));
    Span4Mux_v I__880 (
            .O(N__5849),
            .I(N__5843));
    Odrv4 I__879 (
            .O(N__5846),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__878 (
            .O(N__5843),
            .I(CONSTANT_ONE_NET));
    IoInMux I__877 (
            .O(N__5838),
            .I(N__5835));
    LocalMux I__876 (
            .O(N__5835),
            .I(N__5832));
    IoSpan4Mux I__875 (
            .O(N__5832),
            .I(N__5829));
    Span4Mux_s0_v I__874 (
            .O(N__5829),
            .I(N__5826));
    Sp12to4 I__873 (
            .O(N__5826),
            .I(N__5823));
    Span12Mux_h I__872 (
            .O(N__5823),
            .I(N__5820));
    Span12Mux_v I__871 (
            .O(N__5820),
            .I(N__5817));
    Odrv12 I__870 (
            .O(N__5817),
            .I(CMA_c_5));
    IoInMux I__869 (
            .O(N__5814),
            .I(N__5811));
    LocalMux I__868 (
            .O(N__5811),
            .I(N__5808));
    IoSpan4Mux I__867 (
            .O(N__5808),
            .I(N__5805));
    Span4Mux_s2_v I__866 (
            .O(N__5805),
            .I(N__5801));
    InMux I__865 (
            .O(N__5804),
            .I(N__5798));
    Sp12to4 I__864 (
            .O(N__5801),
            .I(N__5795));
    LocalMux I__863 (
            .O(N__5798),
            .I(N__5792));
    Span12Mux_s8_v I__862 (
            .O(N__5795),
            .I(N__5789));
    Span4Mux_v I__861 (
            .O(N__5792),
            .I(N__5786));
    Span12Mux_v I__860 (
            .O(N__5789),
            .I(N__5783));
    Sp12to4 I__859 (
            .O(N__5786),
            .I(N__5780));
    Span12Mux_h I__858 (
            .O(N__5783),
            .I(N__5777));
    Span12Mux_h I__857 (
            .O(N__5780),
            .I(N__5774));
    Odrv12 I__856 (
            .O(N__5777),
            .I(A_c_11));
    Odrv12 I__855 (
            .O(N__5774),
            .I(A_c_11));
    CascadeMux I__854 (
            .O(N__5769),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ));
    InMux I__853 (
            .O(N__5766),
            .I(N__5763));
    LocalMux I__852 (
            .O(N__5763),
            .I(N__5760));
    Span4Mux_v I__851 (
            .O(N__5760),
            .I(N__5757));
    Span4Mux_v I__850 (
            .O(N__5757),
            .I(N__5754));
    Span4Mux_v I__849 (
            .O(N__5754),
            .I(N__5751));
    Sp12to4 I__848 (
            .O(N__5751),
            .I(N__5748));
    Span12Mux_h I__847 (
            .O(N__5748),
            .I(N__5745));
    Odrv12 I__846 (
            .O(N__5745),
            .I(A_c_17));
    CascadeMux I__845 (
            .O(N__5742),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ));
    InMux I__844 (
            .O(N__5739),
            .I(N__5735));
    InMux I__843 (
            .O(N__5738),
            .I(N__5732));
    LocalMux I__842 (
            .O(N__5735),
            .I(N__5729));
    LocalMux I__841 (
            .O(N__5732),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    Odrv4 I__840 (
            .O(N__5729),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    InMux I__839 (
            .O(N__5724),
            .I(N__5721));
    LocalMux I__838 (
            .O(N__5721),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ));
    InMux I__837 (
            .O(N__5718),
            .I(N__5715));
    LocalMux I__836 (
            .O(N__5715),
            .I(N__5712));
    Span12Mux_v I__835 (
            .O(N__5712),
            .I(N__5709));
    Span12Mux_h I__834 (
            .O(N__5709),
            .I(N__5706));
    Odrv12 I__833 (
            .O(N__5706),
            .I(A_c_14));
    InMux I__832 (
            .O(N__5703),
            .I(N__5700));
    LocalMux I__831 (
            .O(N__5700),
            .I(\U712_CHIP_RAM.N_353 ));
    InMux I__830 (
            .O(N__5697),
            .I(N__5694));
    LocalMux I__829 (
            .O(N__5694),
            .I(N__5691));
    Span12Mux_v I__828 (
            .O(N__5691),
            .I(N__5688));
    Span12Mux_h I__827 (
            .O(N__5688),
            .I(N__5685));
    Odrv12 I__826 (
            .O(N__5685),
            .I(A_c_20));
    CascadeMux I__825 (
            .O(N__5682),
            .I(N__5679));
    InMux I__824 (
            .O(N__5679),
            .I(N__5675));
    InMux I__823 (
            .O(N__5678),
            .I(N__5672));
    LocalMux I__822 (
            .O(N__5675),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    LocalMux I__821 (
            .O(N__5672),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    CascadeMux I__820 (
            .O(N__5667),
            .I(N__5664));
    InMux I__819 (
            .O(N__5664),
            .I(N__5661));
    LocalMux I__818 (
            .O(N__5661),
            .I(\U712_CHIP_RAM.DBENn_7_0_0 ));
    InMux I__817 (
            .O(N__5658),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_1 ));
    InMux I__816 (
            .O(N__5655),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_2 ));
    InMux I__815 (
            .O(N__5652),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_3 ));
    InMux I__814 (
            .O(N__5649),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_4 ));
    InMux I__813 (
            .O(N__5646),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_5 ));
    InMux I__812 (
            .O(N__5643),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_6 ));
    CascadeMux I__811 (
            .O(N__5640),
            .I(N__5631));
    InMux I__810 (
            .O(N__5639),
            .I(N__5624));
    InMux I__809 (
            .O(N__5638),
            .I(N__5624));
    InMux I__808 (
            .O(N__5637),
            .I(N__5624));
    InMux I__807 (
            .O(N__5636),
            .I(N__5621));
    InMux I__806 (
            .O(N__5635),
            .I(N__5618));
    InMux I__805 (
            .O(N__5634),
            .I(N__5613));
    InMux I__804 (
            .O(N__5631),
            .I(N__5613));
    LocalMux I__803 (
            .O(N__5624),
            .I(N__5606));
    LocalMux I__802 (
            .O(N__5621),
            .I(N__5606));
    LocalMux I__801 (
            .O(N__5618),
            .I(N__5606));
    LocalMux I__800 (
            .O(N__5613),
            .I(N__5600));
    Span4Mux_v I__799 (
            .O(N__5606),
            .I(N__5597));
    InMux I__798 (
            .O(N__5605),
            .I(N__5588));
    InMux I__797 (
            .O(N__5604),
            .I(N__5583));
    InMux I__796 (
            .O(N__5603),
            .I(N__5583));
    Span4Mux_h I__795 (
            .O(N__5600),
            .I(N__5578));
    Span4Mux_h I__794 (
            .O(N__5597),
            .I(N__5578));
    InMux I__793 (
            .O(N__5596),
            .I(N__5575));
    InMux I__792 (
            .O(N__5595),
            .I(N__5566));
    InMux I__791 (
            .O(N__5594),
            .I(N__5566));
    InMux I__790 (
            .O(N__5593),
            .I(N__5566));
    InMux I__789 (
            .O(N__5592),
            .I(N__5566));
    InMux I__788 (
            .O(N__5591),
            .I(N__5563));
    LocalMux I__787 (
            .O(N__5588),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__786 (
            .O(N__5583),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__785 (
            .O(N__5578),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__784 (
            .O(N__5575),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__783 (
            .O(N__5566),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__782 (
            .O(N__5563),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__781 (
            .O(N__5550),
            .I(N__5547));
    LocalMux I__780 (
            .O(N__5547),
            .I(N__5544));
    Odrv12 I__779 (
            .O(N__5544),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_0 ));
    CascadeMux I__778 (
            .O(N__5541),
            .I(N__5537));
    InMux I__777 (
            .O(N__5540),
            .I(N__5531));
    InMux I__776 (
            .O(N__5537),
            .I(N__5528));
    InMux I__775 (
            .O(N__5536),
            .I(N__5525));
    InMux I__774 (
            .O(N__5535),
            .I(N__5520));
    InMux I__773 (
            .O(N__5534),
            .I(N__5520));
    LocalMux I__772 (
            .O(N__5531),
            .I(N__5517));
    LocalMux I__771 (
            .O(N__5528),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__770 (
            .O(N__5525),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__769 (
            .O(N__5520),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__768 (
            .O(N__5517),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    InMux I__767 (
            .O(N__5508),
            .I(N__5505));
    LocalMux I__766 (
            .O(N__5505),
            .I(N__5502));
    Odrv12 I__765 (
            .O(N__5502),
            .I(\U712_CHIP_RAM.N_382 ));
    CascadeMux I__764 (
            .O(N__5499),
            .I(N__5494));
    InMux I__763 (
            .O(N__5498),
            .I(N__5490));
    InMux I__762 (
            .O(N__5497),
            .I(N__5487));
    InMux I__761 (
            .O(N__5494),
            .I(N__5482));
    InMux I__760 (
            .O(N__5493),
            .I(N__5482));
    LocalMux I__759 (
            .O(N__5490),
            .I(N__5474));
    LocalMux I__758 (
            .O(N__5487),
            .I(N__5474));
    LocalMux I__757 (
            .O(N__5482),
            .I(N__5474));
    InMux I__756 (
            .O(N__5481),
            .I(N__5471));
    Odrv4 I__755 (
            .O(N__5474),
            .I(\U712_CHIP_RAM.N_534 ));
    LocalMux I__754 (
            .O(N__5471),
            .I(\U712_CHIP_RAM.N_534 ));
    CascadeMux I__753 (
            .O(N__5466),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_cascade_ ));
    CascadeMux I__752 (
            .O(N__5463),
            .I(\U712_REG_SM.N_411_cascade_ ));
    CascadeMux I__751 (
            .O(N__5460),
            .I(\U712_BYTE_ENABLE.N_446_cascade_ ));
    IoInMux I__750 (
            .O(N__5457),
            .I(N__5454));
    LocalMux I__749 (
            .O(N__5454),
            .I(N__5451));
    IoSpan4Mux I__748 (
            .O(N__5451),
            .I(N__5448));
    Span4Mux_s3_v I__747 (
            .O(N__5448),
            .I(N__5445));
    Sp12to4 I__746 (
            .O(N__5445),
            .I(N__5442));
    Span12Mux_s11_v I__745 (
            .O(N__5442),
            .I(N__5439));
    Odrv12 I__744 (
            .O(N__5439),
            .I(N_52_i));
    InMux I__743 (
            .O(N__5436),
            .I(N__5433));
    LocalMux I__742 (
            .O(N__5433),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    CascadeMux I__741 (
            .O(N__5430),
            .I(\U712_CHIP_RAM.N_399_cascade_ ));
    InMux I__740 (
            .O(N__5427),
            .I(N__5424));
    LocalMux I__739 (
            .O(N__5424),
            .I(N__5420));
    InMux I__738 (
            .O(N__5423),
            .I(N__5417));
    Span4Mux_h I__737 (
            .O(N__5420),
            .I(N__5414));
    LocalMux I__736 (
            .O(N__5417),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    Odrv4 I__735 (
            .O(N__5414),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__734 (
            .O(N__5409),
            .I(N__5406));
    LocalMux I__733 (
            .O(N__5406),
            .I(N__5402));
    InMux I__732 (
            .O(N__5405),
            .I(N__5399));
    Span4Mux_h I__731 (
            .O(N__5402),
            .I(N__5396));
    LocalMux I__730 (
            .O(N__5399),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    Odrv4 I__729 (
            .O(N__5396),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    CascadeMux I__728 (
            .O(N__5391),
            .I(N__5388));
    InMux I__727 (
            .O(N__5388),
            .I(N__5385));
    LocalMux I__726 (
            .O(N__5385),
            .I(N__5381));
    InMux I__725 (
            .O(N__5384),
            .I(N__5378));
    Span4Mux_h I__724 (
            .O(N__5381),
            .I(N__5375));
    LocalMux I__723 (
            .O(N__5378),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    Odrv4 I__722 (
            .O(N__5375),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__721 (
            .O(N__5370),
            .I(N__5367));
    LocalMux I__720 (
            .O(N__5367),
            .I(N__5363));
    InMux I__719 (
            .O(N__5366),
            .I(N__5360));
    Span4Mux_v I__718 (
            .O(N__5363),
            .I(N__5357));
    LocalMux I__717 (
            .O(N__5360),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    Odrv4 I__716 (
            .O(N__5357),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__715 (
            .O(N__5352),
            .I(N__5349));
    LocalMux I__714 (
            .O(N__5349),
            .I(N__5346));
    Span4Mux_v I__713 (
            .O(N__5346),
            .I(N__5343));
    Odrv4 I__712 (
            .O(N__5343),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_0_3 ));
    CascadeMux I__711 (
            .O(N__5340),
            .I(N__5337));
    InMux I__710 (
            .O(N__5337),
            .I(N__5334));
    LocalMux I__709 (
            .O(N__5334),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__708 (
            .O(N__5331),
            .I(N__5328));
    LocalMux I__707 (
            .O(N__5328),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1 ));
    InMux I__706 (
            .O(N__5325),
            .I(N__5322));
    LocalMux I__705 (
            .O(N__5322),
            .I(N__5318));
    InMux I__704 (
            .O(N__5321),
            .I(N__5315));
    Span4Mux_v I__703 (
            .O(N__5318),
            .I(N__5312));
    LocalMux I__702 (
            .O(N__5315),
            .I(N__5309));
    Odrv4 I__701 (
            .O(N__5312),
            .I(\U712_CHIP_RAM.N_310 ));
    Odrv4 I__700 (
            .O(N__5309),
            .I(\U712_CHIP_RAM.N_310 ));
    InMux I__699 (
            .O(N__5304),
            .I(N__5301));
    LocalMux I__698 (
            .O(N__5301),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0 ));
    CEMux I__697 (
            .O(N__5298),
            .I(N__5294));
    CEMux I__696 (
            .O(N__5297),
            .I(N__5291));
    LocalMux I__695 (
            .O(N__5294),
            .I(N__5286));
    LocalMux I__694 (
            .O(N__5291),
            .I(N__5286));
    Span4Mux_v I__693 (
            .O(N__5286),
            .I(N__5283));
    Odrv4 I__692 (
            .O(N__5283),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    CascadeMux I__691 (
            .O(N__5280),
            .I(N__5273));
    CascadeMux I__690 (
            .O(N__5279),
            .I(N__5268));
    CascadeMux I__689 (
            .O(N__5278),
            .I(N__5265));
    CascadeMux I__688 (
            .O(N__5277),
            .I(N__5261));
    CascadeMux I__687 (
            .O(N__5276),
            .I(N__5258));
    InMux I__686 (
            .O(N__5273),
            .I(N__5254));
    InMux I__685 (
            .O(N__5272),
            .I(N__5251));
    InMux I__684 (
            .O(N__5271),
            .I(N__5247));
    InMux I__683 (
            .O(N__5268),
            .I(N__5242));
    InMux I__682 (
            .O(N__5265),
            .I(N__5242));
    InMux I__681 (
            .O(N__5264),
            .I(N__5239));
    InMux I__680 (
            .O(N__5261),
            .I(N__5234));
    InMux I__679 (
            .O(N__5258),
            .I(N__5234));
    CascadeMux I__678 (
            .O(N__5257),
            .I(N__5226));
    LocalMux I__677 (
            .O(N__5254),
            .I(N__5219));
    LocalMux I__676 (
            .O(N__5251),
            .I(N__5219));
    InMux I__675 (
            .O(N__5250),
            .I(N__5216));
    LocalMux I__674 (
            .O(N__5247),
            .I(N__5209));
    LocalMux I__673 (
            .O(N__5242),
            .I(N__5209));
    LocalMux I__672 (
            .O(N__5239),
            .I(N__5209));
    LocalMux I__671 (
            .O(N__5234),
            .I(N__5206));
    InMux I__670 (
            .O(N__5233),
            .I(N__5201));
    InMux I__669 (
            .O(N__5232),
            .I(N__5201));
    InMux I__668 (
            .O(N__5231),
            .I(N__5198));
    InMux I__667 (
            .O(N__5230),
            .I(N__5195));
    InMux I__666 (
            .O(N__5229),
            .I(N__5186));
    InMux I__665 (
            .O(N__5226),
            .I(N__5186));
    InMux I__664 (
            .O(N__5225),
            .I(N__5186));
    InMux I__663 (
            .O(N__5224),
            .I(N__5186));
    Odrv4 I__662 (
            .O(N__5219),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__661 (
            .O(N__5216),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__660 (
            .O(N__5209),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv12 I__659 (
            .O(N__5206),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__658 (
            .O(N__5201),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__657 (
            .O(N__5198),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__656 (
            .O(N__5195),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__655 (
            .O(N__5186),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__654 (
            .O(N__5169),
            .I(N__5166));
    LocalMux I__653 (
            .O(N__5166),
            .I(N__5163));
    Odrv4 I__652 (
            .O(N__5163),
            .I(\U712_CHIP_RAM.N_385 ));
    InMux I__651 (
            .O(N__5160),
            .I(N__5146));
    InMux I__650 (
            .O(N__5159),
            .I(N__5146));
    InMux I__649 (
            .O(N__5158),
            .I(N__5146));
    InMux I__648 (
            .O(N__5157),
            .I(N__5141));
    InMux I__647 (
            .O(N__5156),
            .I(N__5141));
    InMux I__646 (
            .O(N__5155),
            .I(N__5134));
    InMux I__645 (
            .O(N__5154),
            .I(N__5134));
    InMux I__644 (
            .O(N__5153),
            .I(N__5134));
    LocalMux I__643 (
            .O(N__5146),
            .I(\U712_CHIP_RAM.N_182 ));
    LocalMux I__642 (
            .O(N__5141),
            .I(\U712_CHIP_RAM.N_182 ));
    LocalMux I__641 (
            .O(N__5134),
            .I(\U712_CHIP_RAM.N_182 ));
    InMux I__640 (
            .O(N__5127),
            .I(N__5123));
    InMux I__639 (
            .O(N__5126),
            .I(N__5120));
    LocalMux I__638 (
            .O(N__5123),
            .I(N__5115));
    LocalMux I__637 (
            .O(N__5120),
            .I(N__5115));
    Odrv4 I__636 (
            .O(N__5115),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__635 (
            .O(N__5112),
            .I(N__5108));
    InMux I__634 (
            .O(N__5111),
            .I(N__5105));
    LocalMux I__633 (
            .O(N__5108),
            .I(N__5102));
    LocalMux I__632 (
            .O(N__5105),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    Odrv4 I__631 (
            .O(N__5102),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__630 (
            .O(N__5097),
            .I(N__5094));
    LocalMux I__629 (
            .O(N__5094),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_0_4 ));
    InMux I__628 (
            .O(N__5091),
            .I(N__5084));
    InMux I__627 (
            .O(N__5090),
            .I(N__5084));
    InMux I__626 (
            .O(N__5089),
            .I(N__5081));
    LocalMux I__625 (
            .O(N__5084),
            .I(\U712_CHIP_RAM.N_191 ));
    LocalMux I__624 (
            .O(N__5081),
            .I(\U712_CHIP_RAM.N_191 ));
    InMux I__623 (
            .O(N__5076),
            .I(N__5072));
    InMux I__622 (
            .O(N__5075),
            .I(N__5069));
    LocalMux I__621 (
            .O(N__5072),
            .I(\U712_CHIP_RAM.N_327 ));
    LocalMux I__620 (
            .O(N__5069),
            .I(\U712_CHIP_RAM.N_327 ));
    InMux I__619 (
            .O(N__5064),
            .I(N__5059));
    InMux I__618 (
            .O(N__5063),
            .I(N__5054));
    InMux I__617 (
            .O(N__5062),
            .I(N__5054));
    LocalMux I__616 (
            .O(N__5059),
            .I(\U712_CHIP_RAM.N_300 ));
    LocalMux I__615 (
            .O(N__5054),
            .I(\U712_CHIP_RAM.N_300 ));
    InMux I__614 (
            .O(N__5049),
            .I(N__5046));
    LocalMux I__613 (
            .O(N__5046),
            .I(\U712_CHIP_RAM.N_370 ));
    CascadeMux I__612 (
            .O(N__5043),
            .I(N__5034));
    InMux I__611 (
            .O(N__5042),
            .I(N__5031));
    InMux I__610 (
            .O(N__5041),
            .I(N__5028));
    InMux I__609 (
            .O(N__5040),
            .I(N__5025));
    InMux I__608 (
            .O(N__5039),
            .I(N__5022));
    InMux I__607 (
            .O(N__5038),
            .I(N__5017));
    InMux I__606 (
            .O(N__5037),
            .I(N__5017));
    InMux I__605 (
            .O(N__5034),
            .I(N__5014));
    LocalMux I__604 (
            .O(N__5031),
            .I(\U712_CHIP_RAM.N_301 ));
    LocalMux I__603 (
            .O(N__5028),
            .I(\U712_CHIP_RAM.N_301 ));
    LocalMux I__602 (
            .O(N__5025),
            .I(\U712_CHIP_RAM.N_301 ));
    LocalMux I__601 (
            .O(N__5022),
            .I(\U712_CHIP_RAM.N_301 ));
    LocalMux I__600 (
            .O(N__5017),
            .I(\U712_CHIP_RAM.N_301 ));
    LocalMux I__599 (
            .O(N__5014),
            .I(\U712_CHIP_RAM.N_301 ));
    CascadeMux I__598 (
            .O(N__5001),
            .I(\U712_CHIP_RAM.N_466_cascade_ ));
    CascadeMux I__597 (
            .O(N__4998),
            .I(\U712_CHIP_RAM.N_299_cascade_ ));
    InMux I__596 (
            .O(N__4995),
            .I(N__4991));
    InMux I__595 (
            .O(N__4994),
            .I(N__4988));
    LocalMux I__594 (
            .O(N__4991),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ));
    LocalMux I__593 (
            .O(N__4988),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ));
    InMux I__592 (
            .O(N__4983),
            .I(N__4980));
    LocalMux I__591 (
            .O(N__4980),
            .I(N__4977));
    Span12Mux_h I__590 (
            .O(N__4977),
            .I(N__4974));
    Span12Mux_v I__589 (
            .O(N__4974),
            .I(N__4971));
    Odrv12 I__588 (
            .O(N__4971),
            .I(A_c_16));
    InMux I__587 (
            .O(N__4968),
            .I(N__4965));
    LocalMux I__586 (
            .O(N__4965),
            .I(\U712_CHIP_RAM.CMA_5_i_0_9 ));
    InMux I__585 (
            .O(N__4962),
            .I(N__4959));
    LocalMux I__584 (
            .O(N__4959),
            .I(N__4956));
    Span4Mux_h I__583 (
            .O(N__4956),
            .I(N__4953));
    Sp12to4 I__582 (
            .O(N__4953),
            .I(N__4950));
    Span12Mux_v I__581 (
            .O(N__4950),
            .I(N__4947));
    Odrv12 I__580 (
            .O(N__4947),
            .I(A_c_19));
    IoInMux I__579 (
            .O(N__4944),
            .I(N__4941));
    LocalMux I__578 (
            .O(N__4941),
            .I(N__4938));
    Span12Mux_s7_h I__577 (
            .O(N__4938),
            .I(N__4935));
    Span12Mux_h I__576 (
            .O(N__4935),
            .I(N__4932));
    Odrv12 I__575 (
            .O(N__4932),
            .I(CMA_c_9));
    SRMux I__574 (
            .O(N__4929),
            .I(N__4926));
    LocalMux I__573 (
            .O(N__4926),
            .I(N__4922));
    InMux I__572 (
            .O(N__4925),
            .I(N__4919));
    Span4Mux_v I__571 (
            .O(N__4922),
            .I(N__4916));
    LocalMux I__570 (
            .O(N__4919),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    Odrv4 I__569 (
            .O(N__4916),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__568 (
            .O(N__4911),
            .I(N__4906));
    InMux I__567 (
            .O(N__4910),
            .I(N__4903));
    InMux I__566 (
            .O(N__4909),
            .I(N__4899));
    LocalMux I__565 (
            .O(N__4906),
            .I(N__4896));
    LocalMux I__564 (
            .O(N__4903),
            .I(N__4893));
    InMux I__563 (
            .O(N__4902),
            .I(N__4890));
    LocalMux I__562 (
            .O(N__4899),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    Odrv4 I__561 (
            .O(N__4896),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    Odrv4 I__560 (
            .O(N__4893),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__559 (
            .O(N__4890),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__558 (
            .O(N__4881),
            .I(N__4878));
    InMux I__557 (
            .O(N__4878),
            .I(N__4875));
    LocalMux I__556 (
            .O(N__4875),
            .I(N__4870));
    InMux I__555 (
            .O(N__4874),
            .I(N__4867));
    InMux I__554 (
            .O(N__4873),
            .I(N__4863));
    Span4Mux_h I__553 (
            .O(N__4870),
            .I(N__4860));
    LocalMux I__552 (
            .O(N__4867),
            .I(N__4857));
    InMux I__551 (
            .O(N__4866),
            .I(N__4854));
    LocalMux I__550 (
            .O(N__4863),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    Odrv4 I__549 (
            .O(N__4860),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    Odrv12 I__548 (
            .O(N__4857),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__547 (
            .O(N__4854),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__546 (
            .O(N__4845),
            .I(N__4842));
    LocalMux I__545 (
            .O(N__4842),
            .I(N__4839));
    Odrv4 I__544 (
            .O(N__4839),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_2 ));
    CascadeMux I__543 (
            .O(N__4836),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_ ));
    CascadeMux I__542 (
            .O(N__4833),
            .I(N__4830));
    InMux I__541 (
            .O(N__4830),
            .I(N__4827));
    LocalMux I__540 (
            .O(N__4827),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_1 ));
    CascadeMux I__539 (
            .O(N__4824),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_3_cascade_ ));
    CascadeMux I__538 (
            .O(N__4821),
            .I(\U712_CHIP_RAM.N_191_cascade_ ));
    CEMux I__537 (
            .O(N__4818),
            .I(N__4815));
    LocalMux I__536 (
            .O(N__4815),
            .I(\U712_CHIP_RAM.N_191_0 ));
    InMux I__535 (
            .O(N__4812),
            .I(N__4809));
    LocalMux I__534 (
            .O(N__4809),
            .I(N__4806));
    Span12Mux_h I__533 (
            .O(N__4806),
            .I(N__4803));
    Span12Mux_v I__532 (
            .O(N__4803),
            .I(N__4800));
    Odrv12 I__531 (
            .O(N__4800),
            .I(A_c_18));
    InMux I__530 (
            .O(N__4797),
            .I(N__4794));
    LocalMux I__529 (
            .O(N__4794),
            .I(N__4790));
    InMux I__528 (
            .O(N__4793),
            .I(N__4787));
    Odrv4 I__527 (
            .O(N__4790),
            .I(\U712_CHIP_RAM.N_315 ));
    LocalMux I__526 (
            .O(N__4787),
            .I(\U712_CHIP_RAM.N_315 ));
    CascadeMux I__525 (
            .O(N__4782),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_ ));
    InMux I__524 (
            .O(N__4779),
            .I(N__4776));
    LocalMux I__523 (
            .O(N__4776),
            .I(\U712_CHIP_RAM.N_336 ));
    InMux I__522 (
            .O(N__4773),
            .I(N__4770));
    LocalMux I__521 (
            .O(N__4770),
            .I(N__4767));
    Odrv4 I__520 (
            .O(N__4767),
            .I(\U712_CHIP_RAM.N_372 ));
    IoInMux I__519 (
            .O(N__4764),
            .I(N__4761));
    LocalMux I__518 (
            .O(N__4761),
            .I(N__4758));
    IoSpan4Mux I__517 (
            .O(N__4758),
            .I(N__4755));
    Span4Mux_s0_h I__516 (
            .O(N__4755),
            .I(N__4752));
    Sp12to4 I__515 (
            .O(N__4752),
            .I(N__4749));
    Span12Mux_h I__514 (
            .O(N__4749),
            .I(N__4746));
    Span12Mux_v I__513 (
            .O(N__4746),
            .I(N__4743));
    Odrv12 I__512 (
            .O(N__4743),
            .I(CMA_c_8));
    InMux I__511 (
            .O(N__4740),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__510 (
            .O(N__4737),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__509 (
            .O(N__4734),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    CascadeMux I__508 (
            .O(N__4731),
            .I(N__4728));
    InMux I__507 (
            .O(N__4728),
            .I(N__4724));
    InMux I__506 (
            .O(N__4727),
            .I(N__4719));
    LocalMux I__505 (
            .O(N__4724),
            .I(N__4716));
    InMux I__504 (
            .O(N__4723),
            .I(N__4711));
    InMux I__503 (
            .O(N__4722),
            .I(N__4711));
    LocalMux I__502 (
            .O(N__4719),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    Odrv4 I__501 (
            .O(N__4716),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__500 (
            .O(N__4711),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__499 (
            .O(N__4704),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__498 (
            .O(N__4701),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__497 (
            .O(N__4698),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__496 (
            .O(N__4695),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    InMux I__495 (
            .O(N__4692),
            .I(N__4687));
    CascadeMux I__494 (
            .O(N__4691),
            .I(N__4683));
    InMux I__493 (
            .O(N__4690),
            .I(N__4680));
    LocalMux I__492 (
            .O(N__4687),
            .I(N__4677));
    InMux I__491 (
            .O(N__4686),
            .I(N__4672));
    InMux I__490 (
            .O(N__4683),
            .I(N__4672));
    LocalMux I__489 (
            .O(N__4680),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    Odrv12 I__488 (
            .O(N__4677),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__487 (
            .O(N__4672),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__486 (
            .O(N__4665),
            .I(N__4662));
    LocalMux I__485 (
            .O(N__4662),
            .I(\U712_CHIP_RAM.LATCH_CLK_6 ));
    CascadeMux I__484 (
            .O(N__4659),
            .I(\U712_CHIP_RAM.N_396_cascade_ ));
    IoInMux I__483 (
            .O(N__4656),
            .I(N__4653));
    LocalMux I__482 (
            .O(N__4653),
            .I(N__4650));
    Span12Mux_s1_v I__481 (
            .O(N__4650),
            .I(N__4647));
    Span12Mux_v I__480 (
            .O(N__4647),
            .I(N__4643));
    InMux I__479 (
            .O(N__4646),
            .I(N__4640));
    Odrv12 I__478 (
            .O(N__4643),
            .I(LATCH_CLK_c));
    LocalMux I__477 (
            .O(N__4640),
            .I(LATCH_CLK_c));
    CascadeMux I__476 (
            .O(N__4635),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_2_0_cascade_ ));
    InMux I__475 (
            .O(N__4632),
            .I(N__4629));
    LocalMux I__474 (
            .O(N__4629),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_2_3 ));
    CascadeMux I__473 (
            .O(N__4626),
            .I(\U712_CHIP_RAM.N_301_cascade_ ));
    CascadeMux I__472 (
            .O(N__4623),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_0_1_cascade_ ));
    CascadeMux I__471 (
            .O(N__4620),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_1_5_cascade_ ));
    InMux I__470 (
            .O(N__4617),
            .I(N__4614));
    LocalMux I__469 (
            .O(N__4614),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_1_4 ));
    CascadeMux I__468 (
            .O(N__4611),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_2_2_cascade_ ));
    InMux I__467 (
            .O(N__4608),
            .I(N__4602));
    InMux I__466 (
            .O(N__4607),
            .I(N__4602));
    LocalMux I__465 (
            .O(N__4602),
            .I(\U712_CHIP_RAM.N_433 ));
    CascadeMux I__464 (
            .O(N__4599),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_4_i_2_cascade_ ));
    InMux I__463 (
            .O(N__4596),
            .I(N__4593));
    LocalMux I__462 (
            .O(N__4593),
            .I(N__4590));
    Odrv4 I__461 (
            .O(N__4590),
            .I(\U712_CHIP_RAM.N_65 ));
    CascadeMux I__460 (
            .O(N__4587),
            .I(\U712_CHIP_RAM.N_173_cascade_ ));
    IoInMux I__459 (
            .O(N__4584),
            .I(N__4581));
    LocalMux I__458 (
            .O(N__4581),
            .I(N__4578));
    Span12Mux_s8_v I__457 (
            .O(N__4578),
            .I(N__4575));
    Odrv12 I__456 (
            .O(N__4575),
            .I(VBENn_c));
    InMux I__455 (
            .O(N__4572),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__454 (
            .O(N__4569),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__453 (
            .O(N__4566),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__452 (
            .O(N__4563),
            .I(N__4539));
    ClkMux I__451 (
            .O(N__4562),
            .I(N__4539));
    ClkMux I__450 (
            .O(N__4561),
            .I(N__4539));
    ClkMux I__449 (
            .O(N__4560),
            .I(N__4539));
    ClkMux I__448 (
            .O(N__4559),
            .I(N__4539));
    ClkMux I__447 (
            .O(N__4558),
            .I(N__4539));
    ClkMux I__446 (
            .O(N__4557),
            .I(N__4539));
    ClkMux I__445 (
            .O(N__4556),
            .I(N__4539));
    GlobalMux I__444 (
            .O(N__4539),
            .I(N__4536));
    gio2CtrlBuf I__443 (
            .O(N__4536),
            .I(C1_c_g));
    InMux I__442 (
            .O(N__4533),
            .I(N__4529));
    InMux I__441 (
            .O(N__4532),
            .I(N__4526));
    LocalMux I__440 (
            .O(N__4529),
            .I(N__4523));
    LocalMux I__439 (
            .O(N__4526),
            .I(N__4520));
    Span4Mux_v I__438 (
            .O(N__4523),
            .I(N__4517));
    Span4Mux_v I__437 (
            .O(N__4520),
            .I(N__4514));
    Span4Mux_h I__436 (
            .O(N__4517),
            .I(N__4511));
    Sp12to4 I__435 (
            .O(N__4514),
            .I(N__4508));
    Sp12to4 I__434 (
            .O(N__4511),
            .I(N__4503));
    Span12Mux_h I__433 (
            .O(N__4508),
            .I(N__4503));
    Odrv12 I__432 (
            .O(N__4503),
            .I(DBRn_c));
    InMux I__431 (
            .O(N__4500),
            .I(N__4497));
    LocalMux I__430 (
            .O(N__4497),
            .I(DBR_SYNCZ0Z_0));
    InMux I__429 (
            .O(N__4494),
            .I(N__4491));
    LocalMux I__428 (
            .O(N__4491),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_1_1 ));
    CascadeMux I__427 (
            .O(N__4488),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_1_0_cascade_ ));
    CascadeMux I__426 (
            .O(N__4485),
            .I(\U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1_cascade_ ));
    CascadeMux I__425 (
            .O(N__4482),
            .I(\U712_CHIP_RAM.N_442_cascade_ ));
    InMux I__424 (
            .O(N__4479),
            .I(N__4473));
    InMux I__423 (
            .O(N__4478),
            .I(N__4473));
    LocalMux I__422 (
            .O(N__4473),
            .I(\U712_CHIP_RAM.CLK_EN_5_0 ));
    InMux I__421 (
            .O(N__4470),
            .I(N__4467));
    LocalMux I__420 (
            .O(N__4467),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__419 (
            .O(N__4464),
            .I(bfn_7_13_0_));
    InMux I__418 (
            .O(N__4461),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__417 (
            .O(N__4458),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__416 (
            .O(N__4455),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__415 (
            .O(N__4452),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    CascadeMux I__414 (
            .O(N__4449),
            .I(N__4446));
    InMux I__413 (
            .O(N__4446),
            .I(N__4443));
    LocalMux I__412 (
            .O(N__4443),
            .I(N__4439));
    InMux I__411 (
            .O(N__4442),
            .I(N__4436));
    Span4Mux_h I__410 (
            .O(N__4439),
            .I(N__4433));
    LocalMux I__409 (
            .O(N__4436),
            .I(N__4430));
    Span4Mux_v I__408 (
            .O(N__4433),
            .I(N__4427));
    Span4Mux_h I__407 (
            .O(N__4430),
            .I(N__4424));
    Odrv4 I__406 (
            .O(N__4427),
            .I(DBRn_c_i));
    Odrv4 I__405 (
            .O(N__4424),
            .I(DBRn_c_i));
    InMux I__404 (
            .O(N__4419),
            .I(N__4416));
    LocalMux I__403 (
            .O(N__4416),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_5 ));
    CascadeMux I__402 (
            .O(N__4413),
            .I(\U712_CHIP_RAM.N_458_cascade_ ));
    CascadeMux I__401 (
            .O(N__4410),
            .I(N__4407));
    InMux I__400 (
            .O(N__4407),
            .I(N__4401));
    InMux I__399 (
            .O(N__4406),
            .I(N__4401));
    LocalMux I__398 (
            .O(N__4401),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ));
    CascadeMux I__397 (
            .O(N__4398),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a2_0_cascade_ ));
    IoInMux I__396 (
            .O(N__4395),
            .I(N__4392));
    LocalMux I__395 (
            .O(N__4392),
            .I(N__4389));
    Span12Mux_s2_h I__394 (
            .O(N__4389),
            .I(N__4386));
    Span12Mux_h I__393 (
            .O(N__4386),
            .I(N__4383));
    Span12Mux_v I__392 (
            .O(N__4383),
            .I(N__4379));
    InMux I__391 (
            .O(N__4382),
            .I(N__4376));
    Odrv12 I__390 (
            .O(N__4379),
            .I(CLK_EN_c));
    LocalMux I__389 (
            .O(N__4376),
            .I(CLK_EN_c));
    IoInMux I__388 (
            .O(N__4371),
            .I(N__4368));
    LocalMux I__387 (
            .O(N__4368),
            .I(N__4365));
    Odrv12 I__386 (
            .O(N__4365),
            .I(DBRn_c_i_0));
    IoInMux I__385 (
            .O(N__4362),
            .I(N__4359));
    LocalMux I__384 (
            .O(N__4359),
            .I(N__4356));
    Span4Mux_s3_v I__383 (
            .O(N__4356),
            .I(N__4353));
    Span4Mux_h I__382 (
            .O(N__4353),
            .I(N__4350));
    Odrv4 I__381 (
            .O(N__4350),
            .I(CLK80_PLL_i_i));
    IoInMux I__380 (
            .O(N__4347),
            .I(N__4344));
    LocalMux I__379 (
            .O(N__4344),
            .I(N__4341));
    IoSpan4Mux I__378 (
            .O(N__4341),
            .I(N__4338));
    Span4Mux_s2_v I__377 (
            .O(N__4338),
            .I(N__4335));
    Sp12to4 I__376 (
            .O(N__4335),
            .I(N__4332));
    Span12Mux_v I__375 (
            .O(N__4332),
            .I(N__4329));
    Odrv12 I__374 (
            .O(N__4329),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .I(N__4559));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__4561));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__4562));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__4557));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .I(N__4556));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__4558));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .I(N__4563));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_12_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__7796),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__9483),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4371),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__8496),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_11_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_11_5  (
            .in0(N__4442),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11220),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_3_1_1.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_3_1_1.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_3_1_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_3_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10770),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_5_12_7.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_5_12_7.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_5_12_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_5_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4533),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_7_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_7_8_2 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_7_8_2  (
            .in0(N__10152),
            .in1(N__11552),
            .in2(N__4449),
            .in3(N__5738),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .ce(),
            .sr(N__11195));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_7_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_7_9_1 .LUT_INIT=16'b0101000010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_7_9_1  (
            .in0(N__5272),
            .in1(N__7754),
            .in2(N__6420),
            .in3(N__7598),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_7_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_7_11_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_5_LC_7_11_1  (
            .in0(N__10958),
            .in1(_gnd_net_),
            .in2(N__4410),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10753),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_11_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_11_2  (
            .in0(N__6081),
            .in1(N__4419),
            .in2(_gnd_net_),
            .in3(N__4406),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_458_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_11_3 .LUT_INIT=16'b1010001010100000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_11_3  (
            .in0(N__10956),
            .in1(N__8708),
            .in2(N__4413),
            .in3(N__7425),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10753),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_7_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_7_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_4_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__10957),
            .in2(_gnd_net_),
            .in3(N__8625),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10753),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_12_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_12_0  (
            .in0(N__7740),
            .in1(N__7599),
            .in2(N__6418),
            .in3(N__5604),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_7_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_7_12_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_7_12_1 .LUT_INIT=16'b1000110011011100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_7_12_1  (
            .in0(N__5038),
            .in1(N__4382),
            .in2(N__4398),
            .in3(N__4479),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10758),
            .ce(),
            .sr(N__11173));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIN5DI_LC_7_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIN5DI_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIN5DI_LC_7_12_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIN5DI_LC_7_12_2  (
            .in0(N__5232),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5536),
            .lcout(\U712_CHIP_RAM.CLK_EN_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_7_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_7_12_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_7_12_3  (
            .in0(N__8934),
            .in1(N__7739),
            .in2(_gnd_net_),
            .in3(N__5233),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_12_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_12_4  (
            .in0(N__4793),
            .in1(N__5603),
            .in2(N__4485),
            .in3(N__5037),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_442_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_12_5 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_12_5  (
            .in0(N__8935),
            .in1(_gnd_net_),
            .in2(N__4482),
            .in3(N__4478),
            .lcout(\U712_CHIP_RAM.N_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_7_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_7_12_7 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_7_12_7  (
            .in0(N__8936),
            .in1(N__7011),
            .in2(_gnd_net_),
            .in3(N__6219),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10758),
            .ce(),
            .sr(N__11173));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_13_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__4470),
            .in2(_gnd_net_),
            .in3(N__4464),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__4560),
            .ce(),
            .sr(N__4929));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_13_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__5366),
            .in2(_gnd_net_),
            .in3(N__4461),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__4560),
            .ce(),
            .sr(N__4929));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_13_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__5405),
            .in2(_gnd_net_),
            .in3(N__4458),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__4560),
            .ce(),
            .sr(N__4929));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_13_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_13_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__5423),
            .in2(_gnd_net_),
            .in3(N__4455),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__4560),
            .ce(),
            .sr(N__4929));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_13_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_13_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__5384),
            .in2(_gnd_net_),
            .in3(N__4452),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__4560),
            .ce(),
            .sr(N__4929));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_13_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__5111),
            .in2(_gnd_net_),
            .in3(N__4572),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__4560),
            .ce(),
            .sr(N__4929));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_13_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_13_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__5127),
            .in2(_gnd_net_),
            .in3(N__4569),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__4560),
            .ce(),
            .sr(N__4929));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_13_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_13_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__6269),
            .in2(_gnd_net_),
            .in3(N__4566),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4560),
            .ce(),
            .sr(N__4929));
    defparam DBR_SYNC_0_LC_7_14_2.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_7_14_2.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_7_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_7_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4532),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10765),
            .ce(),
            .sr(N__11160));
    defparam DBR_SYNC_1_LC_7_14_6.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_7_14_6.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_7_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_7_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4500),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10765),
            .ce(),
            .sr(N__11160));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNIK9021_0_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNIK9021_0_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNIK9021_0_LC_8_8_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNIK9021_0_LC_8_8_0  (
            .in0(N__10071),
            .in1(N__7996),
            .in2(N__9409),
            .in3(N__10017),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_2_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_2_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_2_LC_8_9_0 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_2_LC_8_9_0  (
            .in0(N__5264),
            .in1(N__4692),
            .in2(N__5640),
            .in3(N__4874),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_8_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_8_9_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_8_9_1  (
            .in0(N__6419),
            .in1(N__4910),
            .in2(N__4731),
            .in3(N__5634),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMDsr_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_8_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_8_9_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_8_9_2  (
            .in0(N__4608),
            .in1(N__4494),
            .in2(N__4488),
            .in3(N__5325),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMDsr_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_9_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_9_3 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_9_3  (
            .in0(N__8011),
            .in1(N__5090),
            .in2(N__4620),
            .in3(N__4617),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10738),
            .ce(),
            .sr(N__11188));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_8_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_8_9_5 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_8_9_5  (
            .in0(N__7595),
            .in1(N__4607),
            .in2(N__5280),
            .in3(N__7753),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMDsr_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_8_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_8_9_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_8_9_6 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_8_9_6  (
            .in0(N__5091),
            .in1(N__4632),
            .in2(N__4611),
            .in3(N__10078),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10738),
            .ce(),
            .sr(N__11188));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_8_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_8_10_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_8_10_0  (
            .in0(N__5637),
            .in1(N__7745),
            .in2(N__5278),
            .in3(N__7592),
            .lcout(\U712_CHIP_RAM.N_433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_10_2 .LUT_INIT=16'b1011110110011101;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_10_2  (
            .in0(N__5639),
            .in1(N__7746),
            .in2(N__5279),
            .in3(N__6312),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_4_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_3 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_3  (
            .in0(N__7594),
            .in1(N__5042),
            .in2(N__4599),
            .in3(N__5064),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_173_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_10_4 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_8_10_4  (
            .in0(N__4596),
            .in1(N__11010),
            .in2(N__4587),
            .in3(N__8803),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10743),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_10_5 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_LC_8_10_5  (
            .in0(N__9025),
            .in1(N__7956),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_8_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_8_10_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_8_10_6  (
            .in0(N__5638),
            .in1(N__7744),
            .in2(_gnd_net_),
            .in3(N__5040),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMDsr_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_8_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_8_10_7 .LUT_INIT=16'b1111001111110111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_8_10_7  (
            .in0(N__7593),
            .in1(N__5169),
            .in2(N__4635),
            .in3(N__5321),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILL5O1_0_LC_8_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILL5O1_0_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILL5O1_0_LC_8_11_0 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNILL5O1_0_LC_8_11_0  (
            .in0(N__6378),
            .in1(N__7590),
            .in2(N__5257),
            .in3(N__7697),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIC9HD1_LC_8_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIC9HD1_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIC9HD1_LC_8_11_1 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIC9HD1_LC_8_11_1  (
            .in0(N__5593),
            .in1(N__7691),
            .in2(_gnd_net_),
            .in3(N__7408),
            .lcout(\U712_CHIP_RAM.N_327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_11_2  (
            .in0(N__4866),
            .in1(N__4902),
            .in2(N__4691),
            .in3(N__4722),
            .lcout(\U712_CHIP_RAM.N_301 ),
            .ltout(\U712_CHIP_RAM.N_301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_8_11_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_8_11_3  (
            .in0(N__5592),
            .in1(_gnd_net_),
            .in2(N__4626),
            .in3(N__5224),
            .lcout(\U712_CHIP_RAM.N_534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_0_LC_8_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_0_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_0_LC_8_11_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_0_LC_8_11_4  (
            .in0(N__4686),
            .in1(N__4723),
            .in2(_gnd_net_),
            .in3(N__5594),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_8_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_8_11_5 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_8_11_5  (
            .in0(N__5595),
            .in1(N__5229),
            .in2(_gnd_net_),
            .in3(N__5039),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMDsr_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_11_6 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_11_6  (
            .in0(N__4773),
            .in1(N__7591),
            .in2(N__4623),
            .in3(N__5076),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_LC_8_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_LC_8_11_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__5225),
            .in2(_gnd_net_),
            .in3(N__6377),
            .lcout(\U712_CHIP_RAM.N_300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_12_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_12_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__6397),
            .in2(_gnd_net_),
            .in3(N__8720),
            .lcout(\U712_CHIP_RAM.LATCH_CLK_6 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_12_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_12_1  (
            .in0(N__5158),
            .in1(N__5250),
            .in2(_gnd_net_),
            .in3(N__4740),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__10754),
            .ce(N__5297),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_12_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__7730),
            .in2(_gnd_net_),
            .in3(N__4737),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_12_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_12_3  (
            .in0(N__5159),
            .in1(N__5605),
            .in2(_gnd_net_),
            .in3(N__4734),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__10754),
            .ce(N__5297),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_12_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_12_4  (
            .in0(N__5153),
            .in1(N__4727),
            .in2(_gnd_net_),
            .in3(N__4704),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__10754),
            .ce(N__5297),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_12_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_12_5  (
            .in0(N__5160),
            .in1(N__4909),
            .in2(_gnd_net_),
            .in3(N__4701),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__10754),
            .ce(N__5297),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_12_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_12_6  (
            .in0(N__5154),
            .in1(N__4873),
            .in2(_gnd_net_),
            .in3(N__4698),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__10754),
            .ce(N__5297),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_12_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_12_7  (
            .in0(N__4690),
            .in1(N__5155),
            .in2(_gnd_net_),
            .in3(N__4695),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10754),
            .ce(N__5297),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_13_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_13_0  (
            .in0(N__4797),
            .in1(N__5498),
            .in2(N__7738),
            .in3(N__7545),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_396_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_8_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_8_13_1 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_8_13_1  (
            .in0(N__11006),
            .in1(N__4665),
            .in2(N__4659),
            .in3(N__4646),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10759),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_8_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_8_13_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__5534),
            .in2(_gnd_net_),
            .in3(N__6379),
            .lcout(\U712_CHIP_RAM.N_315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_13_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_13_4  (
            .in0(N__6154),
            .in1(N__10556),
            .in2(_gnd_net_),
            .in3(N__7439),
            .lcout(\U712_CHIP_RAM.N_336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIU7TF5_LC_8_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIU7TF5_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIU7TF5_LC_8_13_5 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIU7TF5_LC_8_13_5  (
            .in0(N__7438),
            .in1(N__6099),
            .in2(N__6456),
            .in3(N__5979),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_8_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_8_13_6 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_8_13_6  (
            .in0(N__5535),
            .in1(N__11007),
            .in2(N__4782),
            .in3(N__4779),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10759),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_13_7 .LUT_INIT=16'b1010100110101011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_13_7  (
            .in0(N__6383),
            .in1(N__5231),
            .in2(N__7583),
            .in3(N__7698),
            .lcout(\U712_CHIP_RAM.N_372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_8_14_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_8_14_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__11008),
            .in2(_gnd_net_),
            .in3(N__5436),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10762),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_8_15_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_8_15_0 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_8_15_0  (
            .in0(N__11009),
            .in1(N__6067),
            .in2(_gnd_net_),
            .in3(N__7215),
            .lcout(\U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_7_1 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_7_1  (
            .in0(N__8012),
            .in1(N__9406),
            .in2(_gnd_net_),
            .in3(N__10028),
            .lcout(\U712_CHIP_RAM.CMA_5_i_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_9_8_2 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_9_8_2  (
            .in0(N__8389),
            .in1(N__8037),
            .in2(N__6900),
            .in3(N__5724),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10731),
            .ce(N__8293),
            .sr(N__11189));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_9_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_9_8_4 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_9_8_4  (
            .in0(N__4968),
            .in1(N__4962),
            .in2(N__9056),
            .in3(N__8028),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10731),
            .ce(N__8293),
            .sr(N__11189));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIDBLK1_3_LC_9_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIDBLK1_3_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIDBLK1_3_LC_9_8_7 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIDBLK1_3_LC_9_8_7  (
            .in0(N__7997),
            .in1(N__4925),
            .in2(N__9410),
            .in3(N__10072),
            .lcout(\U712_CHIP_RAM.un1_CMA25_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__7742),
            .in2(_gnd_net_),
            .in3(N__7379),
            .lcout(\U712_CHIP_RAM.DBENn_7_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_0_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_0_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_0_LC_9_9_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_0_LC_9_9_1  (
            .in0(N__5508),
            .in1(N__4911),
            .in2(N__4881),
            .in3(N__4845),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_0_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_0_LC_9_9_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_0_LC_9_9_2 .LUT_INIT=16'b1111001011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_0_LC_9_9_2  (
            .in0(N__7596),
            .in1(N__7743),
            .in2(N__4836),
            .in3(N__5271),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10734),
            .ce(N__4818),
            .sr(N__11184));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1DB24_2_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1DB24_2_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1DB24_2_LC_9_10_1 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI1DB24_2_LC_9_10_1  (
            .in0(N__6182),
            .in1(N__7741),
            .in2(N__4833),
            .in3(N__5063),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI2MHHA_2_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI2MHHA_2_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI2MHHA_2_LC_9_10_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI2MHHA_2_LC_9_10_2  (
            .in0(N__5550),
            .in1(N__5049),
            .in2(N__4824),
            .in3(N__5041),
            .lcout(\U712_CHIP_RAM.N_191 ),
            .ltout(\U712_CHIP_RAM.N_191_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_0_LC_9_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_0_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_0_LC_9_10_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_0_LC_9_10_3  (
            .in0(N__11219),
            .in1(_gnd_net_),
            .in2(N__4821),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_191_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_9_10_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_9_10_5  (
            .in0(N__4812),
            .in1(N__4995),
            .in2(_gnd_net_),
            .in3(N__7003),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10739),
            .ce(),
            .sr(N__11174));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_10_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_10_6 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_10_6  (
            .in0(N__5097),
            .in1(N__5089),
            .in2(N__9408),
            .in3(N__5352),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10739),
            .ce(),
            .sr(N__11174));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7FAQ2_3_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7FAQ2_3_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7FAQ2_3_LC_9_10_7 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI7FAQ2_3_LC_9_10_7  (
            .in0(N__5635),
            .in1(N__5075),
            .in2(_gnd_net_),
            .in3(N__5062),
            .lcout(\U712_CHIP_RAM.N_370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_9_11_0 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_9_11_0  (
            .in0(N__6183),
            .in1(N__10954),
            .in2(N__7443),
            .in3(N__5978),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_0_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_0_LC_9_11_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_0_LC_9_11_1  (
            .in0(N__5591),
            .in1(N__6375),
            .in2(N__5043),
            .in3(N__5230),
            .lcout(\U712_CHIP_RAM.N_466 ),
            .ltout(\U712_CHIP_RAM.N_466_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_9_11_2 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_9_11_2  (
            .in0(N__7692),
            .in1(_gnd_net_),
            .in2(N__5001),
            .in3(N__7578),
            .lcout(\U712_CHIP_RAM.N_471 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_9_11_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__5540),
            .in2(_gnd_net_),
            .in3(N__6376),
            .lcout(\U712_CHIP_RAM.N_299 ),
            .ltout(\U712_CHIP_RAM.N_299_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_9_11_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_9_11_4  (
            .in0(N__7693),
            .in1(N__7579),
            .in2(N__4998),
            .in3(N__5481),
            .lcout(\U712_CHIP_RAM.N_429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_11_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_11_5  (
            .in0(N__4994),
            .in1(N__4983),
            .in2(_gnd_net_),
            .in3(N__9356),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_11_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_11_6  (
            .in0(N__7694),
            .in1(N__7580),
            .in2(_gnd_net_),
            .in3(N__7371),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_399_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_11_7 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_11_7  (
            .in0(N__10955),
            .in1(N__5497),
            .in2(N__5430),
            .in3(N__6300),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_12_1 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_12_1  (
            .in0(N__5427),
            .in1(N__5409),
            .in2(N__5391),
            .in3(N__5370),
            .lcout(\U712_CHIP_RAM.REFRESH5lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_12_2 .LUT_INIT=16'b0011000011000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_12_2  (
            .in0(N__6243),
            .in1(N__7547),
            .in2(N__5277),
            .in3(N__7708),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_12_3 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_12_3  (
            .in0(N__11000),
            .in1(N__5156),
            .in2(N__5340),
            .in3(N__5331),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10748),
            .ce(N__5298),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_0_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_0_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_0_LC_9_12_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_0_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__7707),
            .in2(_gnd_net_),
            .in3(N__6385),
            .lcout(\U712_CHIP_RAM.N_310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_12_5 .LUT_INIT=16'b0001001011011110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_12_5  (
            .in0(N__5870),
            .in1(N__5157),
            .in2(N__6404),
            .in3(N__5304),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10748),
            .ce(N__5298),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_12_6 .LUT_INIT=16'b1111100111111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_12_6  (
            .in0(N__5636),
            .in1(N__6384),
            .in2(N__5276),
            .in3(N__7546),
            .lcout(\U712_CHIP_RAM.N_385 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_9_13_0 .LUT_INIT=16'b1111110111011101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_9_13_0  (
            .in0(N__11002),
            .in1(N__6279),
            .in2(N__6296),
            .in3(N__5493),
            .lcout(\U712_CHIP_RAM.N_182 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_13_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__5126),
            .in2(_gnd_net_),
            .in3(N__5112),
            .lcout(\U712_CHIP_RAM.REFRESH5lto7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_9_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_9_13_2 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_9_13_2  (
            .in0(N__11003),
            .in1(N__5596),
            .in2(N__7582),
            .in3(N__7695),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_0_LC_9_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_0_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_0_LC_9_13_4 .LUT_INIT=16'b1010101010110001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_0_LC_9_13_4  (
            .in0(N__7540),
            .in1(N__7696),
            .in2(N__5541),
            .in3(N__6389),
            .lcout(\U712_CHIP_RAM.N_382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_13_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_13_5  (
            .in0(N__6390),
            .in1(N__7541),
            .in2(N__5499),
            .in3(N__7737),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_13_6 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__11001),
            .in2(N__5466),
            .in3(N__7556),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10755),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_14_0 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_14_0  (
            .in0(N__7905),
            .in1(N__7191),
            .in2(N__9210),
            .in3(N__7236),
            .lcout(),
            .ltout(\U712_REG_SM.N_411_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_14_1 .LUT_INIT=16'b0000101000000010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_9_14_1  (
            .in0(N__11005),
            .in1(N__9209),
            .in2(N__5463),
            .in3(N__9621),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10760),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_9_14_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_9_14_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_9_14_3  (
            .in0(N__11872),
            .in1(N__8766),
            .in2(_gnd_net_),
            .in3(N__8724),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_446_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_52_i_LC_9_14_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_52_i_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_52_i_LC_9_14_4 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \U712_BYTE_ENABLE.N_52_i_LC_9_14_4  (
            .in0(N__7146),
            .in1(N__7158),
            .in2(N__5460),
            .in3(N__9800),
            .lcout(N_52_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_9_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_9_14_5 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_9_14_5  (
            .in0(N__11004),
            .in1(N__11873),
            .in2(_gnd_net_),
            .in3(N__11927),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10760),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_9_15_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_9_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__6513),
            .in2(N__6558),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBR_COUNT_2_LC_9_15_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_2_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_2_LC_9_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_2_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__6527),
            .in2(_gnd_net_),
            .in3(N__5658),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_1 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_2 ),
            .clk(N__10763),
            .ce(),
            .sr(N__5888));
    defparam \U712_CHIP_RAM.DBR_COUNT_3_LC_9_15_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_3_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_3_LC_9_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_3_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__6791),
            .in2(_gnd_net_),
            .in3(N__5655),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_2 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_3 ),
            .clk(N__10763),
            .ce(),
            .sr(N__5888));
    defparam \U712_CHIP_RAM.DBR_COUNT_4_LC_9_15_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_4_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_4_LC_9_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_4_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__6804),
            .in2(_gnd_net_),
            .in3(N__5652),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_3 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_4 ),
            .clk(N__10763),
            .ce(),
            .sr(N__5888));
    defparam \U712_CHIP_RAM.DBR_COUNT_5_LC_9_15_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_5_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_5_LC_9_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_5_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__6816),
            .in2(_gnd_net_),
            .in3(N__5649),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_4 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_5 ),
            .clk(N__10763),
            .ce(),
            .sr(N__5888));
    defparam \U712_CHIP_RAM.DBR_COUNT_6_LC_9_15_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_6_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_6_LC_9_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_6_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__6540),
            .in2(_gnd_net_),
            .in3(N__5646),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_5 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_6 ),
            .clk(N__10763),
            .ce(),
            .sr(N__5888));
    defparam \U712_CHIP_RAM.DBR_COUNT_7_LC_9_15_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_COUNT_7_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_7_LC_9_15_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_7_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__6777),
            .in2(_gnd_net_),
            .in3(N__5643),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10763),
            .ce(),
            .sr(N__5888));
    defparam \U712_CHIP_RAM.DBR_COUNT_1_LC_9_15_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_COUNT_1_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_1_LC_9_15_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_1_LC_9_15_7  (
            .in0(N__6514),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6557),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10763),
            .ce(),
            .sr(N__5888));
    defparam \U712_CHIP_RAM.DBR_COUNT_0_LC_9_16_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_COUNT_0_LC_9_16_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_0_LC_9_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_0_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6516),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10766),
            .ce(),
            .sr(N__5889));
    defparam CONSTANT_ONE_LUT4_LC_10_2_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_2_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_2_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_10_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_10_7_2 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_10_7_2  (
            .in0(N__5703),
            .in1(N__8390),
            .in2(N__9447),
            .in3(N__6171),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10722),
            .ce(N__8290),
            .sr(N__11190));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_8_2  (
            .in0(N__5804),
            .in1(N__5924),
            .in2(_gnd_net_),
            .in3(N__9439),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_8_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_8_3  (
            .in0(N__9440),
            .in1(N__9038),
            .in2(N__5769),
            .in3(N__9267),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_8_5  (
            .in0(N__9438),
            .in1(N__5678),
            .in2(_gnd_net_),
            .in3(N__5766),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_8_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_8_6  (
            .in0(N__9037),
            .in1(N__9441),
            .in2(N__5742),
            .in3(N__5739),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_7  (
            .in0(N__5718),
            .in1(N__9036),
            .in2(_gnd_net_),
            .in3(N__9960),
            .lcout(\U712_CHIP_RAM.N_353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_9_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_9_0  (
            .in0(N__5697),
            .in1(N__11531),
            .in2(N__5682),
            .in3(N__7007),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10732),
            .ce(),
            .sr(N__11175));
    defparam \U712_CHIP_RAM.DBENn_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_10_9_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_10_9_3 .LUT_INIT=16'b0010111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_10_9_3  (
            .in0(N__8745),
            .in1(N__6201),
            .in2(N__5667),
            .in3(N__9969),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10732),
            .ce(),
            .sr(N__11175));
    defparam \U712_CHIP_RAM.DBDIR_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_10_9_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_10_9_4 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_10_9_4  (
            .in0(N__6162),
            .in1(N__6038),
            .in2(_gnd_net_),
            .in3(N__6114),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10732),
            .ce(),
            .sr(N__11175));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI3LH42_3_LC_10_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI3LH42_3_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI3LH42_3_LC_10_9_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI3LH42_3_LC_10_9_6  (
            .in0(N__11218),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6027),
            .lcout(\U712_CHIP_RAM.un1_CMA25_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_1  (
            .in0(N__6021),
            .in1(N__5987),
            .in2(_gnd_net_),
            .in3(N__9344),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_10_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_10_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_10_10_2  (
            .in0(N__5988),
            .in1(N__6006),
            .in2(_gnd_net_),
            .in3(N__7001),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10735),
            .ce(),
            .sr(N__11168));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIU7TF5_0_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIU7TF5_0_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIU7TF5_0_LC_10_10_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIU7TF5_0_LC_10_10_4  (
            .in0(N__6449),
            .in1(N__6092),
            .in2(N__7450),
            .in3(N__5974),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_10_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_10_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_10_10_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__5958),
            .in2(N__5943),
            .in3(N__8162),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10735),
            .ce(),
            .sr(N__11168));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_10_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_10_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_10_10_6  (
            .in0(N__5925),
            .in1(N__5940),
            .in2(_gnd_net_),
            .in3(N__7000),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10735),
            .ce(),
            .sr(N__11168));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_10_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_10_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_10_10_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_10_10_7  (
            .in0(N__7002),
            .in1(N__5907),
            .in2(_gnd_net_),
            .in3(N__8123),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10735),
            .ce(),
            .sr(N__11168));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_11_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_11_0  (
            .in0(N__7719),
            .in1(N__7367),
            .in2(N__7451),
            .in3(N__7581),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_10_11_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6222),
            .in3(N__6215),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_11_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6192),
            .in3(N__11217),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_11_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_11_3  (
            .in0(N__9004),
            .in1(N__6189),
            .in2(N__9407),
            .in3(N__10101),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_11_4 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_11_4  (
            .in0(N__6241),
            .in1(N__6571),
            .in2(_gnd_net_),
            .in3(N__6441),
            .lcout(\U712_CHIP_RAM.N_319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_11_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_11_5  (
            .in0(N__9003),
            .in1(N__7074),
            .in2(_gnd_net_),
            .in3(N__9930),
            .lcout(\U712_CHIP_RAM.N_359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_10_11_6 .LUT_INIT=16'b0101000011000000;
    LogicCell40 \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_10_11_6  (
            .in0(N__6161),
            .in1(N__10600),
            .in2(N__10877),
            .in3(N__6113),
            .lcout(DMA_WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10740),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIFGNH_LC_10_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIFGNH_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIFGNH_LC_10_11_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIFGNH_LC_10_11_7  (
            .in0(N__6572),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6242),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_12_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_12_0  (
            .in0(N__7241),
            .in1(N__10943),
            .in2(N__6492),
            .in3(N__6080),
            .lcout(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10744),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_10_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_10_12_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__8990),
            .in2(_gnd_net_),
            .in3(N__6448),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_419_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_12_4 .LUT_INIT=16'b1100000011000100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_12_4  (
            .in0(N__7313),
            .in1(N__10942),
            .in2(N__6477),
            .in3(N__6474),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10744),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_10_12_5 .LUT_INIT=16'b0110010000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_10_12_5  (
            .in0(N__7709),
            .in1(N__7548),
            .in2(N__6414),
            .in3(N__6311),
            .lcout(\U712_CHIP_RAM.N_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_12_6 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_12_6  (
            .in0(N__7549),
            .in1(N__7710),
            .in2(_gnd_net_),
            .in3(N__7378),
            .lcout(\U712_CHIP_RAM.N_434 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_10_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_12_7 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_10_12_7  (
            .in0(N__6273),
            .in1(N__6255),
            .in2(N__10996),
            .in3(N__6249),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10744),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_10_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_10_13_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(N__7182),
            .in2(_gnd_net_),
            .in3(N__9139),
            .lcout(\U712_REG_SM.N_322 ),
            .ltout(\U712_REG_SM.N_322_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_13_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_13_1  (
            .in0(N__9237),
            .in1(N__7277),
            .in2(N__6228),
            .in3(N__7903),
            .lcout(\U712_REG_SM.N_410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_13_2 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_13_2  (
            .in0(N__9605),
            .in1(N__9236),
            .in2(_gnd_net_),
            .in3(N__9198),
            .lcout(\U712_REG_SM.N_367 ),
            .ltout(\U712_REG_SM.N_367_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_3 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(N__6644),
            .in2(N__6225),
            .in3(N__7904),
            .lcout(\U712_REG_SM.N_131 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_RNO_0_LC_10_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_RNO_0_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REGENn_RNO_0_LC_10_13_5 .LUT_INIT=16'b0101000000100010;
    LogicCell40 \U712_REG_SM.REGENn_RNO_0_LC_10_13_5  (
            .in0(N__9199),
            .in1(N__7278),
            .in2(N__9147),
            .in3(N__6610),
            .lcout(\U712_REG_SM.REGENn_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_10_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_10_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_10_13_6  (
            .in0(N__9606),
            .in1(N__7183),
            .in2(N__7242),
            .in3(N__9200),
            .lcout(),
            .ltout(\U712_REG_SM.N_408_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_10_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_10_13_7 .LUT_INIT=16'b1110110011100100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_10_13_7  (
            .in0(N__10948),
            .in1(N__7948),
            .in2(N__6660),
            .in3(N__6657),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10749),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_10_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_10_14_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_10_14_0 .LUT_INIT=16'b1100110011001101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_10_14_0  (
            .in0(N__6594),
            .in1(N__6651),
            .in2(N__7911),
            .in3(N__7965),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10756),
            .ce(),
            .sr(N__11156));
    defparam \U712_REG_SM.WRITE_CYCLE_LC_10_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_10_14_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_10_14_1 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_REG_SM.WRITE_CYCLE_LC_10_14_1  (
            .in0(N__10579),
            .in1(N__6645),
            .in2(_gnd_net_),
            .in3(N__8446),
            .lcout(\U712_REG_SM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10756),
            .ce(),
            .sr(N__11156));
    defparam \U712_REG_SM.REGENn_LC_10_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_10_14_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_10_14_2 .LUT_INIT=16'b1010011010100010;
    LogicCell40 \U712_REG_SM.REGENn_LC_10_14_2  (
            .in0(N__6611),
            .in1(N__6633),
            .in2(N__9618),
            .in3(N__7254),
            .lcout(REGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10756),
            .ce(),
            .sr(N__11156));
    defparam \U712_REG_SM.REG_TACK_LC_10_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_10_14_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_10_14_4  (
            .in0(N__6593),
            .in1(N__7875),
            .in2(N__8847),
            .in3(N__6585),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10756),
            .ce(),
            .sr(N__11156));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_10_15_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_10_15_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_10_15_0  (
            .in0(N__6579),
            .in1(N__6553),
            .in2(_gnd_net_),
            .in3(N__6539),
            .lcout(),
            .ltout(\U712_CHIP_RAM.RAM_CYCLE_DISABLE_5_i_a2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_10_15_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_10_15_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_10_15_1  (
            .in0(N__6528),
            .in1(N__6515),
            .in2(N__6495),
            .in3(N__6765),
            .lcout(\U712_CHIP_RAM.N_456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_15_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_15_4 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_15_4  (
            .in0(N__10463),
            .in1(N__9868),
            .in2(_gnd_net_),
            .in3(N__9011),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_10_15_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_10_15_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_10_15_5  (
            .in0(N__6815),
            .in1(N__6803),
            .in2(N__6792),
            .in3(N__6776),
            .lcout(\U712_CHIP_RAM.RAM_CYCLE_DISABLE_5_i_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_10_15_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_10_15_7 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_10_15_7  (
            .in0(N__9012),
            .in1(N__10464),
            .in2(_gnd_net_),
            .in3(N__10421),
            .lcout(\U712_BYTE_ENABLE.N_424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_RNO_0_LC_10_16_2 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_10_16_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_REG_SM.LDSn_RNO_0_LC_10_16_2  (
            .in0(N__9835),
            .in1(N__10405),
            .in2(N__10575),
            .in3(N__10500),
            .lcout(\U712_REG_SM.N_402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_10_19_6 .C_ON=1'b0;
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_10_19_6 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_10_19_6  (
            .in0(N__11868),
            .in1(N__11919),
            .in2(_gnd_net_),
            .in3(N__10619),
            .lcout(DMA_LATCH_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_11_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_11_7_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_11_7_3  (
            .in0(N__8391),
            .in1(N__10092),
            .in2(_gnd_net_),
            .in3(N__9417),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10720),
            .ce(N__8292),
            .sr(N__11185));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_8_0  (
            .in0(N__6719),
            .in1(N__7044),
            .in2(_gnd_net_),
            .in3(N__9419),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_8_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_8_1  (
            .in0(N__9035),
            .in1(N__9442),
            .in2(N__6684),
            .in3(N__9981),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_8_2 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_11_8_2  (
            .in0(N__6879),
            .in1(N__8377),
            .in2(N__6681),
            .in3(N__11298),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10723),
            .ce(N__8300),
            .sr(N__11176));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_11_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_11_8_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__9034),
            .in2(_gnd_net_),
            .in3(N__9418),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_8_5 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_11_8_5  (
            .in0(N__10314),
            .in1(N__8378),
            .in2(N__6894),
            .in3(N__7110),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10723),
            .ce(N__8300),
            .sr(N__11176));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_11_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_11_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_11_9_2  (
            .in0(N__7005),
            .in1(N__7092),
            .in2(_gnd_net_),
            .in3(N__7073),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10728),
            .ce(),
            .sr(N__11169));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_11_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_11_9_3  (
            .in0(N__7059),
            .in1(N__7043),
            .in2(_gnd_net_),
            .in3(N__7004),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10728),
            .ce(),
            .sr(N__11169));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_11_9_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_11_9_5  (
            .in0(N__7029),
            .in1(N__8226),
            .in2(_gnd_net_),
            .in3(N__7006),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10728),
            .ce(),
            .sr(N__11169));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_10_2 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_11_10_2  (
            .in0(N__8375),
            .in1(N__6892),
            .in2(N__10254),
            .in3(N__8106),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10733),
            .ce(N__8301),
            .sr(N__11161));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_11_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_11_10_3 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_11_10_3  (
            .in0(N__8373),
            .in1(N__9255),
            .in2(N__6898),
            .in3(N__8631),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10733),
            .ce(N__8301),
            .sr(N__11161));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_10_6 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_11_10_6  (
            .in0(N__8376),
            .in1(N__6893),
            .in2(N__9948),
            .in3(N__8211),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10733),
            .ce(N__8301),
            .sr(N__11161));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_10_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_11_10_7  (
            .in0(N__8374),
            .in1(N__9246),
            .in2(N__6899),
            .in3(N__6846),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10733),
            .ce(N__8301),
            .sr(N__11161));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_11_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_11_0  (
            .in0(N__7755),
            .in1(N__7597),
            .in2(N__7452),
            .in3(N__7380),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10736),
            .ce(N__7341),
            .sr(N__11157));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_11_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_11_12_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__8429),
            .in2(_gnd_net_),
            .in3(N__7276),
            .lcout(),
            .ltout(\U712_REG_SM.N_401_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_11_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_11_12_1 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_11_12_1  (
            .in0(N__7335),
            .in1(N__7314),
            .in2(N__7281),
            .in3(N__10941),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10741),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_11_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_11_13_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_11_13_2  (
            .in0(N__7270),
            .in1(N__9192),
            .in2(N__9619),
            .in3(N__7253),
            .lcout(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_11_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_11_13_3 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_11_13_3  (
            .in0(N__9194),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7237),
            .lcout(),
            .ltout(\U712_REG_SM.N_324_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_11_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_11_13_4 .LUT_INIT=16'b0010000000100010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_11_13_4  (
            .in0(N__10947),
            .in1(N__7164),
            .in2(N__7194),
            .in3(N__9613),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10745),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_11_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_11_13_6 .LUT_INIT=16'b0000000011111101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_11_13_6  (
            .in0(N__9143),
            .in1(N__9193),
            .in2(N__9620),
            .in3(N__7187),
            .lcout(\U712_REG_SM.STATE_COUNTc_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_170_i_LC_11_14_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_170_i_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_170_i_LC_11_14_0 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \U712_BYTE_ENABLE.N_170_i_LC_11_14_0  (
            .in0(N__7157),
            .in1(N__9801),
            .in2(N__8673),
            .in3(N__7145),
            .lcout(N_170_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_14_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__9197),
            .in2(_gnd_net_),
            .in3(N__9593),
            .lcout(),
            .ltout(\U712_REG_SM.N_325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_14_2 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_11_14_2  (
            .in0(N__10959),
            .in1(N__8448),
            .in2(N__7968),
            .in3(N__9145),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10750),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_14_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_14_3 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_14_3  (
            .in0(N__9234),
            .in1(N__9196),
            .in2(_gnd_net_),
            .in3(N__9592),
            .lcout(\U712_REG_SM.N_302 ),
            .ltout(\U712_REG_SM.N_302_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_14_4 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_11_14_4  (
            .in0(N__10960),
            .in1(N__7910),
            .in2(N__7959),
            .in3(N__9235),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10750),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.N_160_i_LC_11_14_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_160_i_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_160_i_LC_11_14_5 .LUT_INIT=16'b0101010001010000;
    LogicCell40 \U712_BUFFERS.N_160_i_LC_11_14_5  (
            .in0(N__7949),
            .in1(N__11952),
            .in2(N__9055),
            .in3(N__11874),
            .lcout(N_160_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_11_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_11_14_7 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_11_14_7  (
            .in0(N__7909),
            .in1(N__9195),
            .in2(_gnd_net_),
            .in3(N__9591),
            .lcout(\U712_REG_SM.N_404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_11_15_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_11_15_1 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_11_15_1 .LUT_INIT=16'b1111100011111100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_11_15_1  (
            .in0(N__9101),
            .in1(N__7815),
            .in2(N__8664),
            .in3(N__9724),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10757),
            .ce(),
            .sr(N__11154));
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_15_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_15_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7797),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10757),
            .ce(),
            .sr(N__11154));
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_15_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7761),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10757),
            .ce(),
            .sr(N__11154));
    defparam \U712_REG_SM.ASn_ess_RNO_LC_11_16_0 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_11_16_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U712_REG_SM.ASn_ess_RNO_LC_11_16_0  (
            .in0(N__9529),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11216),
            .lcout(\U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_16_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_16_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_16_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_11_16_4  (
            .in0(N__10998),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8100),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10761),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_16_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_16_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__8659),
            .in2(_gnd_net_),
            .in3(N__8099),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_16_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_16_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_11_16_7  (
            .in0(N__9729),
            .in1(_gnd_net_),
            .in2(N__9105),
            .in3(N__10997),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10761),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_LC_11_17_0 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_LC_11_17_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_ess_LC_11_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.ASn_ess_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9617),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10764),
            .ce(N__8067),
            .sr(N__11150));
    defparam \U712_CHIP_RAM.RASn_LC_12_2_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_12_2_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_12_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_12_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8019),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10718),
            .ce(),
            .sr(N__11197));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_8_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_8_0  (
            .in0(N__11733),
            .in1(N__11548),
            .in2(_gnd_net_),
            .in3(N__10147),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11286),
            .ce(N__11255),
            .sr(N__11167));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_8_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_8_1  (
            .in0(N__10148),
            .in1(_gnd_net_),
            .in2(N__11553),
            .in3(N__11042),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11286),
            .ce(N__11255),
            .sr(N__11167));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNIE8IL_0_LC_12_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNIE8IL_0_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNIE8IL_0_LC_12_9_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNIE8IL_0_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__8010),
            .in2(_gnd_net_),
            .in3(N__10027),
            .lcout(\U712_CHIP_RAM.N_309 ),
            .ltout(\U712_CHIP_RAM.N_309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_9_4 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_9_4  (
            .in0(N__9043),
            .in1(N__11792),
            .in2(N__7971),
            .in3(N__9448),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_9_6 .LUT_INIT=16'b0100000000001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_9_6  (
            .in0(N__9044),
            .in1(N__11793),
            .in2(N__8388),
            .in3(N__9449),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_9_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(N__8322),
            .in2(N__8316),
            .in3(N__8145),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10721),
            .ce(N__8291),
            .sr(N__11159));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_0  (
            .in0(N__8241),
            .in1(N__8225),
            .in2(_gnd_net_),
            .in3(N__9452),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_10_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_10_1  (
            .in0(N__9455),
            .in1(N__9047),
            .in2(N__8214),
            .in3(N__11685),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_10_2  (
            .in0(N__8195),
            .in1(N__8163),
            .in2(_gnd_net_),
            .in3(N__9450),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_10_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_10_3  (
            .in0(N__9453),
            .in1(N__9045),
            .in2(N__8148),
            .in3(N__11565),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_10_4  (
            .in0(N__8139),
            .in1(N__8124),
            .in2(_gnd_net_),
            .in3(N__9451),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_10_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_10_5  (
            .in0(N__9454),
            .in1(N__9046),
            .in2(N__8109),
            .in3(N__10164),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_11_0 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_11_0  (
            .in0(N__9039),
            .in1(N__8643),
            .in2(N__9446),
            .in3(N__9936),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_12_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_12_11_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_3_LC_12_11_3  (
            .in0(N__10840),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10779),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10730),
            .ce(),
            .sr(_gnd_net_));
    defparam pll_RNI8MQ3_LC_12_12_4.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_12_12_4.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_12_12_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 pll_RNI8MQ3_LC_12_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9097),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_LC_12_13_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_12_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_12_13_1 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_LC_12_13_1  (
            .in0(N__9684),
            .in1(N__8514),
            .in2(_gnd_net_),
            .in3(N__8859),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10737),
            .ce(),
            .sr(N__11155));
    defparam \U712_REG_SM.C3_SYNC_0_LC_12_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_12_13_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_12_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8477),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10737),
            .ce(),
            .sr(N__11155));
    defparam \U712_REG_SM.C3_SYNC_1_LC_12_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_12_13_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_12_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8454),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10737),
            .ce(),
            .sr(N__11155));
    defparam \U712_REG_SM.START_RST_LC_12_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.START_RST_LC_12_13_6 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_REG_SM.START_RST_LC_12_13_6  (
            .in0(N__8430),
            .in1(N__8447),
            .in2(_gnd_net_),
            .in3(N__9144),
            .lcout(\U712_REG_SM.START_RSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10737),
            .ce(),
            .sr(N__11155));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_12_14_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_12_14_0 .LUT_INIT=16'b0010111100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_12_14_0  (
            .in0(N__9789),
            .in1(N__9869),
            .in2(N__9921),
            .in3(N__9051),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_443_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_54_i_LC_12_14_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_54_i_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_54_i_LC_12_14_1 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \U712_BYTE_ENABLE.N_54_i_LC_12_14_1  (
            .in0(N__8779),
            .in1(N__11951),
            .in2(N__8418),
            .in3(N__8722),
            .lcout(N_54_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_12_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_12_14_2 .LUT_INIT=16'b1101110111001111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_12_14_2  (
            .in0(N__9228),
            .in1(N__9181),
            .in2(N__9146),
            .in3(N__9577),
            .lcout(\U712_REG_SM.un1_REGENn_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_14_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_14_3 .LUT_INIT=16'b0000000000110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_14_3  (
            .in0(N__8814),
            .in1(N__9668),
            .in2(N__8853),
            .in3(N__9720),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_452_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_14_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_14_4 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_12_14_4  (
            .in0(N__9669),
            .in1(N__10961),
            .in2(N__9108),
            .in3(N__9096),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10742),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_12_14_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_12_14_5 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_12_14_5  (
            .in0(N__9870),
            .in1(N__9790),
            .in2(N__9057),
            .in3(N__9920),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_421_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_168_i_LC_12_14_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_168_i_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_168_i_LC_12_14_6 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \U712_BYTE_ENABLE.N_168_i_LC_12_14_6  (
            .in0(N__8721),
            .in1(N__11950),
            .in2(N__8883),
            .in3(N__8778),
            .lcout(N_168_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_12_14_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_12_14_7 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_12_14_7  (
            .in0(N__8813),
            .in1(N__8849),
            .in2(_gnd_net_),
            .in3(N__9667),
            .lcout(\U712_CYCLE_TERM.N_326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_15_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_15_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__8848),
            .in2(_gnd_net_),
            .in3(N__8812),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_12_15_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_12_15_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_12_15_1  (
            .in0(N__11850),
            .in1(N__8780),
            .in2(_gnd_net_),
            .in3(N__8723),
            .lcout(\U712_BYTE_ENABLE.N_425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_12_15_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_12_15_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_12_15_4  (
            .in0(N__10962),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8663),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10747),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_12_16_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_12_16_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_12_16_0 .LUT_INIT=16'b0101010101000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_12_16_0  (
            .in0(N__9728),
            .in1(N__9699),
            .in2(N__9693),
            .in3(N__9680),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10752),
            .ce(),
            .sr(N__11149));
    defparam \U712_REG_SM.LDSn_LC_12_16_2 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_LC_12_16_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.LDSn_LC_12_16_2 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \U712_REG_SM.LDSn_LC_12_16_2  (
            .in0(N__9600),
            .in1(N__9654),
            .in2(N__9638),
            .in3(N__9533),
            .lcout(LDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10752),
            .ce(),
            .sr(N__11149));
    defparam \U712_REG_SM.UDSn_LC_12_16_7 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_LC_12_16_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.UDSn_LC_12_16_7 .LUT_INIT=16'b1010111110101100;
    LogicCell40 \U712_REG_SM.UDSn_LC_12_16_7  (
            .in0(N__9494),
            .in1(N__9601),
            .in2(N__9534),
            .in3(N__9909),
            .lcout(UDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10752),
            .ce(),
            .sr(N__11149));
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_4.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_4.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_19_4 (
            .in0(N__10999),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_i_i_LC_12_20_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_i_i_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_i_i_LC_12_20_7 .LUT_INIT=16'b0000101010110000;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_i_i_LC_12_20_7  (
            .in0(N__9775),
            .in1(N__9867),
            .in2(N__10397),
            .in3(N__10478),
            .lcout(N_166),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CASn_LC_13_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_13_6_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_13_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9456),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10719),
            .ce(),
            .sr(N__11191));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_9_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_9_0  (
            .in0(N__10305),
            .in1(N__11530),
            .in2(_gnd_net_),
            .in3(N__11673),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__11256),
            .sr(N__11170));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_10_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_10_3  (
            .in0(N__11669),
            .in1(N__11495),
            .in2(_gnd_net_),
            .in3(N__10304),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11284),
            .ce(N__11253),
            .sr(N__11162));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_10_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_10_4  (
            .in0(N__11500),
            .in1(N__11732),
            .in2(_gnd_net_),
            .in3(N__11767),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11284),
            .ce(N__11253),
            .sr(N__11162));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_10_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_10_5  (
            .in0(N__10206),
            .in1(N__11496),
            .in2(_gnd_net_),
            .in3(N__10241),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11284),
            .ce(N__11253),
            .sr(N__11162));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_10_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_10_6  (
            .in0(N__10242),
            .in1(_gnd_net_),
            .in2(N__11529),
            .in3(N__11766),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11284),
            .ce(N__11253),
            .sr(N__11162));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_3  (
            .in0(N__10202),
            .in1(N__11490),
            .in2(_gnd_net_),
            .in3(N__10296),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__11251),
            .sr(N__11158));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_11_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_11_6  (
            .in0(N__11778),
            .in1(_gnd_net_),
            .in2(N__11528),
            .in3(N__10240),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__11251),
            .sr(N__11158));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_13_15_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_13_15_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_13_15_1  (
            .in0(N__10509),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10420),
            .lcout(\U712_BYTE_ENABLE.N_298_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDSn_RNO_0_LC_13_16_7 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_13_16_7 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \U712_REG_SM.UDSn_RNO_0_LC_13_16_7  (
            .in0(N__10584),
            .in1(N__9854),
            .in2(N__10422),
            .in3(N__10508),
            .lcout(\U712_REG_SM.N_459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_390_i_LC_13_20_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_390_i_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_390_i_LC_13_20_0 .LUT_INIT=16'b0011110000101000;
    LogicCell40 \U712_BYTE_ENABLE.N_390_i_LC_13_20_0  (
            .in0(N__9793),
            .in1(N__10499),
            .in2(N__10416),
            .in3(N__9873),
            .lcout(N_390_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_389_i_LC_13_20_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_389_i_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_389_i_LC_13_20_2 .LUT_INIT=16'b0011110000010100;
    LogicCell40 \U712_BYTE_ENABLE.N_389_i_LC_13_20_2  (
            .in0(N__9792),
            .in1(N__10498),
            .in2(N__10415),
            .in3(N__9872),
            .lcout(N_389_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_13_20_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_13_20_5 .LUT_INIT=16'b0000011100110000;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_13_20_5  (
            .in0(N__9871),
            .in1(N__9791),
            .in2(N__10507),
            .in3(N__10398),
            .lcout(N_189),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_8_3  (
            .in0(N__11535),
            .in1(N__11610),
            .in2(_gnd_net_),
            .in3(N__11667),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11285),
            .ce(N__11259),
            .sr(N__11186));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_10_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_10_2  (
            .in0(N__10303),
            .in1(N__11494),
            .in2(_gnd_net_),
            .in3(N__10195),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11282),
            .ce(N__11257),
            .sr(N__11171));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_11_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_11_1  (
            .in0(N__10231),
            .in1(N__11470),
            .in2(_gnd_net_),
            .in3(N__10194),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__11252),
            .sr(N__11163));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_11_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_11_3  (
            .in0(N__10133),
            .in1(N__11471),
            .in2(_gnd_net_),
            .in3(N__11731),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__11252),
            .sr(N__11163));
    defparam \U712_CHIP_RAM.CRCSn_LC_15_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_15_6_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_15_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_15_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10091),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10724),
            .ce(),
            .sr(N__11196));
    defparam \U712_CHIP_RAM.WEn_LC_15_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_15_7_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_15_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_15_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10032),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10729),
            .ce(),
            .sr(N__11193));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_8_7  (
            .in0(N__11534),
            .in1(N__11622),
            .in2(_gnd_net_),
            .in3(N__11372),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__11261),
            .sr(N__11192));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_2  (
            .in0(N__11321),
            .in1(N__11533),
            .in2(_gnd_net_),
            .in3(N__11364),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__11260),
            .sr(N__11187));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_10_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_10_2  (
            .in0(N__11532),
            .in1(N__11618),
            .in2(_gnd_net_),
            .in3(N__11371),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11281),
            .ce(N__11258),
            .sr(N__11177));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_11_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_11_1  (
            .in0(N__11777),
            .in1(N__11446),
            .in2(_gnd_net_),
            .in3(N__11730),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__11254),
            .sr(N__11172));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_11_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_11_5  (
            .in0(N__11668),
            .in1(N__11445),
            .in2(_gnd_net_),
            .in3(N__11611),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__11254),
            .sr(N__11172));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_8_5  (
            .in0(N__11539),
            .in1(N__11373),
            .in2(_gnd_net_),
            .in3(N__11325),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11283),
            .ce(N__11262),
            .sr(N__11194));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_16_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_16_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_16_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_16_10_0  (
            .in0(N__10876),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11016),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10746),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_16_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_16_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_16_10_3 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_16_10_3  (
            .in0(N__11058),
            .in1(N__10875),
            .in2(_gnd_net_),
            .in3(N__11043),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10746),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_16_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_16_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_16_11_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_2_LC_16_11_2  (
            .in0(N__10834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10785),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10751),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_24_19_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_24_19_1 .LUT_INIT=16'b0011010101010101;
    LogicCell40 \U712_BUFFERS.DRDDIR_0_m2_LC_24_19_1  (
            .in0(N__10620),
            .in1(N__10583),
            .in2(N__11923),
            .in3(N__11835),
            .lcout(DRDDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

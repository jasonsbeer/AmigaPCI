-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Feb 8 2025 11:14:35

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U109_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U109_TOP
entity U109_TOP is
port (
    AD0 : out std_logic_vector(7 downto 0);
    AD2 : out std_logic_vector(7 downto 0);
    DLL : in std_logic_vector(7 downto 0);
    DUU : in std_logic_vector(7 downto 0);
    AD1 : out std_logic_vector(7 downto 0);
    AD3 : out std_logic_vector(7 downto 0);
    DLM : in std_logic_vector(7 downto 0);
    DUM : in std_logic_vector(7 downto 0);
    PCICYCLEn : out std_logic;
    ADLATCH : out std_logic;
    PCI_DIR : out std_logic;
    ALATCH : out std_logic);
end U109_TOP;

-- Architecture of U109_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U109_TOP is

signal \N__2211\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2200\ : std_logic;
signal \N__2193\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2184\ : std_logic;
signal \N__2183\ : std_logic;
signal \N__2182\ : std_logic;
signal \N__2175\ : std_logic;
signal \N__2174\ : std_logic;
signal \N__2173\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2165\ : std_logic;
signal \N__2164\ : std_logic;
signal \N__2157\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2155\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2147\ : std_logic;
signal \N__2146\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2138\ : std_logic;
signal \N__2137\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2129\ : std_logic;
signal \N__2128\ : std_logic;
signal \N__2121\ : std_logic;
signal \N__2120\ : std_logic;
signal \N__2119\ : std_logic;
signal \N__2112\ : std_logic;
signal \N__2111\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2103\ : std_logic;
signal \N__2102\ : std_logic;
signal \N__2101\ : std_logic;
signal \N__2094\ : std_logic;
signal \N__2093\ : std_logic;
signal \N__2092\ : std_logic;
signal \N__2085\ : std_logic;
signal \N__2084\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2076\ : std_logic;
signal \N__2075\ : std_logic;
signal \N__2074\ : std_logic;
signal \N__2067\ : std_logic;
signal \N__2066\ : std_logic;
signal \N__2065\ : std_logic;
signal \N__2058\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2056\ : std_logic;
signal \N__2049\ : std_logic;
signal \N__2048\ : std_logic;
signal \N__2047\ : std_logic;
signal \N__2040\ : std_logic;
signal \N__2039\ : std_logic;
signal \N__2038\ : std_logic;
signal \N__2031\ : std_logic;
signal \N__2030\ : std_logic;
signal \N__2029\ : std_logic;
signal \N__2022\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2020\ : std_logic;
signal \N__2013\ : std_logic;
signal \N__2012\ : std_logic;
signal \N__2011\ : std_logic;
signal \N__2004\ : std_logic;
signal \N__2003\ : std_logic;
signal \N__2002\ : std_logic;
signal \N__1995\ : std_logic;
signal \N__1994\ : std_logic;
signal \N__1993\ : std_logic;
signal \N__1986\ : std_logic;
signal \N__1985\ : std_logic;
signal \N__1984\ : std_logic;
signal \N__1977\ : std_logic;
signal \N__1976\ : std_logic;
signal \N__1975\ : std_logic;
signal \N__1968\ : std_logic;
signal \N__1967\ : std_logic;
signal \N__1966\ : std_logic;
signal \N__1959\ : std_logic;
signal \N__1958\ : std_logic;
signal \N__1957\ : std_logic;
signal \N__1950\ : std_logic;
signal \N__1949\ : std_logic;
signal \N__1948\ : std_logic;
signal \N__1941\ : std_logic;
signal \N__1940\ : std_logic;
signal \N__1939\ : std_logic;
signal \N__1932\ : std_logic;
signal \N__1931\ : std_logic;
signal \N__1930\ : std_logic;
signal \N__1923\ : std_logic;
signal \N__1922\ : std_logic;
signal \N__1921\ : std_logic;
signal \N__1914\ : std_logic;
signal \N__1913\ : std_logic;
signal \N__1912\ : std_logic;
signal \N__1905\ : std_logic;
signal \N__1904\ : std_logic;
signal \N__1903\ : std_logic;
signal \N__1896\ : std_logic;
signal \N__1895\ : std_logic;
signal \N__1894\ : std_logic;
signal \N__1887\ : std_logic;
signal \N__1886\ : std_logic;
signal \N__1885\ : std_logic;
signal \N__1878\ : std_logic;
signal \N__1877\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1869\ : std_logic;
signal \N__1868\ : std_logic;
signal \N__1867\ : std_logic;
signal \N__1860\ : std_logic;
signal \N__1859\ : std_logic;
signal \N__1858\ : std_logic;
signal \N__1851\ : std_logic;
signal \N__1850\ : std_logic;
signal \N__1849\ : std_logic;
signal \N__1842\ : std_logic;
signal \N__1841\ : std_logic;
signal \N__1840\ : std_logic;
signal \N__1833\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1831\ : std_logic;
signal \N__1824\ : std_logic;
signal \N__1823\ : std_logic;
signal \N__1822\ : std_logic;
signal \N__1815\ : std_logic;
signal \N__1814\ : std_logic;
signal \N__1813\ : std_logic;
signal \N__1806\ : std_logic;
signal \N__1805\ : std_logic;
signal \N__1804\ : std_logic;
signal \N__1797\ : std_logic;
signal \N__1796\ : std_logic;
signal \N__1795\ : std_logic;
signal \N__1788\ : std_logic;
signal \N__1787\ : std_logic;
signal \N__1786\ : std_logic;
signal \N__1779\ : std_logic;
signal \N__1778\ : std_logic;
signal \N__1777\ : std_logic;
signal \N__1770\ : std_logic;
signal \N__1769\ : std_logic;
signal \N__1768\ : std_logic;
signal \N__1761\ : std_logic;
signal \N__1760\ : std_logic;
signal \N__1759\ : std_logic;
signal \N__1752\ : std_logic;
signal \N__1751\ : std_logic;
signal \N__1750\ : std_logic;
signal \N__1743\ : std_logic;
signal \N__1742\ : std_logic;
signal \N__1741\ : std_logic;
signal \N__1734\ : std_logic;
signal \N__1733\ : std_logic;
signal \N__1732\ : std_logic;
signal \N__1725\ : std_logic;
signal \N__1724\ : std_logic;
signal \N__1723\ : std_logic;
signal \N__1716\ : std_logic;
signal \N__1715\ : std_logic;
signal \N__1714\ : std_logic;
signal \N__1707\ : std_logic;
signal \N__1706\ : std_logic;
signal \N__1705\ : std_logic;
signal \N__1698\ : std_logic;
signal \N__1697\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1689\ : std_logic;
signal \N__1688\ : std_logic;
signal \N__1687\ : std_logic;
signal \N__1680\ : std_logic;
signal \N__1679\ : std_logic;
signal \N__1678\ : std_logic;
signal \N__1671\ : std_logic;
signal \N__1670\ : std_logic;
signal \N__1669\ : std_logic;
signal \N__1662\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1660\ : std_logic;
signal \N__1653\ : std_logic;
signal \N__1652\ : std_logic;
signal \N__1651\ : std_logic;
signal \N__1644\ : std_logic;
signal \N__1643\ : std_logic;
signal \N__1642\ : std_logic;
signal \N__1635\ : std_logic;
signal \N__1634\ : std_logic;
signal \N__1633\ : std_logic;
signal \N__1626\ : std_logic;
signal \N__1625\ : std_logic;
signal \N__1624\ : std_logic;
signal \N__1617\ : std_logic;
signal \N__1616\ : std_logic;
signal \N__1615\ : std_logic;
signal \N__1608\ : std_logic;
signal \N__1607\ : std_logic;
signal \N__1606\ : std_logic;
signal \N__1589\ : std_logic;
signal \N__1586\ : std_logic;
signal \N__1583\ : std_logic;
signal \N__1580\ : std_logic;
signal \N__1577\ : std_logic;
signal \N__1574\ : std_logic;
signal \N__1571\ : std_logic;
signal \N__1568\ : std_logic;
signal \N__1565\ : std_logic;
signal \N__1562\ : std_logic;
signal \N__1559\ : std_logic;
signal \N__1556\ : std_logic;
signal \N__1553\ : std_logic;
signal \N__1550\ : std_logic;
signal \N__1547\ : std_logic;
signal \N__1544\ : std_logic;
signal \N__1541\ : std_logic;
signal \N__1538\ : std_logic;
signal \N__1535\ : std_logic;
signal \N__1532\ : std_logic;
signal \N__1529\ : std_logic;
signal \N__1526\ : std_logic;
signal \N__1523\ : std_logic;
signal \N__1520\ : std_logic;
signal \N__1517\ : std_logic;
signal \N__1514\ : std_logic;
signal \N__1511\ : std_logic;
signal \N__1508\ : std_logic;
signal \N__1505\ : std_logic;
signal \N__1502\ : std_logic;
signal \N__1499\ : std_logic;
signal \N__1496\ : std_logic;
signal \N__1493\ : std_logic;
signal \N__1490\ : std_logic;
signal \N__1487\ : std_logic;
signal \N__1484\ : std_logic;
signal \N__1481\ : std_logic;
signal \N__1478\ : std_logic;
signal \N__1475\ : std_logic;
signal \N__1472\ : std_logic;
signal \N__1469\ : std_logic;
signal \N__1466\ : std_logic;
signal \N__1463\ : std_logic;
signal \N__1460\ : std_logic;
signal \N__1457\ : std_logic;
signal \N__1454\ : std_logic;
signal \N__1451\ : std_logic;
signal \N__1448\ : std_logic;
signal \N__1445\ : std_logic;
signal \N__1442\ : std_logic;
signal \N__1439\ : std_logic;
signal \N__1436\ : std_logic;
signal \N__1433\ : std_logic;
signal \N__1430\ : std_logic;
signal \N__1427\ : std_logic;
signal \N__1424\ : std_logic;
signal \N__1421\ : std_logic;
signal \N__1418\ : std_logic;
signal \N__1415\ : std_logic;
signal \N__1412\ : std_logic;
signal \N__1409\ : std_logic;
signal \N__1406\ : std_logic;
signal \N__1403\ : std_logic;
signal \N__1400\ : std_logic;
signal \N__1397\ : std_logic;
signal \N__1394\ : std_logic;
signal \N__1391\ : std_logic;
signal \N__1388\ : std_logic;
signal \N__1385\ : std_logic;
signal \N__1382\ : std_logic;
signal \N__1379\ : std_logic;
signal \N__1376\ : std_logic;
signal \N__1373\ : std_logic;
signal \N__1370\ : std_logic;
signal \N__1367\ : std_logic;
signal \N__1364\ : std_logic;
signal \N__1361\ : std_logic;
signal \N__1358\ : std_logic;
signal \N__1355\ : std_logic;
signal \N__1352\ : std_logic;
signal \N__1349\ : std_logic;
signal \N__1346\ : std_logic;
signal \N__1343\ : std_logic;
signal \N__1340\ : std_logic;
signal \N__1337\ : std_logic;
signal \N__1334\ : std_logic;
signal \N__1331\ : std_logic;
signal \N__1328\ : std_logic;
signal \N__1325\ : std_logic;
signal \N__1322\ : std_logic;
signal \N__1319\ : std_logic;
signal \N__1316\ : std_logic;
signal \N__1313\ : std_logic;
signal \N__1310\ : std_logic;
signal \N__1307\ : std_logic;
signal \N__1304\ : std_logic;
signal \N__1301\ : std_logic;
signal \N__1298\ : std_logic;
signal \N__1295\ : std_logic;
signal \N__1292\ : std_logic;
signal \N__1289\ : std_logic;
signal \N__1286\ : std_logic;
signal \N__1283\ : std_logic;
signal \N__1280\ : std_logic;
signal \N__1277\ : std_logic;
signal \N__1274\ : std_logic;
signal \N__1271\ : std_logic;
signal \N__1268\ : std_logic;
signal \N__1265\ : std_logic;
signal \N__1262\ : std_logic;
signal \N__1259\ : std_logic;
signal \N__1256\ : std_logic;
signal \N__1253\ : std_logic;
signal \N__1250\ : std_logic;
signal \N__1247\ : std_logic;
signal \N__1244\ : std_logic;
signal \N__1241\ : std_logic;
signal \N__1238\ : std_logic;
signal \N__1235\ : std_logic;
signal \N__1232\ : std_logic;
signal \N__1229\ : std_logic;
signal \N__1226\ : std_logic;
signal \N__1223\ : std_logic;
signal \N__1220\ : std_logic;
signal \N__1217\ : std_logic;
signal \N__1214\ : std_logic;
signal \N__1211\ : std_logic;
signal \N__1208\ : std_logic;
signal \N__1205\ : std_logic;
signal \N__1202\ : std_logic;
signal \N__1199\ : std_logic;
signal \N__1196\ : std_logic;
signal \N__1193\ : std_logic;
signal \N__1190\ : std_logic;
signal \N__1187\ : std_logic;
signal \N__1184\ : std_logic;
signal \N__1181\ : std_logic;
signal \N__1178\ : std_logic;
signal \N__1175\ : std_logic;
signal \N__1172\ : std_logic;
signal \N__1169\ : std_logic;
signal \N__1166\ : std_logic;
signal \N__1163\ : std_logic;
signal \N__1160\ : std_logic;
signal \N__1157\ : std_logic;
signal \N__1154\ : std_logic;
signal \N__1151\ : std_logic;
signal \N__1148\ : std_logic;
signal \N__1145\ : std_logic;
signal \N__1142\ : std_logic;
signal \N__1139\ : std_logic;
signal \N__1136\ : std_logic;
signal \N__1133\ : std_logic;
signal \N__1130\ : std_logic;
signal \N__1127\ : std_logic;
signal \N__1124\ : std_logic;
signal \N__1121\ : std_logic;
signal \N__1118\ : std_logic;
signal \N__1115\ : std_logic;
signal \N__1112\ : std_logic;
signal \N__1109\ : std_logic;
signal \N__1106\ : std_logic;
signal \N__1103\ : std_logic;
signal \N__1100\ : std_logic;
signal \N__1097\ : std_logic;
signal \N__1094\ : std_logic;
signal \N__1091\ : std_logic;
signal \N__1088\ : std_logic;
signal \N__1085\ : std_logic;
signal \N__1082\ : std_logic;
signal \N__1079\ : std_logic;
signal \N__1076\ : std_logic;
signal \N__1073\ : std_logic;
signal \N__1070\ : std_logic;
signal \N__1067\ : std_logic;
signal \N__1064\ : std_logic;
signal \N__1061\ : std_logic;
signal \N__1058\ : std_logic;
signal \N__1055\ : std_logic;
signal \N__1052\ : std_logic;
signal \N__1049\ : std_logic;
signal \N__1046\ : std_logic;
signal \N__1043\ : std_logic;
signal \N__1040\ : std_logic;
signal \N__1037\ : std_logic;
signal \N__1034\ : std_logic;
signal \N__1031\ : std_logic;
signal \N__1028\ : std_logic;
signal \N__1025\ : std_logic;
signal \N__1022\ : std_logic;
signal \N__1019\ : std_logic;
signal \N__1016\ : std_logic;
signal \N__1013\ : std_logic;
signal \N__1010\ : std_logic;
signal \N__1007\ : std_logic;
signal \N__1004\ : std_logic;
signal \N__1001\ : std_logic;
signal \N__998\ : std_logic;
signal \N__995\ : std_logic;
signal \N__992\ : std_logic;
signal \N__989\ : std_logic;
signal \N__986\ : std_logic;
signal \N__983\ : std_logic;
signal \N__980\ : std_logic;
signal \N__977\ : std_logic;
signal \N__974\ : std_logic;
signal \N__971\ : std_logic;
signal \N__968\ : std_logic;
signal \N__965\ : std_logic;
signal \N__962\ : std_logic;
signal \N__959\ : std_logic;
signal \N__956\ : std_logic;
signal \N__953\ : std_logic;
signal \N__950\ : std_logic;
signal \N__947\ : std_logic;
signal \N__944\ : std_logic;
signal \N__941\ : std_logic;
signal \N__938\ : std_logic;
signal \N__935\ : std_logic;
signal \N__932\ : std_logic;
signal \N__929\ : std_logic;
signal \N__926\ : std_logic;
signal \N__923\ : std_logic;
signal \N__920\ : std_logic;
signal \N__917\ : std_logic;
signal \N__914\ : std_logic;
signal \N__911\ : std_logic;
signal \N__908\ : std_logic;
signal \N__905\ : std_logic;
signal \N__902\ : std_logic;
signal \N__899\ : std_logic;
signal \N__896\ : std_logic;
signal \N__893\ : std_logic;
signal \N__890\ : std_logic;
signal \N__887\ : std_logic;
signal \N__884\ : std_logic;
signal \N__881\ : std_logic;
signal \N__878\ : std_logic;
signal \N__875\ : std_logic;
signal \N__872\ : std_logic;
signal \N__869\ : std_logic;
signal \N__866\ : std_logic;
signal \N__863\ : std_logic;
signal \N__860\ : std_logic;
signal \N__857\ : std_logic;
signal \N__854\ : std_logic;
signal \N__851\ : std_logic;
signal \N__848\ : std_logic;
signal \N__845\ : std_logic;
signal \N__842\ : std_logic;
signal \N__839\ : std_logic;
signal \N__836\ : std_logic;
signal \N__833\ : std_logic;
signal \N__830\ : std_logic;
signal \N__827\ : std_logic;
signal \N__824\ : std_logic;
signal \N__821\ : std_logic;
signal \N__818\ : std_logic;
signal \N__815\ : std_logic;
signal \N__812\ : std_logic;
signal \N__809\ : std_logic;
signal \N__806\ : std_logic;
signal \N__803\ : std_logic;
signal \N__800\ : std_logic;
signal \AD0_c_2\ : std_logic;
signal \AD3_c_0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \AD1_c_6\ : std_logic;
signal \AD3_c_6\ : std_logic;
signal \AD2_c_3\ : std_logic;
signal \AD0_c_3\ : std_logic;
signal \AD1_c_0\ : std_logic;
signal \AD3_c_4\ : std_logic;
signal \AD2_c_4\ : std_logic;
signal \AD2_c_5\ : std_logic;
signal \AD3_c_3\ : std_logic;
signal \AD0_c_1\ : std_logic;
signal \GNDG0\ : std_logic;
signal \AD1_c_2\ : std_logic;
signal \AD2_c_6\ : std_logic;
signal \AD0_c_4\ : std_logic;
signal \AD1_c_5\ : std_logic;
signal \AD2_c_7\ : std_logic;
signal \AD3_c_1\ : std_logic;
signal \AD1_c_3\ : std_logic;
signal \AD0_c_7\ : std_logic;
signal \AD2_c_0\ : std_logic;
signal \AD3_c_5\ : std_logic;
signal \AD0_c_6\ : std_logic;
signal \AD1_c_7\ : std_logic;
signal \AD3_c_7\ : std_logic;
signal \AD2_c_1\ : std_logic;
signal \AD0_c_5\ : std_logic;
signal \AD2_c_2\ : std_logic;
signal \AD1_c_4\ : std_logic;
signal \AD0_c_0\ : std_logic;
signal \AD1_c_1\ : std_logic;
signal \AD3_c_2\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \AD3_wire\ : std_logic_vector(7 downto 0);
signal \DUM_wire\ : std_logic_vector(7 downto 0);
signal \DUU_wire\ : std_logic_vector(7 downto 0);
signal \AD1_wire\ : std_logic_vector(7 downto 0);
signal \DLM_wire\ : std_logic_vector(7 downto 0);
signal \AD0_wire\ : std_logic_vector(7 downto 0);
signal \AD2_wire\ : std_logic_vector(7 downto 0);
signal \DLL_wire\ : std_logic_vector(7 downto 0);
signal \PCI_DIR_wire\ : std_logic;
signal \ADLATCH_wire\ : std_logic;
signal \ALATCH_wire\ : std_logic;
signal \PCICYCLEn_wire\ : std_logic;

begin
    AD3 <= \AD3_wire\;
    \DUM_wire\ <= DUM;
    \DUU_wire\ <= DUU;
    AD1 <= \AD1_wire\;
    \DLM_wire\ <= DLM;
    AD0 <= \AD0_wire\;
    AD2 <= \AD2_wire\;
    \DLL_wire\ <= DLL;
    PCI_DIR <= \PCI_DIR_wire\;
    ADLATCH <= \ADLATCH_wire\;
    ALATCH <= \ALATCH_wire\;
    PCICYCLEn <= \PCICYCLEn_wire\;

    \AD3_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2211\,
            DIN => \N__2210\,
            DOUT => \N__2209\,
            PACKAGEPIN => \AD3_wire\(2)
        );

    \AD3_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2211\,
            PADOUT => \N__2210\,
            PADIN => \N__2209\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1562\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUM_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2202\,
            DIN => \N__2201\,
            DOUT => \N__2200\,
            PACKAGEPIN => \DUM_wire\(1)
        );

    \DUM_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2202\,
            PADOUT => \N__2201\,
            PADIN => \N__2200\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD1_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUU_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2193\,
            DIN => \N__2192\,
            DOUT => \N__2191\,
            PACKAGEPIN => \DUU_wire\(0)
        );

    \DUU_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2193\,
            PADOUT => \N__2192\,
            PADIN => \N__2191\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD0_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD1_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2184\,
            DIN => \N__2183\,
            DOUT => \N__2182\,
            PACKAGEPIN => \AD1_wire\(4)
        );

    \AD1_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2184\,
            PADOUT => \N__2183\,
            PADIN => \N__2182\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1313\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLM_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2175\,
            DIN => \N__2174\,
            DOUT => \N__2173\,
            PACKAGEPIN => \DLM_wire\(2)
        );

    \DLM_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2175\,
            PADOUT => \N__2174\,
            PADIN => \N__2173\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD2_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD0_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2166\,
            DIN => \N__2165\,
            DOUT => \N__2164\,
            PACKAGEPIN => \AD0_wire\(5)
        );

    \AD0_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2166\,
            PADOUT => \N__2165\,
            PADIN => \N__2164\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1364\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD2_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2157\,
            DIN => \N__2156\,
            DOUT => \N__2155\,
            PACKAGEPIN => \AD2_wire\(1)
        );

    \AD2_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2157\,
            PADOUT => \N__2156\,
            PADIN => \N__2155\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1391\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLL_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2148\,
            DIN => \N__2147\,
            DOUT => \N__2146\,
            PACKAGEPIN => \DLL_wire\(7)
        );

    \DLL_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2148\,
            PADOUT => \N__2147\,
            PADIN => \N__2146\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD3_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUM_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2139\,
            DIN => \N__2138\,
            DOUT => \N__2137\,
            PACKAGEPIN => \DUM_wire\(7)
        );

    \DUM_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2139\,
            PADOUT => \N__2138\,
            PADIN => \N__2137\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD1_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUU_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2130\,
            DIN => \N__2129\,
            DOUT => \N__2128\,
            PACKAGEPIN => \DUU_wire\(6)
        );

    \DUU_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2130\,
            PADOUT => \N__2129\,
            PADIN => \N__2128\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD0_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD3_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2121\,
            DIN => \N__2120\,
            DOUT => \N__2119\,
            PACKAGEPIN => \AD3_wire\(5)
        );

    \AD3_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2121\,
            PADOUT => \N__2120\,
            PADIN => \N__2119\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1478\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLM_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2112\,
            DIN => \N__2111\,
            DOUT => \N__2110\,
            PACKAGEPIN => \DLM_wire\(0)
        );

    \DLM_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2112\,
            PADOUT => \N__2111\,
            PADIN => \N__2110\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD2_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD0_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2103\,
            DIN => \N__2102\,
            DOUT => \N__2101\,
            PACKAGEPIN => \AD0_wire\(7)
        );

    \AD0_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2103\,
            PADOUT => \N__2102\,
            PADIN => \N__2101\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1526\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD1_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2094\,
            DIN => \N__2093\,
            DOUT => \N__2092\,
            PACKAGEPIN => \AD1_wire\(3)
        );

    \AD1_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2094\,
            PADOUT => \N__2093\,
            PADIN => \N__2092\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1121\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLL_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2085\,
            DIN => \N__2084\,
            DOUT => \N__2083\,
            PACKAGEPIN => \DLL_wire\(1)
        );

    \DLL_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2085\,
            PADOUT => \N__2084\,
            PADIN => \N__2083\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD3_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLM_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2076\,
            DIN => \N__2075\,
            DOUT => \N__2074\,
            PACKAGEPIN => \DLM_wire\(7)
        );

    \DLM_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2076\,
            PADOUT => \N__2075\,
            PADIN => \N__2074\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD2_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUM_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2067\,
            DIN => \N__2066\,
            DOUT => \N__2065\,
            PACKAGEPIN => \DUM_wire\(5)
        );

    \DUM_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2067\,
            PADOUT => \N__2066\,
            PADIN => \N__2065\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD1_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUU_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2058\,
            DIN => \N__2057\,
            DOUT => \N__2056\,
            PACKAGEPIN => \DUU_wire\(4)
        );

    \DUU_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2058\,
            PADOUT => \N__2057\,
            PADIN => \N__2056\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD0_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD2_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2049\,
            DIN => \N__2048\,
            DOUT => \N__2047\,
            PACKAGEPIN => \AD2_wire\(6)
        );

    \AD2_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2049\,
            PADOUT => \N__2048\,
            PADIN => \N__2047\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1238\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD3_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2040\,
            DIN => \N__2039\,
            DOUT => \N__2038\,
            PACKAGEPIN => \AD3_wire\(7)
        );

    \AD3_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2040\,
            PADOUT => \N__2039\,
            PADIN => \N__2038\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1412\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUM_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2031\,
            DIN => \N__2030\,
            DOUT => \N__2029\,
            PACKAGEPIN => \DUM_wire\(2)
        );

    \DUM_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2031\,
            PADOUT => \N__2030\,
            PADIN => \N__2029\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD1_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PCI_DIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2022\,
            DIN => \N__2021\,
            DOUT => \N__2020\,
            PACKAGEPIN => \PCI_DIR_wire\
        );

    \PCI_DIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2022\,
            PADOUT => \N__2021\,
            PADIN => \N__2020\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD0_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2013\,
            DIN => \N__2012\,
            DOUT => \N__2011\,
            PACKAGEPIN => \AD0_wire\(1)
        );

    \AD0_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2013\,
            PADOUT => \N__2012\,
            PADIN => \N__2011\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__941\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD1_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2004\,
            DIN => \N__2003\,
            DOUT => \N__2002\,
            PACKAGEPIN => \AD1_wire\(1)
        );

    \AD1_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2004\,
            PADOUT => \N__2003\,
            PADIN => \N__2002\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1589\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLL_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1995\,
            DIN => \N__1994\,
            DOUT => \N__1993\,
            PACKAGEPIN => \DLL_wire\(3)
        );

    \DLL_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1995\,
            PADOUT => \N__1994\,
            PADIN => \N__1993\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD3_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLM_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1986\,
            DIN => \N__1985\,
            DOUT => \N__1984\,
            PACKAGEPIN => \DLM_wire\(5)
        );

    \DLM_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1986\,
            PADOUT => \N__1985\,
            PADIN => \N__1984\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD2_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD2_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1977\,
            DIN => \N__1976\,
            DOUT => \N__1975\,
            PACKAGEPIN => \AD2_wire\(4)
        );

    \AD2_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1977\,
            PADOUT => \N__1976\,
            PADIN => \N__1975\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1019\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD3_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1968\,
            DIN => \N__1967\,
            DOUT => \N__1966\,
            PACKAGEPIN => \AD3_wire\(1)
        );

    \AD3_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1968\,
            PADOUT => \N__1967\,
            PADIN => \N__1966\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1145\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLL_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1959\,
            DIN => \N__1958\,
            DOUT => \N__1957\,
            PACKAGEPIN => \DLL_wire\(4)
        );

    \DLL_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1959\,
            PADOUT => \N__1958\,
            PADIN => \N__1957\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD3_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUM_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1950\,
            DIN => \N__1949\,
            DOUT => \N__1948\,
            PACKAGEPIN => \DUM_wire\(0)
        );

    \DUM_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1950\,
            PADOUT => \N__1949\,
            PADIN => \N__1948\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD1_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUU_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1941\,
            DIN => \N__1940\,
            DOUT => \N__1939\,
            PACKAGEPIN => \DUU_wire\(3)
        );

    \DUU_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1941\,
            PADOUT => \N__1940\,
            PADIN => \N__1939\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD0_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD0_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1932\,
            DIN => \N__1931\,
            DOUT => \N__1930\,
            PACKAGEPIN => \AD0_wire\(3)
        );

    \AD0_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1932\,
            PADOUT => \N__1931\,
            PADIN => \N__1930\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1094\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD1_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1923\,
            DIN => \N__1922\,
            DOUT => \N__1921\,
            PACKAGEPIN => \AD1_wire\(7)
        );

    \AD1_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1923\,
            PADOUT => \N__1922\,
            PADIN => \N__1921\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1427\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLM_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1914\,
            DIN => \N__1913\,
            DOUT => \N__1912\,
            PACKAGEPIN => \DLM_wire\(3)
        );

    \DLM_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1914\,
            PADOUT => \N__1913\,
            PADIN => \N__1912\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD2_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD2_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1905\,
            DIN => \N__1904\,
            DOUT => \N__1903\,
            PACKAGEPIN => \AD2_wire\(2)
        );

    \AD2_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1905\,
            PADOUT => \N__1904\,
            PADIN => \N__1903\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1340\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD3_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1896\,
            DIN => \N__1895\,
            DOUT => \N__1894\,
            PACKAGEPIN => \AD3_wire\(3)
        );

    \AD3_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1896\,
            PADOUT => \N__1895\,
            PADIN => \N__1894\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__968\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLL_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1887\,
            DIN => \N__1886\,
            DOUT => \N__1885\,
            PACKAGEPIN => \DLL_wire\(6)
        );

    \DLL_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1887\,
            PADOUT => \N__1886\,
            PADIN => \N__1885\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD3_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUM_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1878\,
            DIN => \N__1877\,
            DOUT => \N__1876\,
            PACKAGEPIN => \DUM_wire\(6)
        );

    \DUM_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1878\,
            PADOUT => \N__1877\,
            PADIN => \N__1876\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD1_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUU_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1869\,
            DIN => \N__1868\,
            DOUT => \N__1867\,
            PACKAGEPIN => \DUU_wire\(1)
        );

    \DUU_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1869\,
            PADOUT => \N__1868\,
            PADIN => \N__1867\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD0_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD1_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1860\,
            DIN => \N__1859\,
            DOUT => \N__1858\,
            PACKAGEPIN => \AD1_wire\(5)
        );

    \AD1_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1860\,
            PADOUT => \N__1859\,
            PADIN => \N__1858\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1190\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD3_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1851\,
            DIN => \N__1850\,
            DOUT => \N__1849\,
            PACKAGEPIN => \AD3_wire\(4)
        );

    \AD3_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1851\,
            PADOUT => \N__1850\,
            PADIN => \N__1849\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1049\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADLATCH_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1842\,
            DIN => \N__1841\,
            DOUT => \N__1840\,
            PACKAGEPIN => \ADLATCH_wire\
        );

    \ADLATCH_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1842\,
            PADOUT => \N__1841\,
            PADIN => \N__1840\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLM_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1833\,
            DIN => \N__1832\,
            DOUT => \N__1831\,
            PACKAGEPIN => \DLM_wire\(1)
        );

    \DLM_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1833\,
            PADOUT => \N__1832\,
            PADIN => \N__1831\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD2_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD0_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1824\,
            DIN => \N__1823\,
            DOUT => \N__1822\,
            PACKAGEPIN => \AD0_wire\(4)
        );

    \AD0_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1824\,
            PADOUT => \N__1823\,
            PADIN => \N__1822\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1214\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD1_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1815\,
            DIN => \N__1814\,
            DOUT => \N__1813\,
            PACKAGEPIN => \AD1_wire\(2)
        );

    \AD1_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1815\,
            PADOUT => \N__1814\,
            PADIN => \N__1813\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1265\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD2_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1806\,
            DIN => \N__1805\,
            DOUT => \N__1804\,
            PACKAGEPIN => \AD2_wire\(0)
        );

    \AD2_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1806\,
            PADOUT => \N__1805\,
            PADIN => \N__1804\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1499\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ALATCH_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1797\,
            DIN => \N__1796\,
            DOUT => \N__1795\,
            PACKAGEPIN => \ALATCH_wire\
        );

    \ALATCH_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1797\,
            PADOUT => \N__1796\,
            PADIN => \N__1795\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLL_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1788\,
            DIN => \N__1787\,
            DOUT => \N__1786\,
            PACKAGEPIN => \DLL_wire\(0)
        );

    \DLL_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1788\,
            PADOUT => \N__1787\,
            PADIN => \N__1786\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD3_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUM_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1779\,
            DIN => \N__1778\,
            DOUT => \N__1777\,
            PACKAGEPIN => \DUM_wire\(4)
        );

    \DUM_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1779\,
            PADOUT => \N__1778\,
            PADIN => \N__1777\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD1_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUU_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1770\,
            DIN => \N__1769\,
            DOUT => \N__1768\,
            PACKAGEPIN => \DUU_wire\(7)
        );

    \DUU_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1770\,
            PADOUT => \N__1769\,
            PADIN => \N__1768\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD0_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD2_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1761\,
            DIN => \N__1760\,
            DOUT => \N__1759\,
            PACKAGEPIN => \AD2_wire\(7)
        );

    \AD2_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1761\,
            PADOUT => \N__1760\,
            PADIN => \N__1759\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1169\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD3_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1752\,
            DIN => \N__1751\,
            DOUT => \N__1750\,
            PACKAGEPIN => \AD3_wire\(6)
        );

    \AD3_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1752\,
            PADOUT => \N__1751\,
            PADIN => \N__1750\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__893\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD0_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1743\,
            DIN => \N__1742\,
            DOUT => \N__1741\,
            PACKAGEPIN => \AD0_wire\(6)
        );

    \AD0_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1743\,
            PADOUT => \N__1742\,
            PADIN => \N__1741\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1448\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD1_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1734\,
            DIN => \N__1733\,
            DOUT => \N__1732\,
            PACKAGEPIN => \AD1_wire\(0)
        );

    \AD1_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1734\,
            PADOUT => \N__1733\,
            PADIN => \N__1732\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1076\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLL_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1725\,
            DIN => \N__1724\,
            DOUT => \N__1723\,
            PACKAGEPIN => \DLL_wire\(2)
        );

    \DLL_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1725\,
            PADOUT => \N__1724\,
            PADIN => \N__1723\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD3_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLM_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1716\,
            DIN => \N__1715\,
            DOUT => \N__1714\,
            PACKAGEPIN => \DLM_wire\(6)
        );

    \DLM_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1716\,
            PADOUT => \N__1715\,
            PADIN => \N__1714\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD2_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUU_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1707\,
            DIN => \N__1706\,
            DOUT => \N__1705\,
            PACKAGEPIN => \DUU_wire\(5)
        );

    \DUU_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1707\,
            PADOUT => \N__1706\,
            PADIN => \N__1705\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD0_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD2_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1698\,
            DIN => \N__1697\,
            DOUT => \N__1696\,
            PACKAGEPIN => \AD2_wire\(5)
        );

    \AD2_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1698\,
            PADOUT => \N__1697\,
            PADIN => \N__1696\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__995\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD3_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1689\,
            DIN => \N__1688\,
            DOUT => \N__1687\,
            PACKAGEPIN => \AD3_wire\(0)
        );

    \AD3_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1689\,
            PADOUT => \N__1688\,
            PADIN => \N__1687\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__845\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUM_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1680\,
            DIN => \N__1679\,
            DOUT => \N__1678\,
            PACKAGEPIN => \DUM_wire\(3)
        );

    \DUM_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1680\,
            PADOUT => \N__1679\,
            PADIN => \N__1678\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD1_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DUU_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1671\,
            DIN => \N__1670\,
            DOUT => \N__1669\,
            PACKAGEPIN => \DUU_wire\(2)
        );

    \DUU_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1671\,
            PADOUT => \N__1670\,
            PADIN => \N__1669\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD0_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PCICYCLEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1662\,
            DIN => \N__1661\,
            DOUT => \N__1660\,
            PACKAGEPIN => \PCICYCLEn_wire\
        );

    \PCICYCLEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1662\,
            PADOUT => \N__1661\,
            PADIN => \N__1660\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1538\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD0_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1653\,
            DIN => \N__1652\,
            DOUT => \N__1651\,
            PACKAGEPIN => \AD0_wire\(0)
        );

    \AD0_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1653\,
            PADOUT => \N__1652\,
            PADIN => \N__1651\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1292\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD1_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1644\,
            DIN => \N__1643\,
            DOUT => \N__1642\,
            PACKAGEPIN => \AD1_wire\(6)
        );

    \AD1_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1644\,
            PADOUT => \N__1643\,
            PADIN => \N__1642\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__914\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLM_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1635\,
            DIN => \N__1634\,
            DOUT => \N__1633\,
            PACKAGEPIN => \DLM_wire\(4)
        );

    \DLM_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1635\,
            PADOUT => \N__1634\,
            PADIN => \N__1633\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD2_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD2_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1626\,
            DIN => \N__1625\,
            DOUT => \N__1624\,
            PACKAGEPIN => \AD2_wire\(3)
        );

    \AD2_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1626\,
            PADOUT => \N__1625\,
            PADIN => \N__1624\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__863\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DLL_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1617\,
            DIN => \N__1616\,
            DOUT => \N__1615\,
            PACKAGEPIN => \DLL_wire\(5)
        );

    \DLL_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1617\,
            PADOUT => \N__1616\,
            PADIN => \N__1615\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AD3_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AD0_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1608\,
            DIN => \N__1607\,
            DOUT => \N__1606\,
            PACKAGEPIN => \AD0_wire\(2)
        );

    \AD0_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1608\,
            PADOUT => \N__1607\,
            PADIN => \N__1606\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__821\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__335\ : IoInMux
    port map (
            O => \N__1589\,
            I => \N__1586\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__1586\,
            I => \N__1583\
        );

    \I__333\ : Span4Mux_s1_v
    port map (
            O => \N__1583\,
            I => \N__1580\
        );

    \I__332\ : Span4Mux_v
    port map (
            O => \N__1580\,
            I => \N__1577\
        );

    \I__331\ : Sp12to4
    port map (
            O => \N__1577\,
            I => \N__1574\
        );

    \I__330\ : Span12Mux_h
    port map (
            O => \N__1574\,
            I => \N__1571\
        );

    \I__329\ : Span12Mux_v
    port map (
            O => \N__1571\,
            I => \N__1568\
        );

    \I__328\ : Span12Mux_h
    port map (
            O => \N__1568\,
            I => \N__1565\
        );

    \I__327\ : Odrv12
    port map (
            O => \N__1565\,
            I => \AD1_c_1\
        );

    \I__326\ : IoInMux
    port map (
            O => \N__1562\,
            I => \N__1559\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__1559\,
            I => \N__1556\
        );

    \I__324\ : IoSpan4Mux
    port map (
            O => \N__1556\,
            I => \N__1553\
        );

    \I__323\ : Span4Mux_s3_h
    port map (
            O => \N__1553\,
            I => \N__1550\
        );

    \I__322\ : Sp12to4
    port map (
            O => \N__1550\,
            I => \N__1547\
        );

    \I__321\ : Span12Mux_v
    port map (
            O => \N__1547\,
            I => \N__1544\
        );

    \I__320\ : Span12Mux_v
    port map (
            O => \N__1544\,
            I => \N__1541\
        );

    \I__319\ : Odrv12
    port map (
            O => \N__1541\,
            I => \AD3_c_2\
        );

    \I__318\ : IoInMux
    port map (
            O => \N__1538\,
            I => \N__1535\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__1535\,
            I => \N__1532\
        );

    \I__316\ : Span4Mux_s3_h
    port map (
            O => \N__1532\,
            I => \N__1529\
        );

    \I__315\ : Odrv4
    port map (
            O => \N__1529\,
            I => \CONSTANT_ONE_NET\
        );

    \I__314\ : IoInMux
    port map (
            O => \N__1526\,
            I => \N__1523\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__1523\,
            I => \N__1520\
        );

    \I__312\ : IoSpan4Mux
    port map (
            O => \N__1520\,
            I => \N__1517\
        );

    \I__311\ : Span4Mux_s2_v
    port map (
            O => \N__1517\,
            I => \N__1514\
        );

    \I__310\ : Span4Mux_v
    port map (
            O => \N__1514\,
            I => \N__1511\
        );

    \I__309\ : Sp12to4
    port map (
            O => \N__1511\,
            I => \N__1508\
        );

    \I__308\ : Span12Mux_v
    port map (
            O => \N__1508\,
            I => \N__1505\
        );

    \I__307\ : Span12Mux_v
    port map (
            O => \N__1505\,
            I => \N__1502\
        );

    \I__306\ : Odrv12
    port map (
            O => \N__1502\,
            I => \AD0_c_7\
        );

    \I__305\ : IoInMux
    port map (
            O => \N__1499\,
            I => \N__1496\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__1496\,
            I => \N__1493\
        );

    \I__303\ : Span12Mux_s4_v
    port map (
            O => \N__1493\,
            I => \N__1490\
        );

    \I__302\ : Span12Mux_h
    port map (
            O => \N__1490\,
            I => \N__1487\
        );

    \I__301\ : Span12Mux_v
    port map (
            O => \N__1487\,
            I => \N__1484\
        );

    \I__300\ : Span12Mux_v
    port map (
            O => \N__1484\,
            I => \N__1481\
        );

    \I__299\ : Odrv12
    port map (
            O => \N__1481\,
            I => \AD2_c_0\
        );

    \I__298\ : IoInMux
    port map (
            O => \N__1478\,
            I => \N__1475\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__1475\,
            I => \N__1472\
        );

    \I__296\ : IoSpan4Mux
    port map (
            O => \N__1472\,
            I => \N__1469\
        );

    \I__295\ : Span4Mux_s3_h
    port map (
            O => \N__1469\,
            I => \N__1466\
        );

    \I__294\ : Sp12to4
    port map (
            O => \N__1466\,
            I => \N__1463\
        );

    \I__293\ : Span12Mux_v
    port map (
            O => \N__1463\,
            I => \N__1460\
        );

    \I__292\ : Span12Mux_v
    port map (
            O => \N__1460\,
            I => \N__1457\
        );

    \I__291\ : Span12Mux_h
    port map (
            O => \N__1457\,
            I => \N__1454\
        );

    \I__290\ : Span12Mux_h
    port map (
            O => \N__1454\,
            I => \N__1451\
        );

    \I__289\ : Odrv12
    port map (
            O => \N__1451\,
            I => \AD3_c_5\
        );

    \I__288\ : IoInMux
    port map (
            O => \N__1448\,
            I => \N__1445\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__1445\,
            I => \N__1442\
        );

    \I__286\ : Span4Mux_s2_v
    port map (
            O => \N__1442\,
            I => \N__1439\
        );

    \I__285\ : Sp12to4
    port map (
            O => \N__1439\,
            I => \N__1436\
        );

    \I__284\ : Span12Mux_h
    port map (
            O => \N__1436\,
            I => \N__1433\
        );

    \I__283\ : Span12Mux_h
    port map (
            O => \N__1433\,
            I => \N__1430\
        );

    \I__282\ : Odrv12
    port map (
            O => \N__1430\,
            I => \AD0_c_6\
        );

    \I__281\ : IoInMux
    port map (
            O => \N__1427\,
            I => \N__1424\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__1424\,
            I => \N__1421\
        );

    \I__279\ : Span12Mux_s11_v
    port map (
            O => \N__1421\,
            I => \N__1418\
        );

    \I__278\ : Span12Mux_h
    port map (
            O => \N__1418\,
            I => \N__1415\
        );

    \I__277\ : Odrv12
    port map (
            O => \N__1415\,
            I => \AD1_c_7\
        );

    \I__276\ : IoInMux
    port map (
            O => \N__1412\,
            I => \N__1409\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__1409\,
            I => \N__1406\
        );

    \I__274\ : Span12Mux_s9_h
    port map (
            O => \N__1406\,
            I => \N__1403\
        );

    \I__273\ : Span12Mux_v
    port map (
            O => \N__1403\,
            I => \N__1400\
        );

    \I__272\ : Span12Mux_v
    port map (
            O => \N__1400\,
            I => \N__1397\
        );

    \I__271\ : Span12Mux_h
    port map (
            O => \N__1397\,
            I => \N__1394\
        );

    \I__270\ : Odrv12
    port map (
            O => \N__1394\,
            I => \AD3_c_7\
        );

    \I__269\ : IoInMux
    port map (
            O => \N__1391\,
            I => \N__1388\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__1388\,
            I => \N__1385\
        );

    \I__267\ : IoSpan4Mux
    port map (
            O => \N__1385\,
            I => \N__1382\
        );

    \I__266\ : Span4Mux_s2_v
    port map (
            O => \N__1382\,
            I => \N__1379\
        );

    \I__265\ : Span4Mux_v
    port map (
            O => \N__1379\,
            I => \N__1376\
        );

    \I__264\ : Sp12to4
    port map (
            O => \N__1376\,
            I => \N__1373\
        );

    \I__263\ : Span12Mux_v
    port map (
            O => \N__1373\,
            I => \N__1370\
        );

    \I__262\ : Span12Mux_v
    port map (
            O => \N__1370\,
            I => \N__1367\
        );

    \I__261\ : Odrv12
    port map (
            O => \N__1367\,
            I => \AD2_c_1\
        );

    \I__260\ : IoInMux
    port map (
            O => \N__1364\,
            I => \N__1361\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__1361\,
            I => \N__1358\
        );

    \I__258\ : IoSpan4Mux
    port map (
            O => \N__1358\,
            I => \N__1355\
        );

    \I__257\ : Span4Mux_s2_v
    port map (
            O => \N__1355\,
            I => \N__1352\
        );

    \I__256\ : Sp12to4
    port map (
            O => \N__1352\,
            I => \N__1349\
        );

    \I__255\ : Span12Mux_h
    port map (
            O => \N__1349\,
            I => \N__1346\
        );

    \I__254\ : Span12Mux_h
    port map (
            O => \N__1346\,
            I => \N__1343\
        );

    \I__253\ : Odrv12
    port map (
            O => \N__1343\,
            I => \AD0_c_5\
        );

    \I__252\ : IoInMux
    port map (
            O => \N__1340\,
            I => \N__1337\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__1337\,
            I => \N__1334\
        );

    \I__250\ : IoSpan4Mux
    port map (
            O => \N__1334\,
            I => \N__1331\
        );

    \I__249\ : Span4Mux_s1_v
    port map (
            O => \N__1331\,
            I => \N__1328\
        );

    \I__248\ : Span4Mux_v
    port map (
            O => \N__1328\,
            I => \N__1325\
        );

    \I__247\ : Sp12to4
    port map (
            O => \N__1325\,
            I => \N__1322\
        );

    \I__246\ : Span12Mux_v
    port map (
            O => \N__1322\,
            I => \N__1319\
        );

    \I__245\ : Span12Mux_v
    port map (
            O => \N__1319\,
            I => \N__1316\
        );

    \I__244\ : Odrv12
    port map (
            O => \N__1316\,
            I => \AD2_c_2\
        );

    \I__243\ : IoInMux
    port map (
            O => \N__1313\,
            I => \N__1310\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__1310\,
            I => \N__1307\
        );

    \I__241\ : Span12Mux_s3_v
    port map (
            O => \N__1307\,
            I => \N__1304\
        );

    \I__240\ : Span12Mux_v
    port map (
            O => \N__1304\,
            I => \N__1301\
        );

    \I__239\ : Span12Mux_h
    port map (
            O => \N__1301\,
            I => \N__1298\
        );

    \I__238\ : Span12Mux_h
    port map (
            O => \N__1298\,
            I => \N__1295\
        );

    \I__237\ : Odrv12
    port map (
            O => \N__1295\,
            I => \AD1_c_4\
        );

    \I__236\ : IoInMux
    port map (
            O => \N__1292\,
            I => \N__1289\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__1289\,
            I => \N__1286\
        );

    \I__234\ : IoSpan4Mux
    port map (
            O => \N__1286\,
            I => \N__1283\
        );

    \I__233\ : Span4Mux_s1_h
    port map (
            O => \N__1283\,
            I => \N__1280\
        );

    \I__232\ : Sp12to4
    port map (
            O => \N__1280\,
            I => \N__1277\
        );

    \I__231\ : Span12Mux_s11_v
    port map (
            O => \N__1277\,
            I => \N__1274\
        );

    \I__230\ : Span12Mux_h
    port map (
            O => \N__1274\,
            I => \N__1271\
        );

    \I__229\ : Span12Mux_h
    port map (
            O => \N__1271\,
            I => \N__1268\
        );

    \I__228\ : Odrv12
    port map (
            O => \N__1268\,
            I => \AD0_c_0\
        );

    \I__227\ : IoInMux
    port map (
            O => \N__1265\,
            I => \N__1262\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1262\,
            I => \N__1259\
        );

    \I__225\ : Span4Mux_s0_v
    port map (
            O => \N__1259\,
            I => \N__1256\
        );

    \I__224\ : Span4Mux_v
    port map (
            O => \N__1256\,
            I => \N__1253\
        );

    \I__223\ : Sp12to4
    port map (
            O => \N__1253\,
            I => \N__1250\
        );

    \I__222\ : Span12Mux_h
    port map (
            O => \N__1250\,
            I => \N__1247\
        );

    \I__221\ : Span12Mux_v
    port map (
            O => \N__1247\,
            I => \N__1244\
        );

    \I__220\ : Span12Mux_h
    port map (
            O => \N__1244\,
            I => \N__1241\
        );

    \I__219\ : Odrv12
    port map (
            O => \N__1241\,
            I => \AD1_c_2\
        );

    \I__218\ : IoInMux
    port map (
            O => \N__1238\,
            I => \N__1235\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__1235\,
            I => \N__1232\
        );

    \I__216\ : IoSpan4Mux
    port map (
            O => \N__1232\,
            I => \N__1229\
        );

    \I__215\ : Span4Mux_s2_v
    port map (
            O => \N__1229\,
            I => \N__1226\
        );

    \I__214\ : Sp12to4
    port map (
            O => \N__1226\,
            I => \N__1223\
        );

    \I__213\ : Span12Mux_s10_v
    port map (
            O => \N__1223\,
            I => \N__1220\
        );

    \I__212\ : Span12Mux_v
    port map (
            O => \N__1220\,
            I => \N__1217\
        );

    \I__211\ : Odrv12
    port map (
            O => \N__1217\,
            I => \AD2_c_6\
        );

    \I__210\ : IoInMux
    port map (
            O => \N__1214\,
            I => \N__1211\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__1211\,
            I => \N__1208\
        );

    \I__208\ : IoSpan4Mux
    port map (
            O => \N__1208\,
            I => \N__1205\
        );

    \I__207\ : Span4Mux_s3_v
    port map (
            O => \N__1205\,
            I => \N__1202\
        );

    \I__206\ : Sp12to4
    port map (
            O => \N__1202\,
            I => \N__1199\
        );

    \I__205\ : Span12Mux_h
    port map (
            O => \N__1199\,
            I => \N__1196\
        );

    \I__204\ : Span12Mux_h
    port map (
            O => \N__1196\,
            I => \N__1193\
        );

    \I__203\ : Odrv12
    port map (
            O => \N__1193\,
            I => \AD0_c_4\
        );

    \I__202\ : IoInMux
    port map (
            O => \N__1190\,
            I => \N__1187\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__1187\,
            I => \N__1184\
        );

    \I__200\ : Span4Mux_s1_v
    port map (
            O => \N__1184\,
            I => \N__1181\
        );

    \I__199\ : Sp12to4
    port map (
            O => \N__1181\,
            I => \N__1178\
        );

    \I__198\ : Span12Mux_h
    port map (
            O => \N__1178\,
            I => \N__1175\
        );

    \I__197\ : Span12Mux_v
    port map (
            O => \N__1175\,
            I => \N__1172\
        );

    \I__196\ : Odrv12
    port map (
            O => \N__1172\,
            I => \AD1_c_5\
        );

    \I__195\ : IoInMux
    port map (
            O => \N__1169\,
            I => \N__1166\
        );

    \I__194\ : LocalMux
    port map (
            O => \N__1166\,
            I => \N__1163\
        );

    \I__193\ : Span4Mux_s3_v
    port map (
            O => \N__1163\,
            I => \N__1160\
        );

    \I__192\ : IoSpan4Mux
    port map (
            O => \N__1160\,
            I => \N__1157\
        );

    \I__191\ : IoSpan4Mux
    port map (
            O => \N__1157\,
            I => \N__1154\
        );

    \I__190\ : IoSpan4Mux
    port map (
            O => \N__1154\,
            I => \N__1151\
        );

    \I__189\ : IoSpan4Mux
    port map (
            O => \N__1151\,
            I => \N__1148\
        );

    \I__188\ : Odrv4
    port map (
            O => \N__1148\,
            I => \AD2_c_7\
        );

    \I__187\ : IoInMux
    port map (
            O => \N__1145\,
            I => \N__1142\
        );

    \I__186\ : LocalMux
    port map (
            O => \N__1142\,
            I => \N__1139\
        );

    \I__185\ : Span4Mux_s3_v
    port map (
            O => \N__1139\,
            I => \N__1136\
        );

    \I__184\ : Sp12to4
    port map (
            O => \N__1136\,
            I => \N__1133\
        );

    \I__183\ : Span12Mux_s3_h
    port map (
            O => \N__1133\,
            I => \N__1130\
        );

    \I__182\ : Span12Mux_v
    port map (
            O => \N__1130\,
            I => \N__1127\
        );

    \I__181\ : Span12Mux_v
    port map (
            O => \N__1127\,
            I => \N__1124\
        );

    \I__180\ : Odrv12
    port map (
            O => \N__1124\,
            I => \AD3_c_1\
        );

    \I__179\ : IoInMux
    port map (
            O => \N__1121\,
            I => \N__1118\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__1118\,
            I => \N__1115\
        );

    \I__177\ : IoSpan4Mux
    port map (
            O => \N__1115\,
            I => \N__1112\
        );

    \I__176\ : Span4Mux_s2_v
    port map (
            O => \N__1112\,
            I => \N__1109\
        );

    \I__175\ : Span4Mux_v
    port map (
            O => \N__1109\,
            I => \N__1106\
        );

    \I__174\ : Sp12to4
    port map (
            O => \N__1106\,
            I => \N__1103\
        );

    \I__173\ : Span12Mux_v
    port map (
            O => \N__1103\,
            I => \N__1100\
        );

    \I__172\ : Span12Mux_h
    port map (
            O => \N__1100\,
            I => \N__1097\
        );

    \I__171\ : Odrv12
    port map (
            O => \N__1097\,
            I => \AD1_c_3\
        );

    \I__170\ : IoInMux
    port map (
            O => \N__1094\,
            I => \N__1091\
        );

    \I__169\ : LocalMux
    port map (
            O => \N__1091\,
            I => \N__1088\
        );

    \I__168\ : Span12Mux_s4_v
    port map (
            O => \N__1088\,
            I => \N__1085\
        );

    \I__167\ : Span12Mux_h
    port map (
            O => \N__1085\,
            I => \N__1082\
        );

    \I__166\ : Span12Mux_h
    port map (
            O => \N__1082\,
            I => \N__1079\
        );

    \I__165\ : Odrv12
    port map (
            O => \N__1079\,
            I => \AD0_c_3\
        );

    \I__164\ : IoInMux
    port map (
            O => \N__1076\,
            I => \N__1073\
        );

    \I__163\ : LocalMux
    port map (
            O => \N__1073\,
            I => \N__1070\
        );

    \I__162\ : IoSpan4Mux
    port map (
            O => \N__1070\,
            I => \N__1067\
        );

    \I__161\ : Span4Mux_s3_h
    port map (
            O => \N__1067\,
            I => \N__1064\
        );

    \I__160\ : Sp12to4
    port map (
            O => \N__1064\,
            I => \N__1061\
        );

    \I__159\ : Span12Mux_v
    port map (
            O => \N__1061\,
            I => \N__1058\
        );

    \I__158\ : Span12Mux_h
    port map (
            O => \N__1058\,
            I => \N__1055\
        );

    \I__157\ : Span12Mux_h
    port map (
            O => \N__1055\,
            I => \N__1052\
        );

    \I__156\ : Odrv12
    port map (
            O => \N__1052\,
            I => \AD1_c_0\
        );

    \I__155\ : IoInMux
    port map (
            O => \N__1049\,
            I => \N__1046\
        );

    \I__154\ : LocalMux
    port map (
            O => \N__1046\,
            I => \N__1043\
        );

    \I__153\ : IoSpan4Mux
    port map (
            O => \N__1043\,
            I => \N__1040\
        );

    \I__152\ : Span4Mux_s2_h
    port map (
            O => \N__1040\,
            I => \N__1037\
        );

    \I__151\ : Sp12to4
    port map (
            O => \N__1037\,
            I => \N__1034\
        );

    \I__150\ : Span12Mux_h
    port map (
            O => \N__1034\,
            I => \N__1031\
        );

    \I__149\ : Span12Mux_v
    port map (
            O => \N__1031\,
            I => \N__1028\
        );

    \I__148\ : Span12Mux_v
    port map (
            O => \N__1028\,
            I => \N__1025\
        );

    \I__147\ : Span12Mux_h
    port map (
            O => \N__1025\,
            I => \N__1022\
        );

    \I__146\ : Odrv12
    port map (
            O => \N__1022\,
            I => \AD3_c_4\
        );

    \I__145\ : IoInMux
    port map (
            O => \N__1019\,
            I => \N__1016\
        );

    \I__144\ : LocalMux
    port map (
            O => \N__1016\,
            I => \N__1013\
        );

    \I__143\ : IoSpan4Mux
    port map (
            O => \N__1013\,
            I => \N__1010\
        );

    \I__142\ : Span4Mux_s2_v
    port map (
            O => \N__1010\,
            I => \N__1007\
        );

    \I__141\ : Sp12to4
    port map (
            O => \N__1007\,
            I => \N__1004\
        );

    \I__140\ : Span12Mux_v
    port map (
            O => \N__1004\,
            I => \N__1001\
        );

    \I__139\ : Span12Mux_v
    port map (
            O => \N__1001\,
            I => \N__998\
        );

    \I__138\ : Odrv12
    port map (
            O => \N__998\,
            I => \AD2_c_4\
        );

    \I__137\ : IoInMux
    port map (
            O => \N__995\,
            I => \N__992\
        );

    \I__136\ : LocalMux
    port map (
            O => \N__992\,
            I => \N__989\
        );

    \I__135\ : IoSpan4Mux
    port map (
            O => \N__989\,
            I => \N__986\
        );

    \I__134\ : Span4Mux_s0_v
    port map (
            O => \N__986\,
            I => \N__983\
        );

    \I__133\ : Span4Mux_v
    port map (
            O => \N__983\,
            I => \N__980\
        );

    \I__132\ : Sp12to4
    port map (
            O => \N__980\,
            I => \N__977\
        );

    \I__131\ : Span12Mux_v
    port map (
            O => \N__977\,
            I => \N__974\
        );

    \I__130\ : Span12Mux_v
    port map (
            O => \N__974\,
            I => \N__971\
        );

    \I__129\ : Odrv12
    port map (
            O => \N__971\,
            I => \AD2_c_5\
        );

    \I__128\ : IoInMux
    port map (
            O => \N__968\,
            I => \N__965\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__965\,
            I => \N__962\
        );

    \I__126\ : Span4Mux_s3_v
    port map (
            O => \N__962\,
            I => \N__959\
        );

    \I__125\ : Span4Mux_v
    port map (
            O => \N__959\,
            I => \N__956\
        );

    \I__124\ : Sp12to4
    port map (
            O => \N__956\,
            I => \N__953\
        );

    \I__123\ : Span12Mux_s0_h
    port map (
            O => \N__953\,
            I => \N__950\
        );

    \I__122\ : Span12Mux_v
    port map (
            O => \N__950\,
            I => \N__947\
        );

    \I__121\ : Span12Mux_v
    port map (
            O => \N__947\,
            I => \N__944\
        );

    \I__120\ : Odrv12
    port map (
            O => \N__944\,
            I => \AD3_c_3\
        );

    \I__119\ : IoInMux
    port map (
            O => \N__941\,
            I => \N__938\
        );

    \I__118\ : LocalMux
    port map (
            O => \N__938\,
            I => \N__935\
        );

    \I__117\ : IoSpan4Mux
    port map (
            O => \N__935\,
            I => \N__932\
        );

    \I__116\ : IoSpan4Mux
    port map (
            O => \N__932\,
            I => \N__929\
        );

    \I__115\ : Span4Mux_s2_h
    port map (
            O => \N__929\,
            I => \N__926\
        );

    \I__114\ : Sp12to4
    port map (
            O => \N__926\,
            I => \N__923\
        );

    \I__113\ : Span12Mux_h
    port map (
            O => \N__923\,
            I => \N__920\
        );

    \I__112\ : Span12Mux_h
    port map (
            O => \N__920\,
            I => \N__917\
        );

    \I__111\ : Odrv12
    port map (
            O => \N__917\,
            I => \AD0_c_1\
        );

    \I__110\ : IoInMux
    port map (
            O => \N__914\,
            I => \N__911\
        );

    \I__109\ : LocalMux
    port map (
            O => \N__911\,
            I => \N__908\
        );

    \I__108\ : Span4Mux_s0_v
    port map (
            O => \N__908\,
            I => \N__905\
        );

    \I__107\ : Sp12to4
    port map (
            O => \N__905\,
            I => \N__902\
        );

    \I__106\ : Span12Mux_h
    port map (
            O => \N__902\,
            I => \N__899\
        );

    \I__105\ : Span12Mux_v
    port map (
            O => \N__899\,
            I => \N__896\
        );

    \I__104\ : Odrv12
    port map (
            O => \N__896\,
            I => \AD1_c_6\
        );

    \I__103\ : IoInMux
    port map (
            O => \N__893\,
            I => \N__890\
        );

    \I__102\ : LocalMux
    port map (
            O => \N__890\,
            I => \N__887\
        );

    \I__101\ : IoSpan4Mux
    port map (
            O => \N__887\,
            I => \N__884\
        );

    \I__100\ : Span4Mux_s2_h
    port map (
            O => \N__884\,
            I => \N__881\
        );

    \I__99\ : Sp12to4
    port map (
            O => \N__881\,
            I => \N__878\
        );

    \I__98\ : Span12Mux_h
    port map (
            O => \N__878\,
            I => \N__875\
        );

    \I__97\ : Span12Mux_v
    port map (
            O => \N__875\,
            I => \N__872\
        );

    \I__96\ : Span12Mux_v
    port map (
            O => \N__872\,
            I => \N__869\
        );

    \I__95\ : Span12Mux_h
    port map (
            O => \N__869\,
            I => \N__866\
        );

    \I__94\ : Odrv12
    port map (
            O => \N__866\,
            I => \AD3_c_6\
        );

    \I__93\ : IoInMux
    port map (
            O => \N__863\,
            I => \N__860\
        );

    \I__92\ : LocalMux
    port map (
            O => \N__860\,
            I => \N__857\
        );

    \I__91\ : Span12Mux_s3_v
    port map (
            O => \N__857\,
            I => \N__854\
        );

    \I__90\ : Span12Mux_v
    port map (
            O => \N__854\,
            I => \N__851\
        );

    \I__89\ : Span12Mux_v
    port map (
            O => \N__851\,
            I => \N__848\
        );

    \I__88\ : Odrv12
    port map (
            O => \N__848\,
            I => \AD2_c_3\
        );

    \I__87\ : IoInMux
    port map (
            O => \N__845\,
            I => \N__842\
        );

    \I__86\ : LocalMux
    port map (
            O => \N__842\,
            I => \N__839\
        );

    \I__85\ : IoSpan4Mux
    port map (
            O => \N__839\,
            I => \N__836\
        );

    \I__84\ : Span4Mux_s3_v
    port map (
            O => \N__836\,
            I => \N__833\
        );

    \I__83\ : Sp12to4
    port map (
            O => \N__833\,
            I => \N__830\
        );

    \I__82\ : Span12Mux_s11_v
    port map (
            O => \N__830\,
            I => \N__827\
        );

    \I__81\ : Span12Mux_v
    port map (
            O => \N__827\,
            I => \N__824\
        );

    \I__80\ : Odrv12
    port map (
            O => \N__824\,
            I => \AD3_c_0\
        );

    \I__79\ : IoInMux
    port map (
            O => \N__821\,
            I => \N__818\
        );

    \I__78\ : LocalMux
    port map (
            O => \N__818\,
            I => \N__815\
        );

    \I__77\ : Span4Mux_s1_v
    port map (
            O => \N__815\,
            I => \N__812\
        );

    \I__76\ : Span4Mux_v
    port map (
            O => \N__812\,
            I => \N__809\
        );

    \I__75\ : Sp12to4
    port map (
            O => \N__809\,
            I => \N__806\
        );

    \I__74\ : Span12Mux_h
    port map (
            O => \N__806\,
            I => \N__803\
        );

    \I__73\ : Span12Mux_h
    port map (
            O => \N__803\,
            I => \N__800\
        );

    \I__72\ : Odrv12
    port map (
            O => \N__800\,
            I => \AD0_c_2\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 15 2024 12:53:28

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    CMA,
    DRA,
    A,
    TSn,
    CLMBEn,
    AWEn,
    RESETn,
    CASn,
    BANK0,
    VBENn,
    CUMBEn,
    CLKRAM,
    C3,
    ASn,
    LDSn,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    DBRn,
    CLK40C,
    CLK40_IN,
    REGSPACEn,
    RAMENn,
    RASn,
    TACKn,
    CLKEN,
    C1);

    input [1:0] SIZ;
    output [10:0] CMA;
    input [9:0] DRA;
    input [20:0] A;
    input TSn;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CASn;
    output BANK0;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    input C3;
    output ASn;
    output LDSn;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    input DBRn;
    output CLK40C;
    input CLK40_IN;
    input REGSPACEn;
    output RAMENn;
    output RASn;
    output TACKn;
    output CLKEN;
    input C1;

    wire N__10331;
    wire N__10330;
    wire N__10329;
    wire N__10322;
    wire N__10321;
    wire N__10320;
    wire N__10313;
    wire N__10312;
    wire N__10311;
    wire N__10304;
    wire N__10303;
    wire N__10302;
    wire N__10295;
    wire N__10294;
    wire N__10293;
    wire N__10286;
    wire N__10285;
    wire N__10284;
    wire N__10277;
    wire N__10276;
    wire N__10275;
    wire N__10268;
    wire N__10267;
    wire N__10266;
    wire N__10259;
    wire N__10258;
    wire N__10257;
    wire N__10250;
    wire N__10249;
    wire N__10248;
    wire N__10241;
    wire N__10240;
    wire N__10239;
    wire N__10232;
    wire N__10231;
    wire N__10230;
    wire N__10223;
    wire N__10222;
    wire N__10221;
    wire N__10214;
    wire N__10213;
    wire N__10212;
    wire N__10205;
    wire N__10204;
    wire N__10203;
    wire N__10196;
    wire N__10195;
    wire N__10194;
    wire N__10187;
    wire N__10186;
    wire N__10185;
    wire N__10178;
    wire N__10177;
    wire N__10176;
    wire N__10169;
    wire N__10168;
    wire N__10167;
    wire N__10160;
    wire N__10159;
    wire N__10158;
    wire N__10151;
    wire N__10150;
    wire N__10149;
    wire N__10142;
    wire N__10141;
    wire N__10140;
    wire N__10133;
    wire N__10132;
    wire N__10131;
    wire N__10124;
    wire N__10123;
    wire N__10122;
    wire N__10115;
    wire N__10114;
    wire N__10113;
    wire N__10106;
    wire N__10105;
    wire N__10104;
    wire N__10097;
    wire N__10096;
    wire N__10095;
    wire N__10088;
    wire N__10087;
    wire N__10086;
    wire N__10079;
    wire N__10078;
    wire N__10077;
    wire N__10070;
    wire N__10069;
    wire N__10068;
    wire N__10061;
    wire N__10060;
    wire N__10059;
    wire N__10052;
    wire N__10051;
    wire N__10050;
    wire N__10043;
    wire N__10042;
    wire N__10041;
    wire N__10034;
    wire N__10033;
    wire N__10032;
    wire N__10025;
    wire N__10024;
    wire N__10023;
    wire N__10016;
    wire N__10015;
    wire N__10014;
    wire N__10007;
    wire N__10006;
    wire N__10005;
    wire N__9998;
    wire N__9997;
    wire N__9996;
    wire N__9989;
    wire N__9988;
    wire N__9987;
    wire N__9980;
    wire N__9979;
    wire N__9978;
    wire N__9971;
    wire N__9970;
    wire N__9969;
    wire N__9962;
    wire N__9961;
    wire N__9960;
    wire N__9953;
    wire N__9952;
    wire N__9951;
    wire N__9944;
    wire N__9943;
    wire N__9942;
    wire N__9935;
    wire N__9934;
    wire N__9933;
    wire N__9926;
    wire N__9925;
    wire N__9924;
    wire N__9917;
    wire N__9916;
    wire N__9915;
    wire N__9908;
    wire N__9907;
    wire N__9906;
    wire N__9899;
    wire N__9898;
    wire N__9897;
    wire N__9890;
    wire N__9889;
    wire N__9888;
    wire N__9881;
    wire N__9880;
    wire N__9879;
    wire N__9872;
    wire N__9871;
    wire N__9870;
    wire N__9863;
    wire N__9862;
    wire N__9861;
    wire N__9854;
    wire N__9853;
    wire N__9852;
    wire N__9845;
    wire N__9844;
    wire N__9843;
    wire N__9836;
    wire N__9835;
    wire N__9834;
    wire N__9827;
    wire N__9826;
    wire N__9825;
    wire N__9818;
    wire N__9817;
    wire N__9816;
    wire N__9809;
    wire N__9808;
    wire N__9807;
    wire N__9800;
    wire N__9799;
    wire N__9798;
    wire N__9791;
    wire N__9790;
    wire N__9789;
    wire N__9782;
    wire N__9781;
    wire N__9780;
    wire N__9773;
    wire N__9772;
    wire N__9771;
    wire N__9764;
    wire N__9763;
    wire N__9762;
    wire N__9755;
    wire N__9754;
    wire N__9753;
    wire N__9746;
    wire N__9745;
    wire N__9744;
    wire N__9737;
    wire N__9736;
    wire N__9735;
    wire N__9728;
    wire N__9727;
    wire N__9726;
    wire N__9719;
    wire N__9718;
    wire N__9717;
    wire N__9710;
    wire N__9709;
    wire N__9708;
    wire N__9701;
    wire N__9700;
    wire N__9699;
    wire N__9692;
    wire N__9691;
    wire N__9690;
    wire N__9683;
    wire N__9682;
    wire N__9681;
    wire N__9674;
    wire N__9673;
    wire N__9672;
    wire N__9665;
    wire N__9664;
    wire N__9663;
    wire N__9656;
    wire N__9655;
    wire N__9654;
    wire N__9647;
    wire N__9646;
    wire N__9645;
    wire N__9638;
    wire N__9637;
    wire N__9636;
    wire N__9629;
    wire N__9628;
    wire N__9627;
    wire N__9620;
    wire N__9619;
    wire N__9618;
    wire N__9601;
    wire N__9598;
    wire N__9595;
    wire N__9592;
    wire N__9591;
    wire N__9588;
    wire N__9585;
    wire N__9582;
    wire N__9577;
    wire N__9574;
    wire N__9573;
    wire N__9572;
    wire N__9571;
    wire N__9570;
    wire N__9569;
    wire N__9568;
    wire N__9567;
    wire N__9566;
    wire N__9565;
    wire N__9564;
    wire N__9563;
    wire N__9562;
    wire N__9561;
    wire N__9560;
    wire N__9559;
    wire N__9558;
    wire N__9557;
    wire N__9556;
    wire N__9555;
    wire N__9554;
    wire N__9553;
    wire N__9552;
    wire N__9551;
    wire N__9550;
    wire N__9549;
    wire N__9548;
    wire N__9547;
    wire N__9546;
    wire N__9545;
    wire N__9544;
    wire N__9543;
    wire N__9542;
    wire N__9541;
    wire N__9540;
    wire N__9539;
    wire N__9538;
    wire N__9535;
    wire N__9534;
    wire N__9533;
    wire N__9532;
    wire N__9531;
    wire N__9530;
    wire N__9529;
    wire N__9528;
    wire N__9527;
    wire N__9526;
    wire N__9525;
    wire N__9524;
    wire N__9523;
    wire N__9522;
    wire N__9421;
    wire N__9418;
    wire N__9417;
    wire N__9416;
    wire N__9415;
    wire N__9414;
    wire N__9413;
    wire N__9412;
    wire N__9411;
    wire N__9410;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9381;
    wire N__9380;
    wire N__9379;
    wire N__9378;
    wire N__9377;
    wire N__9376;
    wire N__9375;
    wire N__9374;
    wire N__9371;
    wire N__9370;
    wire N__9369;
    wire N__9368;
    wire N__9367;
    wire N__9366;
    wire N__9365;
    wire N__9364;
    wire N__9363;
    wire N__9360;
    wire N__9359;
    wire N__9358;
    wire N__9357;
    wire N__9356;
    wire N__9355;
    wire N__9354;
    wire N__9353;
    wire N__9352;
    wire N__9351;
    wire N__9350;
    wire N__9349;
    wire N__9346;
    wire N__9345;
    wire N__9344;
    wire N__9341;
    wire N__9340;
    wire N__9339;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9331;
    wire N__9330;
    wire N__9329;
    wire N__9328;
    wire N__9325;
    wire N__9324;
    wire N__9323;
    wire N__9322;
    wire N__9321;
    wire N__9320;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9192;
    wire N__9189;
    wire N__9184;
    wire N__9181;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9173;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9159;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9142;
    wire N__9141;
    wire N__9140;
    wire N__9139;
    wire N__9136;
    wire N__9133;
    wire N__9130;
    wire N__9127;
    wire N__9126;
    wire N__9125;
    wire N__9124;
    wire N__9123;
    wire N__9122;
    wire N__9119;
    wire N__9114;
    wire N__9111;
    wire N__9102;
    wire N__9099;
    wire N__9094;
    wire N__9085;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9063;
    wire N__9060;
    wire N__9059;
    wire N__9058;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9045;
    wire N__9042;
    wire N__9037;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9012;
    wire N__9007;
    wire N__9004;
    wire N__9003;
    wire N__9000;
    wire N__8997;
    wire N__8994;
    wire N__8991;
    wire N__8988;
    wire N__8985;
    wire N__8982;
    wire N__8979;
    wire N__8976;
    wire N__8973;
    wire N__8968;
    wire N__8965;
    wire N__8962;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8935;
    wire N__8934;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8887;
    wire N__8886;
    wire N__8883;
    wire N__8880;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8866;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8847;
    wire N__8844;
    wire N__8839;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8820;
    wire N__8819;
    wire N__8818;
    wire N__8817;
    wire N__8816;
    wire N__8813;
    wire N__8812;
    wire N__8811;
    wire N__8808;
    wire N__8805;
    wire N__8802;
    wire N__8801;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8787;
    wire N__8782;
    wire N__8781;
    wire N__8778;
    wire N__8773;
    wire N__8770;
    wire N__8769;
    wire N__8768;
    wire N__8761;
    wire N__8758;
    wire N__8755;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8738;
    wire N__8733;
    wire N__8722;
    wire N__8719;
    wire N__8716;
    wire N__8713;
    wire N__8710;
    wire N__8707;
    wire N__8704;
    wire N__8703;
    wire N__8702;
    wire N__8701;
    wire N__8700;
    wire N__8699;
    wire N__8696;
    wire N__8695;
    wire N__8692;
    wire N__8691;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8680;
    wire N__8677;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8644;
    wire N__8641;
    wire N__8638;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8622;
    wire N__8617;
    wire N__8616;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8598;
    wire N__8589;
    wire N__8584;
    wire N__8575;
    wire N__8566;
    wire N__8563;
    wire N__8560;
    wire N__8557;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8541;
    wire N__8540;
    wire N__8539;
    wire N__8538;
    wire N__8535;
    wire N__8534;
    wire N__8531;
    wire N__8530;
    wire N__8527;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8517;
    wire N__8516;
    wire N__8515;
    wire N__8512;
    wire N__8511;
    wire N__8510;
    wire N__8507;
    wire N__8500;
    wire N__8497;
    wire N__8494;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8472;
    wire N__8469;
    wire N__8468;
    wire N__8467;
    wire N__8460;
    wire N__8457;
    wire N__8448;
    wire N__8443;
    wire N__8440;
    wire N__8431;
    wire N__8428;
    wire N__8425;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8388;
    wire N__8385;
    wire N__8380;
    wire N__8377;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8365;
    wire N__8364;
    wire N__8363;
    wire N__8358;
    wire N__8355;
    wire N__8350;
    wire N__8349;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8328;
    wire N__8323;
    wire N__8322;
    wire N__8321;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8309;
    wire N__8302;
    wire N__8299;
    wire N__8298;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8271;
    wire N__8268;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8251;
    wire N__8250;
    wire N__8249;
    wire N__8248;
    wire N__8245;
    wire N__8240;
    wire N__8235;
    wire N__8232;
    wire N__8229;
    wire N__8218;
    wire N__8215;
    wire N__8214;
    wire N__8211;
    wire N__8208;
    wire N__8205;
    wire N__8200;
    wire N__8199;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8179;
    wire N__8178;
    wire N__8175;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8163;
    wire N__8160;
    wire N__8155;
    wire N__8150;
    wire N__8147;
    wire N__8142;
    wire N__8139;
    wire N__8136;
    wire N__8131;
    wire N__8128;
    wire N__8127;
    wire N__8124;
    wire N__8123;
    wire N__8122;
    wire N__8121;
    wire N__8120;
    wire N__8119;
    wire N__8118;
    wire N__8117;
    wire N__8116;
    wire N__8113;
    wire N__8110;
    wire N__8109;
    wire N__8106;
    wire N__8105;
    wire N__8104;
    wire N__8103;
    wire N__8100;
    wire N__8099;
    wire N__8098;
    wire N__8097;
    wire N__8096;
    wire N__8093;
    wire N__8092;
    wire N__8091;
    wire N__8090;
    wire N__8089;
    wire N__8088;
    wire N__8079;
    wire N__8076;
    wire N__8075;
    wire N__8070;
    wire N__8067;
    wire N__8066;
    wire N__8065;
    wire N__8062;
    wire N__8057;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8043;
    wire N__8040;
    wire N__8037;
    wire N__8028;
    wire N__8025;
    wire N__8024;
    wire N__8023;
    wire N__8020;
    wire N__8017;
    wire N__8014;
    wire N__8009;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7980;
    wire N__7977;
    wire N__7974;
    wire N__7971;
    wire N__7962;
    wire N__7953;
    wire N__7944;
    wire N__7933;
    wire N__7930;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7917;
    wire N__7914;
    wire N__7911;
    wire N__7908;
    wire N__7905;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7887;
    wire N__7884;
    wire N__7883;
    wire N__7882;
    wire N__7881;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7867;
    wire N__7864;
    wire N__7855;
    wire N__7854;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7844;
    wire N__7841;
    wire N__7840;
    wire N__7839;
    wire N__7836;
    wire N__7833;
    wire N__7830;
    wire N__7825;
    wire N__7816;
    wire N__7815;
    wire N__7812;
    wire N__7809;
    wire N__7808;
    wire N__7803;
    wire N__7800;
    wire N__7799;
    wire N__7798;
    wire N__7797;
    wire N__7796;
    wire N__7795;
    wire N__7792;
    wire N__7789;
    wire N__7784;
    wire N__7781;
    wire N__7780;
    wire N__7777;
    wire N__7774;
    wire N__7767;
    wire N__7764;
    wire N__7761;
    wire N__7758;
    wire N__7755;
    wire N__7754;
    wire N__7753;
    wire N__7752;
    wire N__7747;
    wire N__7744;
    wire N__7739;
    wire N__7734;
    wire N__7731;
    wire N__7728;
    wire N__7719;
    wire N__7716;
    wire N__7713;
    wire N__7708;
    wire N__7707;
    wire N__7706;
    wire N__7703;
    wire N__7702;
    wire N__7701;
    wire N__7696;
    wire N__7693;
    wire N__7688;
    wire N__7685;
    wire N__7684;
    wire N__7683;
    wire N__7682;
    wire N__7681;
    wire N__7680;
    wire N__7679;
    wire N__7678;
    wire N__7677;
    wire N__7674;
    wire N__7669;
    wire N__7664;
    wire N__7661;
    wire N__7654;
    wire N__7649;
    wire N__7646;
    wire N__7633;
    wire N__7630;
    wire N__7629;
    wire N__7628;
    wire N__7625;
    wire N__7624;
    wire N__7621;
    wire N__7616;
    wire N__7615;
    wire N__7612;
    wire N__7611;
    wire N__7610;
    wire N__7609;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7592;
    wire N__7589;
    wire N__7576;
    wire N__7575;
    wire N__7572;
    wire N__7571;
    wire N__7570;
    wire N__7569;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7543;
    wire N__7542;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7525;
    wire N__7524;
    wire N__7523;
    wire N__7522;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7514;
    wire N__7513;
    wire N__7510;
    wire N__7507;
    wire N__7502;
    wire N__7499;
    wire N__7494;
    wire N__7483;
    wire N__7480;
    wire N__7477;
    wire N__7474;
    wire N__7471;
    wire N__7468;
    wire N__7467;
    wire N__7464;
    wire N__7461;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7435;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7411;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7399;
    wire N__7396;
    wire N__7395;
    wire N__7394;
    wire N__7393;
    wire N__7392;
    wire N__7389;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7379;
    wire N__7376;
    wire N__7373;
    wire N__7368;
    wire N__7365;
    wire N__7362;
    wire N__7359;
    wire N__7354;
    wire N__7351;
    wire N__7348;
    wire N__7345;
    wire N__7342;
    wire N__7339;
    wire N__7330;
    wire N__7329;
    wire N__7326;
    wire N__7323;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7309;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7293;
    wire N__7290;
    wire N__7287;
    wire N__7284;
    wire N__7281;
    wire N__7278;
    wire N__7275;
    wire N__7272;
    wire N__7269;
    wire N__7264;
    wire N__7261;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7251;
    wire N__7248;
    wire N__7245;
    wire N__7240;
    wire N__7237;
    wire N__7236;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7219;
    wire N__7218;
    wire N__7217;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7207;
    wire N__7204;
    wire N__7199;
    wire N__7198;
    wire N__7197;
    wire N__7194;
    wire N__7193;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7181;
    wire N__7178;
    wire N__7173;
    wire N__7162;
    wire N__7159;
    wire N__7156;
    wire N__7153;
    wire N__7150;
    wire N__7147;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7134;
    wire N__7131;
    wire N__7128;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7116;
    wire N__7113;
    wire N__7112;
    wire N__7111;
    wire N__7108;
    wire N__7105;
    wire N__7102;
    wire N__7099;
    wire N__7090;
    wire N__7089;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7066;
    wire N__7065;
    wire N__7062;
    wire N__7061;
    wire N__7060;
    wire N__7055;
    wire N__7052;
    wire N__7049;
    wire N__7042;
    wire N__7041;
    wire N__7036;
    wire N__7033;
    wire N__7030;
    wire N__7027;
    wire N__7026;
    wire N__7025;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7015;
    wire N__7014;
    wire N__7009;
    wire N__7006;
    wire N__7003;
    wire N__7000;
    wire N__6991;
    wire N__6990;
    wire N__6985;
    wire N__6982;
    wire N__6981;
    wire N__6978;
    wire N__6977;
    wire N__6976;
    wire N__6975;
    wire N__6974;
    wire N__6973;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6963;
    wire N__6960;
    wire N__6959;
    wire N__6958;
    wire N__6957;
    wire N__6956;
    wire N__6955;
    wire N__6954;
    wire N__6951;
    wire N__6948;
    wire N__6947;
    wire N__6944;
    wire N__6941;
    wire N__6938;
    wire N__6935;
    wire N__6932;
    wire N__6929;
    wire N__6926;
    wire N__6921;
    wire N__6916;
    wire N__6907;
    wire N__6886;
    wire N__6885;
    wire N__6882;
    wire N__6879;
    wire N__6874;
    wire N__6873;
    wire N__6872;
    wire N__6869;
    wire N__6868;
    wire N__6865;
    wire N__6864;
    wire N__6863;
    wire N__6862;
    wire N__6861;
    wire N__6858;
    wire N__6857;
    wire N__6856;
    wire N__6855;
    wire N__6854;
    wire N__6853;
    wire N__6848;
    wire N__6847;
    wire N__6846;
    wire N__6843;
    wire N__6838;
    wire N__6837;
    wire N__6834;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6820;
    wire N__6817;
    wire N__6814;
    wire N__6811;
    wire N__6808;
    wire N__6807;
    wire N__6806;
    wire N__6805;
    wire N__6804;
    wire N__6801;
    wire N__6796;
    wire N__6791;
    wire N__6788;
    wire N__6781;
    wire N__6776;
    wire N__6771;
    wire N__6762;
    wire N__6745;
    wire N__6744;
    wire N__6743;
    wire N__6740;
    wire N__6735;
    wire N__6732;
    wire N__6729;
    wire N__6726;
    wire N__6723;
    wire N__6720;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6708;
    wire N__6703;
    wire N__6702;
    wire N__6697;
    wire N__6696;
    wire N__6693;
    wire N__6690;
    wire N__6687;
    wire N__6684;
    wire N__6679;
    wire N__6676;
    wire N__6673;
    wire N__6670;
    wire N__6669;
    wire N__6666;
    wire N__6665;
    wire N__6662;
    wire N__6657;
    wire N__6652;
    wire N__6651;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6616;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6585;
    wire N__6584;
    wire N__6579;
    wire N__6576;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6549;
    wire N__6546;
    wire N__6543;
    wire N__6540;
    wire N__6537;
    wire N__6534;
    wire N__6531;
    wire N__6528;
    wire N__6525;
    wire N__6522;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6504;
    wire N__6501;
    wire N__6498;
    wire N__6493;
    wire N__6490;
    wire N__6487;
    wire N__6486;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6426;
    wire N__6423;
    wire N__6420;
    wire N__6415;
    wire N__6412;
    wire N__6411;
    wire N__6408;
    wire N__6405;
    wire N__6404;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6388;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6380;
    wire N__6379;
    wire N__6378;
    wire N__6377;
    wire N__6372;
    wire N__6369;
    wire N__6366;
    wire N__6363;
    wire N__6360;
    wire N__6355;
    wire N__6352;
    wire N__6343;
    wire N__6340;
    wire N__6337;
    wire N__6336;
    wire N__6333;
    wire N__6330;
    wire N__6327;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6312;
    wire N__6309;
    wire N__6306;
    wire N__6305;
    wire N__6300;
    wire N__6297;
    wire N__6292;
    wire N__6289;
    wire N__6288;
    wire N__6285;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6271;
    wire N__6268;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6247;
    wire N__6244;
    wire N__6241;
    wire N__6240;
    wire N__6237;
    wire N__6234;
    wire N__6229;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6193;
    wire N__6190;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6175;
    wire N__6172;
    wire N__6169;
    wire N__6166;
    wire N__6163;
    wire N__6160;
    wire N__6157;
    wire N__6154;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6124;
    wire N__6123;
    wire N__6120;
    wire N__6117;
    wire N__6114;
    wire N__6111;
    wire N__6106;
    wire N__6103;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6081;
    wire N__6078;
    wire N__6075;
    wire N__6070;
    wire N__6069;
    wire N__6066;
    wire N__6063;
    wire N__6058;
    wire N__6055;
    wire N__6054;
    wire N__6053;
    wire N__6050;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6037;
    wire N__6034;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__5998;
    wire N__5995;
    wire N__5992;
    wire N__5989;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5977;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5947;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5881;
    wire N__5878;
    wire N__5875;
    wire N__5872;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5856;
    wire N__5853;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5815;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5788;
    wire N__5785;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5772;
    wire N__5771;
    wire N__5770;
    wire N__5769;
    wire N__5768;
    wire N__5765;
    wire N__5756;
    wire N__5753;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5713;
    wire N__5710;
    wire N__5709;
    wire N__5706;
    wire N__5703;
    wire N__5698;
    wire N__5695;
    wire N__5694;
    wire N__5691;
    wire N__5688;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5676;
    wire N__5673;
    wire N__5670;
    wire N__5667;
    wire N__5662;
    wire N__5659;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5647;
    wire N__5644;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5616;
    wire N__5613;
    wire N__5610;
    wire N__5605;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5565;
    wire N__5560;
    wire N__5557;
    wire N__5554;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5509;
    wire N__5508;
    wire N__5507;
    wire N__5506;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5478;
    wire N__5477;
    wire N__5476;
    wire N__5475;
    wire N__5470;
    wire N__5467;
    wire N__5462;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5448;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5436;
    wire N__5435;
    wire N__5434;
    wire N__5431;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5403;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5236;
    wire N__5233;
    wire N__5230;
    wire N__5227;
    wire N__5224;
    wire N__5221;
    wire N__5218;
    wire N__5215;
    wire N__5212;
    wire N__5209;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5191;
    wire N__5188;
    wire N__5185;
    wire N__5184;
    wire N__5181;
    wire N__5178;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5148;
    wire N__5145;
    wire N__5142;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5130;
    wire N__5127;
    wire N__5124;
    wire N__5121;
    wire N__5118;
    wire N__5113;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5101;
    wire N__5098;
    wire N__5095;
    wire N__5092;
    wire N__5089;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5044;
    wire N__5043;
    wire N__5040;
    wire N__5039;
    wire N__5038;
    wire N__5037;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5017;
    wire N__5014;
    wire N__5007;
    wire N__5002;
    wire N__4999;
    wire N__4996;
    wire N__4993;
    wire N__4990;
    wire N__4987;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4948;
    wire N__4945;
    wire N__4940;
    wire N__4937;
    wire N__4930;
    wire N__4929;
    wire N__4926;
    wire N__4923;
    wire N__4918;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4906;
    wire N__4903;
    wire N__4902;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4879;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4852;
    wire N__4849;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4822;
    wire N__4819;
    wire N__4816;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4804;
    wire N__4801;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4777;
    wire N__4774;
    wire N__4771;
    wire N__4768;
    wire N__4765;
    wire N__4762;
    wire N__4759;
    wire N__4756;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4744;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4734;
    wire N__4733;
    wire N__4730;
    wire N__4727;
    wire N__4724;
    wire N__4717;
    wire N__4714;
    wire N__4713;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4680;
    wire N__4677;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4659;
    wire N__4654;
    wire N__4653;
    wire N__4652;
    wire N__4647;
    wire N__4644;
    wire N__4639;
    wire N__4636;
    wire N__4633;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4615;
    wire N__4612;
    wire N__4609;
    wire N__4606;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4573;
    wire N__4570;
    wire N__4567;
    wire N__4564;
    wire N__4561;
    wire N__4558;
    wire N__4555;
    wire N__4552;
    wire N__4549;
    wire N__4546;
    wire N__4543;
    wire N__4540;
    wire N__4537;
    wire N__4534;
    wire N__4531;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4474;
    wire N__4471;
    wire N__4470;
    wire N__4467;
    wire N__4464;
    wire N__4459;
    wire N__4456;
    wire N__4455;
    wire N__4454;
    wire N__4451;
    wire N__4446;
    wire N__4441;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4429;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4401;
    wire N__4398;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4381;
    wire N__4378;
    wire N__4377;
    wire N__4372;
    wire N__4369;
    wire N__4366;
    wire N__4363;
    wire N__4360;
    wire N__4357;
    wire N__4354;
    wire N__4353;
    wire N__4348;
    wire N__4345;
    wire N__4344;
    wire N__4343;
    wire N__4336;
    wire N__4333;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4316;
    wire N__4311;
    wire N__4308;
    wire N__4303;
    wire N__4300;
    wire N__4297;
    wire N__4294;
    wire N__4291;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4267;
    wire N__4266;
    wire N__4265;
    wire N__4264;
    wire N__4263;
    wire N__4258;
    wire N__4253;
    wire N__4250;
    wire N__4243;
    wire N__4242;
    wire N__4241;
    wire N__4240;
    wire N__4239;
    wire N__4236;
    wire N__4229;
    wire N__4226;
    wire N__4219;
    wire N__4216;
    wire N__4215;
    wire N__4214;
    wire N__4213;
    wire N__4210;
    wire N__4205;
    wire N__4202;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4188;
    wire N__4185;
    wire N__4184;
    wire N__4179;
    wire N__4176;
    wire N__4171;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4159;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4144;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4129;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4117;
    wire N__4114;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4102;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire N__4083;
    wire N__4082;
    wire N__4079;
    wire N__4074;
    wire N__4069;
    wire N__4066;
    wire N__4065;
    wire N__4064;
    wire N__4061;
    wire N__4056;
    wire N__4051;
    wire N__4048;
    wire N__4045;
    wire N__4042;
    wire N__4041;
    wire N__4038;
    wire N__4035;
    wire N__4030;
    wire N__4027;
    wire N__4024;
    wire N__4023;
    wire N__4022;
    wire N__4021;
    wire N__4020;
    wire N__4019;
    wire N__4018;
    wire N__4017;
    wire N__4014;
    wire N__4009;
    wire N__4006;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3986;
    wire N__3979;
    wire N__3978;
    wire N__3977;
    wire N__3976;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3958;
    wire N__3957;
    wire N__3956;
    wire N__3953;
    wire N__3952;
    wire N__3951;
    wire N__3948;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3928;
    wire N__3925;
    wire N__3924;
    wire N__3923;
    wire N__3922;
    wire N__3919;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3900;
    wire N__3897;
    wire N__3894;
    wire N__3889;
    wire N__3886;
    wire N__3885;
    wire N__3884;
    wire N__3883;
    wire N__3874;
    wire N__3871;
    wire N__3870;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3853;
    wire N__3852;
    wire N__3849;
    wire N__3846;
    wire N__3843;
    wire N__3840;
    wire N__3835;
    wire N__3834;
    wire N__3833;
    wire N__3832;
    wire N__3829;
    wire N__3826;
    wire N__3823;
    wire N__3818;
    wire N__3813;
    wire N__3808;
    wire N__3805;
    wire N__3802;
    wire N__3799;
    wire N__3796;
    wire N__3793;
    wire N__3790;
    wire N__3787;
    wire N__3784;
    wire N__3781;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3773;
    wire N__3770;
    wire N__3767;
    wire N__3764;
    wire N__3757;
    wire N__3754;
    wire N__3753;
    wire N__3750;
    wire N__3747;
    wire N__3742;
    wire N__3739;
    wire N__3736;
    wire N__3733;
    wire N__3730;
    wire N__3727;
    wire N__3724;
    wire N__3723;
    wire N__3720;
    wire N__3717;
    wire N__3712;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3696;
    wire N__3691;
    wire N__3688;
    wire N__3685;
    wire N__3682;
    wire N__3679;
    wire N__3676;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3664;
    wire N__3661;
    wire N__3658;
    wire N__3655;
    wire N__3652;
    wire N__3649;
    wire N__3646;
    wire N__3643;
    wire N__3640;
    wire N__3637;
    wire N__3634;
    wire N__3631;
    wire N__3628;
    wire N__3625;
    wire N__3622;
    wire N__3619;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3607;
    wire N__3604;
    wire N__3601;
    wire N__3598;
    wire N__3595;
    wire N__3592;
    wire N__3589;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_OUT_i_i;
    wire CLK40_OUT_i_i;
    wire \U712_REG_SM.N_120 ;
    wire C3_c;
    wire N_677_i;
    wire TACK_EN_i_ess;
    wire \U712_REG_SM.N_86 ;
    wire \U712_REG_SM.N_68_cascade_ ;
    wire \U712_REG_SM.N_73_cascade_ ;
    wire TACK_OUTn;
    wire C1_c;
    wire CLK40_OUT_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.N_45_0_0_en_cascade_ ;
    wire \U712_CYCLE_TERM.N_45_0_0_en_0 ;
    wire VBENn_c;
    wire \U712_REG_SM.N_73 ;
    wire \U712_REG_SM.un1_STATE_COUNT_5_0_1_cascade_ ;
    wire CPU_TACKm;
    wire \U712_REG_SM.STATE_COUNTZ0Z_5 ;
    wire \U712_REG_SM.N_173_0_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.N_54_cascade_ ;
    wire \U712_REG_SM.un1_STATE_COUNT_5_0_1 ;
    wire REG_TACK;
    wire \U712_REG_SM.N_162_0_cascade_ ;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_2 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_165_0_cascade_ ;
    wire \U712_REG_SM.C1_SYNCZ0Z_2 ;
    wire \U712_CHIP_RAM.CPU_TACK_6 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0 ;
    wire A_c_3;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_ ;
    wire A_c_10;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_a3_0 ;
    wire \U712_REG_SM.DS_EN_0_sqmuxa_1_cascade_ ;
    wire \U712_REG_SM.N_68 ;
    wire \U712_REG_SM.N_188_cascade_ ;
    wire \U712_REG_SM.N_162_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire ASn_c;
    wire REGSPACEn_c;
    wire \U712_REG_SM.DS_EN_0_sqmuxa_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire TSn_c;
    wire RAMENn_c;
    wire \U712_REG_SM.N_171_0 ;
    wire SIZ_c_0;
    wire \U712_REG_SM.LDS_OUT_2_0_0 ;
    wire \U712_REG_SM.UDS_OUT_2_0_0 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.N_33 ;
    wire CMA_c_1;
    wire CMA_c_2;
    wire A_c_4;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_ ;
    wire A_c_11;
    wire \U712_CHIP_RAM.N_34 ;
    wire A_c_7;
    wire A_c_14;
    wire A_c_15;
    wire A_c_8;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_6_cascade_ ;
    wire A_c_5;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_ ;
    wire A_c_12;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_REG_SM.N_167_0 ;
    wire \U712_REG_SM.N_117 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.RnW_m ;
    wire \U712_REG_SM.un1_LDS_OUT_0_sqmuxa_1_0 ;
    wire DBRn_c;
    wire U712_REG_SM_DBR_SYNC_0;
    wire U712_REG_SM_DBR_SYNC_1;
    wire SIZ_c_1;
    wire \U712_REG_SM.UDS_OUTZ0 ;
    wire U712_REG_SM_un1_UDSn_i;
    wire RESETn_c_i;
    wire A_c_9;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_ ;
    wire A_c_2;
    wire \U712_CHIP_RAM.N_32 ;
    wire \U712_CHIP_RAM.N_37 ;
    wire CMA_c_5;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_5 ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.N_35 ;
    wire CMA_c_3;
    wire A_c_6;
    wire A_c_13;
    wire \U712_CHIP_RAM.N_36_cascade_ ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_ns_1_2 ;
    wire \U712_CHIP_RAM.N_61_cascade_ ;
    wire \U712_CHIP_RAM.N_65_cascade_ ;
    wire \U712_CHIP_RAM.N_104_1 ;
    wire \U712_CHIP_RAM.N_51 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER16_2_0_cascade_ ;
    wire \U712_CHIP_RAM.N_99_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_cascade_ ;
    wire \U712_CHIP_RAM.N_67_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER18_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_m2_3_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_7 ;
    wire \U712_BYTE_ENABLE.un2_CUMBEnZ0_cascade_ ;
    wire CUMBEn_c;
    wire \U712_BYTE_ENABLE.LLBE_0_0_tz ;
    wire \U712_BYTE_ENABLE.un2_CLLBEnZ0_cascade_ ;
    wire CLLBEn_c;
    wire \U712_BYTE_ENABLE.un2_CLMBEnZ0_cascade_ ;
    wire CLMBEn_c;
    wire A_c_1;
    wire A_c_0;
    wire \U712_BYTE_ENABLE.LW_TRANS_0 ;
    wire \U712_BYTE_ENABLE.un2_CUUBEnZ0_cascade_ ;
    wire DBENn_c;
    wire CUUBEn_c;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ;
    wire bfn_14_4_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire A_c_17;
    wire \U712_CHIP_RAM.CMA_5_0_8_cascade_ ;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.N_38 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire A_c_19;
    wire CMA_c_9;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_4 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER18_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.N_158_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_ns_1_1 ;
    wire \U712_CHIP_RAM.N_132 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_i ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_5_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER18_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0 ;
    wire \U712_REG_SM.DS_ENZ0 ;
    wire \U712_REG_SM.LDS_OUTZ0 ;
    wire U712_REG_SM_un1_LDSn_i;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire CMA_c_7;
    wire A_c_18;
    wire A_c_16;
    wire \U712_CHIP_RAM.N_39 ;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_1_a3_0 ;
    wire \U712_CHIP_RAM.un1_CMA31_0_i ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6 ;
    wire \U712_REG_SM.N_173_0 ;
    wire \U712_REG_SM.N_183_1 ;
    wire \U712_REG_SM.N_165_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.un1_DBR_SYNC ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_2_1 ;
    wire \U712_CHIP_RAM.N_108 ;
    wire \U712_CHIP_RAM.N_77_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4 ;
    wire \U712_CHIP_RAM.N_80 ;
    wire \U712_CHIP_RAM.N_77 ;
    wire \U712_CHIP_RAM.N_80_cascade_ ;
    wire \U712_CHIP_RAM.N_50_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.N_60 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER39_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER39_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_50 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire CASLn_c;
    wire CASUn_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire DBDIR_c;
    wire DRDDIR_0_i;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.un1_CMA31_0_i_0 ;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.N_65 ;
    wire \U712_CHIP_RAM.N_78 ;
    wire \U712_CHIP_RAM.N_67 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_cascade_ ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_5 ;
    wire \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.REFRESH_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_135 ;
    wire \U712_CHIP_RAM.N_122 ;
    wire \U712_CHIP_RAM.N_135_cascade_ ;
    wire \U712_CHIP_RAM.N_121 ;
    wire \U712_CHIP_RAM.N_66 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_2_cascade_ ;
    wire \U712_CHIP_RAM.N_61 ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire RnW_c;
    wire CPU_CYCLEm;
    wire AWEn_c;
    wire \U712_CHIP_RAM.N_47 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_63 ;
    wire RESETn_c;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_63_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER46 ;
    wire \U712_CHIP_RAM.N_127 ;
    wire \U712_CHIP_RAM.N_124 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.N_107 ;
    wire REG_CYCLEm;
    wire DMA_CYCLEm;
    wire DRDENn_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire WEn_c;
    wire RAS0n_c;
    wire RAS1n_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire CLK80_OUT;
    wire RESETn_c_i_g;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_OUT_i),
            .REFERENCECLK(N__3610),
            .RESETB(N__9217),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_OUT),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__10331),
            .DIN(N__10330),
            .DOUT(N__10329),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__10331),
            .PADOUT(N__10330),
            .PADIN(N__10329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5788),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__10322),
            .DIN(N__10321),
            .DOUT(N__10320),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__10322),
            .PADOUT(N__10321),
            .PADIN(N__10320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__10313),
            .DIN(N__10312),
            .DOUT(N__10311),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__10313),
            .PADOUT(N__10312),
            .PADIN(N__10311),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8566),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__10304),
            .DIN(N__10303),
            .DOUT(N__10302),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__10304),
            .PADOUT(N__10303),
            .PADIN(N__10302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7435),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__10295),
            .DIN(N__10294),
            .DOUT(N__10293),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__10295),
            .PADOUT(N__10294),
            .PADIN(N__10293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKEN_obuf_iopad (
            .OE(N__10286),
            .DIN(N__10285),
            .DOUT(N__10284),
            .PACKAGEPIN(CLKEN));
    defparam CLKEN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKEN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKEN_obuf_preio (
            .PADOEN(N__10286),
            .PADOUT(N__10285),
            .PADIN(N__10284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9213),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__10277),
            .DIN(N__10276),
            .DOUT(N__10275),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__10277),
            .PADOUT(N__10276),
            .PADIN(N__10275),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__10268),
            .DIN(N__10267),
            .DOUT(N__10266),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__10268),
            .PADOUT(N__10267),
            .PADIN(N__10266),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__10259),
            .DIN(N__10258),
            .DOUT(N__10257),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__10259),
            .PADOUT(N__10258),
            .PADIN(N__10257),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__10250),
            .DIN(N__10249),
            .DOUT(N__10248),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__10250),
            .PADOUT(N__10249),
            .PADIN(N__10248),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__10241),
            .DIN(N__10240),
            .DOUT(N__10239),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__10241),
            .PADOUT(N__10240),
            .PADIN(N__10239),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__10232),
            .DIN(N__10231),
            .DOUT(N__10230),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__10232),
            .PADOUT(N__10231),
            .PADIN(N__10230),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6205),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__10223),
            .DIN(N__10222),
            .DOUT(N__10221),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__10223),
            .PADOUT(N__10222),
            .PADIN(N__10221),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4290),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__10214),
            .DIN(N__10213),
            .DOUT(N__10212),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__10214),
            .PADOUT(N__10213),
            .PADIN(N__10212),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__10205),
            .DIN(N__10204),
            .DOUT(N__10203),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__10205),
            .PADOUT(N__10204),
            .PADIN(N__10203),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__10196),
            .DIN(N__10195),
            .DOUT(N__10194),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__10196),
            .PADOUT(N__10195),
            .PADIN(N__10194),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3799),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__10187),
            .DIN(N__10186),
            .DOUT(N__10185),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__10187),
            .PADOUT(N__10186),
            .PADIN(N__10185),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__10178),
            .DIN(N__10177),
            .DOUT(N__10176),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__10178),
            .PADOUT(N__10177),
            .PADIN(N__10176),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__10169),
            .DIN(N__10168),
            .DOUT(N__10167),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__10169),
            .PADOUT(N__10168),
            .PADIN(N__10167),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4615),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__10160),
            .DIN(N__10159),
            .DOUT(N__10158),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__10160),
            .PADOUT(N__10159),
            .PADIN(N__10158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__10151),
            .DIN(N__10150),
            .DOUT(N__10149),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__10151),
            .PADOUT(N__10150),
            .PADIN(N__10149),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8839),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__10142),
            .DIN(N__10141),
            .DOUT(N__10140),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__10142),
            .PADOUT(N__10141),
            .PADIN(N__10140),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__10133),
            .DIN(N__10132),
            .DOUT(N__10131),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__10133),
            .PADOUT(N__10132),
            .PADIN(N__10131),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__10124),
            .DIN(N__10123),
            .DOUT(N__10122),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__10124),
            .PADOUT(N__10123),
            .PADIN(N__10122),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__10115),
            .DIN(N__10114),
            .DOUT(N__10113),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__10115),
            .PADOUT(N__10114),
            .PADIN(N__10113),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__10106),
            .DIN(N__10105),
            .DOUT(N__10104),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__10106),
            .PADOUT(N__10105),
            .PADIN(N__10104),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__10097),
            .DIN(N__10096),
            .DOUT(N__10095),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__10097),
            .PADOUT(N__10096),
            .PADIN(N__10095),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__10088),
            .DIN(N__10087),
            .DOUT(N__10086),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__10088),
            .PADOUT(N__10087),
            .PADIN(N__10086),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__10079),
            .DIN(N__10078),
            .DOUT(N__10077),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__10079),
            .PADOUT(N__10078),
            .PADIN(N__10077),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__10070),
            .DIN(N__10069),
            .DOUT(N__10068),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__10070),
            .PADOUT(N__10069),
            .PADIN(N__10068),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__10061),
            .DIN(N__10060),
            .DOUT(N__10059),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__10061),
            .PADOUT(N__10060),
            .PADIN(N__10059),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__10052),
            .DIN(N__10051),
            .DOUT(N__10050),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__10052),
            .PADOUT(N__10051),
            .PADIN(N__10050),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5932),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__10043),
            .DIN(N__10042),
            .DOUT(N__10041),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__10043),
            .PADOUT(N__10042),
            .PADIN(N__10041),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__10034),
            .DIN(N__10033),
            .DOUT(N__10032),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__10034),
            .PADOUT(N__10033),
            .PADIN(N__10032),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__10025),
            .DIN(N__10024),
            .DOUT(N__10023),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__10025),
            .PADOUT(N__10024),
            .PADIN(N__10023),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__10016),
            .DIN(N__10015),
            .DOUT(N__10014),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__10016),
            .PADOUT(N__10015),
            .PADIN(N__10014),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__10007),
            .DIN(N__10006),
            .DOUT(N__10005),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__10007),
            .PADOUT(N__10006),
            .PADIN(N__10005),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3685),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__9998),
            .DIN(N__9997),
            .DOUT(N__9996),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__9998),
            .PADOUT(N__9997),
            .PADIN(N__9996),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6271),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__9989),
            .DIN(N__9988),
            .DOUT(N__9987),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__9989),
            .PADOUT(N__9988),
            .PADIN(N__9987),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__9980),
            .DIN(N__9979),
            .DOUT(N__9978),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__9980),
            .PADOUT(N__9979),
            .PADIN(N__9978),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8722),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__9971),
            .DIN(N__9970),
            .DOUT(N__9969),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__9971),
            .PADOUT(N__9970),
            .PADIN(N__9969),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__9962),
            .DIN(N__9961),
            .DOUT(N__9960),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__9962),
            .PADOUT(N__9961),
            .PADIN(N__9960),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__9953),
            .DIN(N__9952),
            .DOUT(N__9951),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__9953),
            .PADOUT(N__9952),
            .PADIN(N__9951),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3625),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__9944),
            .DIN(N__9943),
            .DOUT(N__9942),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__9944),
            .PADOUT(N__9943),
            .PADIN(N__9942),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__9935),
            .DIN(N__9934),
            .DOUT(N__9933),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__9935),
            .PADOUT(N__9934),
            .PADIN(N__9933),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4429),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__9926),
            .DIN(N__9925),
            .DOUT(N__9924),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__9926),
            .PADOUT(N__9925),
            .PADIN(N__9924),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5368),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__9917),
            .DIN(N__9916),
            .DOUT(N__9915),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__9917),
            .PADOUT(N__9916),
            .PADIN(N__9915),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__9908),
            .DIN(N__9907),
            .DOUT(N__9906),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__9908),
            .PADOUT(N__9907),
            .PADIN(N__9906),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_0_iopad (
            .OE(N__9899),
            .DIN(N__9898),
            .DOUT(N__9897),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__9899),
            .PADOUT(N__9898),
            .PADIN(N__9897),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__9890),
            .DIN(N__9889),
            .DOUT(N__9888),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__9890),
            .PADOUT(N__9889),
            .PADIN(N__9888),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7414),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__9881),
            .DIN(N__9880),
            .DOUT(N__9879),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__9881),
            .PADOUT(N__9880),
            .PADIN(N__9879),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__9872),
            .DIN(N__9871),
            .DOUT(N__9870),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__9872),
            .PADOUT(N__9871),
            .PADIN(N__9870),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5302),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__9863),
            .DIN(N__9862),
            .DOUT(N__9861),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__9863),
            .PADOUT(N__9862),
            .PADIN(N__9861),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9085),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__9854),
            .DIN(N__9853),
            .DOUT(N__9852),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__9854),
            .PADOUT(N__9853),
            .PADIN(N__9852),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5554),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__9845),
            .DIN(N__9844),
            .DOUT(N__9843),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__9845),
            .PADOUT(N__9844),
            .PADIN(N__9843),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5881),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__9836),
            .DIN(N__9835),
            .DOUT(N__9834),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__9836),
            .PADOUT(N__9835),
            .PADIN(N__9834),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4428),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__9827),
            .DIN(N__9826),
            .DOUT(N__9825),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__9827),
            .PADOUT(N__9826),
            .PADIN(N__9825),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__9818),
            .DIN(N__9817),
            .DOUT(N__9816),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__9818),
            .PADOUT(N__9817),
            .PADIN(N__9816),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__9809),
            .DIN(N__9808),
            .DOUT(N__9807),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__9809),
            .PADOUT(N__9808),
            .PADIN(N__9807),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5530),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__9800),
            .DIN(N__9799),
            .DOUT(N__9798),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__9800),
            .PADOUT(N__9799),
            .PADIN(N__9798),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8431),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__9791),
            .DIN(N__9790),
            .DOUT(N__9789),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__9791),
            .PADOUT(N__9790),
            .PADIN(N__9789),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7477),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__9782),
            .DIN(N__9781),
            .DOUT(N__9780),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__9782),
            .PADOUT(N__9781),
            .PADIN(N__9780),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5590),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__9773),
            .DIN(N__9772),
            .DOUT(N__9771),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__9773),
            .PADOUT(N__9772),
            .PADIN(N__9771),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__9764),
            .DIN(N__9763),
            .DOUT(N__9762),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__9764),
            .PADOUT(N__9763),
            .PADIN(N__9762),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__9755),
            .DIN(N__9754),
            .DOUT(N__9753),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__9755),
            .PADOUT(N__9754),
            .PADIN(N__9753),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__9746),
            .DIN(N__9745),
            .DOUT(N__9744),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__9746),
            .PADOUT(N__9745),
            .PADIN(N__9744),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__9737),
            .DIN(N__9736),
            .DOUT(N__9735),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__9737),
            .PADOUT(N__9736),
            .PADIN(N__9735),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4594),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__9728),
            .DIN(N__9727),
            .DOUT(N__9726),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__9728),
            .PADOUT(N__9727),
            .PADIN(N__9726),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__9719),
            .DIN(N__9718),
            .DOUT(N__9717),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__9719),
            .PADOUT(N__9718),
            .PADIN(N__9717),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5746),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__9710),
            .DIN(N__9709),
            .DOUT(N__9708),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__9710),
            .PADOUT(N__9709),
            .PADIN(N__9708),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3649),
            .DIN0(),
            .DOUT0(N__3736),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__9701),
            .DIN(N__9700),
            .DOUT(N__9699),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__9701),
            .PADOUT(N__9700),
            .PADIN(N__9699),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4582),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__9692),
            .DIN(N__9691),
            .DOUT(N__9690),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__9692),
            .PADOUT(N__9691),
            .PADIN(N__9690),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__9683),
            .DIN(N__9682),
            .DOUT(N__9681),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__9683),
            .PADOUT(N__9682),
            .PADIN(N__9681),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__9674),
            .DIN(N__9673),
            .DOUT(N__9672),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__9674),
            .PADOUT(N__9673),
            .PADIN(N__9672),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5962),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__9665),
            .DIN(N__9664),
            .DOUT(N__9663),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__9665),
            .PADOUT(N__9664),
            .PADIN(N__9663),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__9656),
            .DIN(N__9655),
            .DOUT(N__9654),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__9656),
            .PADOUT(N__9655),
            .PADIN(N__9654),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__9647),
            .DIN(N__9646),
            .DOUT(N__9645),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__9647),
            .PADOUT(N__9646),
            .PADIN(N__9645),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__9638),
            .DIN(N__9637),
            .DOUT(N__9636),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__9638),
            .PADOUT(N__9637),
            .PADIN(N__9636),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__9629),
            .DIN(N__9628),
            .DOUT(N__9627),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__9629),
            .PADOUT(N__9628),
            .PADIN(N__9627),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5206),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__9620),
            .DIN(N__9619),
            .DOUT(N__9618),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__9620),
            .PADOUT(N__9619),
            .PADIN(N__9618),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4852),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2307 (
            .O(N__9601),
            .I(N__9598));
    LocalMux I__2306 (
            .O(N__9598),
            .I(N__9595));
    Odrv12 I__2305 (
            .O(N__9595),
            .I(RAS1n_c));
    InMux I__2304 (
            .O(N__9592),
            .I(N__9588));
    InMux I__2303 (
            .O(N__9591),
            .I(N__9585));
    LocalMux I__2302 (
            .O(N__9588),
            .I(N__9582));
    LocalMux I__2301 (
            .O(N__9585),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    Odrv4 I__2300 (
            .O(N__9582),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2299 (
            .O(N__9577),
            .I(N__9574));
    LocalMux I__2298 (
            .O(N__9574),
            .I(N__9535));
    ClkMux I__2297 (
            .O(N__9573),
            .I(N__9421));
    ClkMux I__2296 (
            .O(N__9572),
            .I(N__9421));
    ClkMux I__2295 (
            .O(N__9571),
            .I(N__9421));
    ClkMux I__2294 (
            .O(N__9570),
            .I(N__9421));
    ClkMux I__2293 (
            .O(N__9569),
            .I(N__9421));
    ClkMux I__2292 (
            .O(N__9568),
            .I(N__9421));
    ClkMux I__2291 (
            .O(N__9567),
            .I(N__9421));
    ClkMux I__2290 (
            .O(N__9566),
            .I(N__9421));
    ClkMux I__2289 (
            .O(N__9565),
            .I(N__9421));
    ClkMux I__2288 (
            .O(N__9564),
            .I(N__9421));
    ClkMux I__2287 (
            .O(N__9563),
            .I(N__9421));
    ClkMux I__2286 (
            .O(N__9562),
            .I(N__9421));
    ClkMux I__2285 (
            .O(N__9561),
            .I(N__9421));
    ClkMux I__2284 (
            .O(N__9560),
            .I(N__9421));
    ClkMux I__2283 (
            .O(N__9559),
            .I(N__9421));
    ClkMux I__2282 (
            .O(N__9558),
            .I(N__9421));
    ClkMux I__2281 (
            .O(N__9557),
            .I(N__9421));
    ClkMux I__2280 (
            .O(N__9556),
            .I(N__9421));
    ClkMux I__2279 (
            .O(N__9555),
            .I(N__9421));
    ClkMux I__2278 (
            .O(N__9554),
            .I(N__9421));
    ClkMux I__2277 (
            .O(N__9553),
            .I(N__9421));
    ClkMux I__2276 (
            .O(N__9552),
            .I(N__9421));
    ClkMux I__2275 (
            .O(N__9551),
            .I(N__9421));
    ClkMux I__2274 (
            .O(N__9550),
            .I(N__9421));
    ClkMux I__2273 (
            .O(N__9549),
            .I(N__9421));
    ClkMux I__2272 (
            .O(N__9548),
            .I(N__9421));
    ClkMux I__2271 (
            .O(N__9547),
            .I(N__9421));
    ClkMux I__2270 (
            .O(N__9546),
            .I(N__9421));
    ClkMux I__2269 (
            .O(N__9545),
            .I(N__9421));
    ClkMux I__2268 (
            .O(N__9544),
            .I(N__9421));
    ClkMux I__2267 (
            .O(N__9543),
            .I(N__9421));
    ClkMux I__2266 (
            .O(N__9542),
            .I(N__9421));
    ClkMux I__2265 (
            .O(N__9541),
            .I(N__9421));
    ClkMux I__2264 (
            .O(N__9540),
            .I(N__9421));
    ClkMux I__2263 (
            .O(N__9539),
            .I(N__9421));
    ClkMux I__2262 (
            .O(N__9538),
            .I(N__9421));
    Glb2LocalMux I__2261 (
            .O(N__9535),
            .I(N__9421));
    ClkMux I__2260 (
            .O(N__9534),
            .I(N__9421));
    ClkMux I__2259 (
            .O(N__9533),
            .I(N__9421));
    ClkMux I__2258 (
            .O(N__9532),
            .I(N__9421));
    ClkMux I__2257 (
            .O(N__9531),
            .I(N__9421));
    ClkMux I__2256 (
            .O(N__9530),
            .I(N__9421));
    ClkMux I__2255 (
            .O(N__9529),
            .I(N__9421));
    ClkMux I__2254 (
            .O(N__9528),
            .I(N__9421));
    ClkMux I__2253 (
            .O(N__9527),
            .I(N__9421));
    ClkMux I__2252 (
            .O(N__9526),
            .I(N__9421));
    ClkMux I__2251 (
            .O(N__9525),
            .I(N__9421));
    ClkMux I__2250 (
            .O(N__9524),
            .I(N__9421));
    ClkMux I__2249 (
            .O(N__9523),
            .I(N__9421));
    ClkMux I__2248 (
            .O(N__9522),
            .I(N__9421));
    GlobalMux I__2247 (
            .O(N__9421),
            .I(CLK80_OUT));
    InMux I__2246 (
            .O(N__9418),
            .I(N__9406));
    InMux I__2245 (
            .O(N__9417),
            .I(N__9403));
    InMux I__2244 (
            .O(N__9416),
            .I(N__9400));
    InMux I__2243 (
            .O(N__9415),
            .I(N__9391));
    InMux I__2242 (
            .O(N__9414),
            .I(N__9391));
    InMux I__2241 (
            .O(N__9413),
            .I(N__9391));
    InMux I__2240 (
            .O(N__9412),
            .I(N__9391));
    InMux I__2239 (
            .O(N__9411),
            .I(N__9388));
    InMux I__2238 (
            .O(N__9410),
            .I(N__9385));
    InMux I__2237 (
            .O(N__9409),
            .I(N__9382));
    LocalMux I__2236 (
            .O(N__9406),
            .I(N__9371));
    LocalMux I__2235 (
            .O(N__9403),
            .I(N__9360));
    LocalMux I__2234 (
            .O(N__9400),
            .I(N__9346));
    LocalMux I__2233 (
            .O(N__9391),
            .I(N__9341));
    LocalMux I__2232 (
            .O(N__9388),
            .I(N__9335));
    LocalMux I__2231 (
            .O(N__9385),
            .I(N__9332));
    LocalMux I__2230 (
            .O(N__9382),
            .I(N__9325));
    SRMux I__2229 (
            .O(N__9381),
            .I(N__9223));
    SRMux I__2228 (
            .O(N__9380),
            .I(N__9223));
    SRMux I__2227 (
            .O(N__9379),
            .I(N__9223));
    SRMux I__2226 (
            .O(N__9378),
            .I(N__9223));
    SRMux I__2225 (
            .O(N__9377),
            .I(N__9223));
    SRMux I__2224 (
            .O(N__9376),
            .I(N__9223));
    SRMux I__2223 (
            .O(N__9375),
            .I(N__9223));
    SRMux I__2222 (
            .O(N__9374),
            .I(N__9223));
    Glb2LocalMux I__2221 (
            .O(N__9371),
            .I(N__9223));
    SRMux I__2220 (
            .O(N__9370),
            .I(N__9223));
    SRMux I__2219 (
            .O(N__9369),
            .I(N__9223));
    SRMux I__2218 (
            .O(N__9368),
            .I(N__9223));
    SRMux I__2217 (
            .O(N__9367),
            .I(N__9223));
    SRMux I__2216 (
            .O(N__9366),
            .I(N__9223));
    SRMux I__2215 (
            .O(N__9365),
            .I(N__9223));
    SRMux I__2214 (
            .O(N__9364),
            .I(N__9223));
    SRMux I__2213 (
            .O(N__9363),
            .I(N__9223));
    Glb2LocalMux I__2212 (
            .O(N__9360),
            .I(N__9223));
    SRMux I__2211 (
            .O(N__9359),
            .I(N__9223));
    SRMux I__2210 (
            .O(N__9358),
            .I(N__9223));
    SRMux I__2209 (
            .O(N__9357),
            .I(N__9223));
    SRMux I__2208 (
            .O(N__9356),
            .I(N__9223));
    SRMux I__2207 (
            .O(N__9355),
            .I(N__9223));
    SRMux I__2206 (
            .O(N__9354),
            .I(N__9223));
    SRMux I__2205 (
            .O(N__9353),
            .I(N__9223));
    SRMux I__2204 (
            .O(N__9352),
            .I(N__9223));
    SRMux I__2203 (
            .O(N__9351),
            .I(N__9223));
    SRMux I__2202 (
            .O(N__9350),
            .I(N__9223));
    SRMux I__2201 (
            .O(N__9349),
            .I(N__9223));
    Glb2LocalMux I__2200 (
            .O(N__9346),
            .I(N__9223));
    SRMux I__2199 (
            .O(N__9345),
            .I(N__9223));
    SRMux I__2198 (
            .O(N__9344),
            .I(N__9223));
    Glb2LocalMux I__2197 (
            .O(N__9341),
            .I(N__9223));
    SRMux I__2196 (
            .O(N__9340),
            .I(N__9223));
    SRMux I__2195 (
            .O(N__9339),
            .I(N__9223));
    SRMux I__2194 (
            .O(N__9338),
            .I(N__9223));
    Glb2LocalMux I__2193 (
            .O(N__9335),
            .I(N__9223));
    Glb2LocalMux I__2192 (
            .O(N__9332),
            .I(N__9223));
    SRMux I__2191 (
            .O(N__9331),
            .I(N__9223));
    SRMux I__2190 (
            .O(N__9330),
            .I(N__9223));
    SRMux I__2189 (
            .O(N__9329),
            .I(N__9223));
    SRMux I__2188 (
            .O(N__9328),
            .I(N__9223));
    Glb2LocalMux I__2187 (
            .O(N__9325),
            .I(N__9223));
    SRMux I__2186 (
            .O(N__9324),
            .I(N__9223));
    SRMux I__2185 (
            .O(N__9323),
            .I(N__9223));
    SRMux I__2184 (
            .O(N__9322),
            .I(N__9223));
    SRMux I__2183 (
            .O(N__9321),
            .I(N__9223));
    SRMux I__2182 (
            .O(N__9320),
            .I(N__9223));
    GlobalMux I__2181 (
            .O(N__9223),
            .I(N__9220));
    gio2CtrlBuf I__2180 (
            .O(N__9220),
            .I(RESETn_c_i_g));
    IoInMux I__2179 (
            .O(N__9217),
            .I(N__9214));
    LocalMux I__2178 (
            .O(N__9214),
            .I(N__9210));
    IoInMux I__2177 (
            .O(N__9213),
            .I(N__9207));
    Span4Mux_s3_v I__2176 (
            .O(N__9210),
            .I(N__9204));
    LocalMux I__2175 (
            .O(N__9207),
            .I(N__9201));
    Span4Mux_v I__2174 (
            .O(N__9204),
            .I(N__9198));
    Span4Mux_s3_h I__2173 (
            .O(N__9201),
            .I(N__9195));
    Span4Mux_h I__2172 (
            .O(N__9198),
            .I(N__9192));
    Span4Mux_h I__2171 (
            .O(N__9195),
            .I(N__9189));
    Odrv4 I__2170 (
            .O(N__9192),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2169 (
            .O(N__9189),
            .I(CONSTANT_ONE_NET));
    InMux I__2168 (
            .O(N__9184),
            .I(N__9181));
    LocalMux I__2167 (
            .O(N__9181),
            .I(N__9177));
    InMux I__2166 (
            .O(N__9180),
            .I(N__9174));
    Span4Mux_h I__2165 (
            .O(N__9177),
            .I(N__9168));
    LocalMux I__2164 (
            .O(N__9174),
            .I(N__9168));
    InMux I__2163 (
            .O(N__9173),
            .I(N__9165));
    Span4Mux_v I__2162 (
            .O(N__9168),
            .I(N__9162));
    LocalMux I__2161 (
            .O(N__9165),
            .I(N__9159));
    Sp12to4 I__2160 (
            .O(N__9162),
            .I(N__9155));
    Span4Mux_v I__2159 (
            .O(N__9159),
            .I(N__9152));
    InMux I__2158 (
            .O(N__9158),
            .I(N__9149));
    Odrv12 I__2157 (
            .O(N__9155),
            .I(REG_CYCLEm));
    Odrv4 I__2156 (
            .O(N__9152),
            .I(REG_CYCLEm));
    LocalMux I__2155 (
            .O(N__9149),
            .I(REG_CYCLEm));
    InMux I__2154 (
            .O(N__9142),
            .I(N__9136));
    InMux I__2153 (
            .O(N__9141),
            .I(N__9133));
    InMux I__2152 (
            .O(N__9140),
            .I(N__9130));
    InMux I__2151 (
            .O(N__9139),
            .I(N__9127));
    LocalMux I__2150 (
            .O(N__9136),
            .I(N__9119));
    LocalMux I__2149 (
            .O(N__9133),
            .I(N__9114));
    LocalMux I__2148 (
            .O(N__9130),
            .I(N__9114));
    LocalMux I__2147 (
            .O(N__9127),
            .I(N__9111));
    InMux I__2146 (
            .O(N__9126),
            .I(N__9102));
    InMux I__2145 (
            .O(N__9125),
            .I(N__9102));
    InMux I__2144 (
            .O(N__9124),
            .I(N__9102));
    InMux I__2143 (
            .O(N__9123),
            .I(N__9102));
    InMux I__2142 (
            .O(N__9122),
            .I(N__9099));
    Span4Mux_v I__2141 (
            .O(N__9119),
            .I(N__9094));
    Span4Mux_v I__2140 (
            .O(N__9114),
            .I(N__9094));
    Odrv4 I__2139 (
            .O(N__9111),
            .I(DMA_CYCLEm));
    LocalMux I__2138 (
            .O(N__9102),
            .I(DMA_CYCLEm));
    LocalMux I__2137 (
            .O(N__9099),
            .I(DMA_CYCLEm));
    Odrv4 I__2136 (
            .O(N__9094),
            .I(DMA_CYCLEm));
    IoInMux I__2135 (
            .O(N__9085),
            .I(N__9082));
    LocalMux I__2134 (
            .O(N__9082),
            .I(N__9079));
    IoSpan4Mux I__2133 (
            .O(N__9079),
            .I(N__9076));
    Sp12to4 I__2132 (
            .O(N__9076),
            .I(N__9073));
    Span12Mux_v I__2131 (
            .O(N__9073),
            .I(N__9070));
    Span12Mux_h I__2130 (
            .O(N__9070),
            .I(N__9067));
    Odrv12 I__2129 (
            .O(N__9067),
            .I(DRDENn_c));
    CEMux I__2128 (
            .O(N__9064),
            .I(N__9060));
    CEMux I__2127 (
            .O(N__9063),
            .I(N__9055));
    LocalMux I__2126 (
            .O(N__9060),
            .I(N__9052));
    CEMux I__2125 (
            .O(N__9059),
            .I(N__9049));
    CEMux I__2124 (
            .O(N__9058),
            .I(N__9046));
    LocalMux I__2123 (
            .O(N__9055),
            .I(N__9042));
    Span4Mux_h I__2122 (
            .O(N__9052),
            .I(N__9037));
    LocalMux I__2121 (
            .O(N__9049),
            .I(N__9037));
    LocalMux I__2120 (
            .O(N__9046),
            .I(N__9034));
    CEMux I__2119 (
            .O(N__9045),
            .I(N__9031));
    Span4Mux_v I__2118 (
            .O(N__9042),
            .I(N__9028));
    Span4Mux_v I__2117 (
            .O(N__9037),
            .I(N__9023));
    Span4Mux_v I__2116 (
            .O(N__9034),
            .I(N__9023));
    LocalMux I__2115 (
            .O(N__9031),
            .I(N__9020));
    Span4Mux_h I__2114 (
            .O(N__9028),
            .I(N__9017));
    Span4Mux_h I__2113 (
            .O(N__9023),
            .I(N__9012));
    Span4Mux_v I__2112 (
            .O(N__9020),
            .I(N__9012));
    Odrv4 I__2111 (
            .O(N__9017),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    Odrv4 I__2110 (
            .O(N__9012),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    InMux I__2109 (
            .O(N__9007),
            .I(N__9004));
    LocalMux I__2108 (
            .O(N__9004),
            .I(N__9000));
    InMux I__2107 (
            .O(N__9003),
            .I(N__8997));
    Span4Mux_v I__2106 (
            .O(N__9000),
            .I(N__8994));
    LocalMux I__2105 (
            .O(N__8997),
            .I(N__8991));
    Sp12to4 I__2104 (
            .O(N__8994),
            .I(N__8988));
    Span4Mux_h I__2103 (
            .O(N__8991),
            .I(N__8985));
    Span12Mux_h I__2102 (
            .O(N__8988),
            .I(N__8982));
    Sp12to4 I__2101 (
            .O(N__8985),
            .I(N__8979));
    Span12Mux_v I__2100 (
            .O(N__8982),
            .I(N__8976));
    Span12Mux_v I__2099 (
            .O(N__8979),
            .I(N__8973));
    Odrv12 I__2098 (
            .O(N__8976),
            .I(DRA_c_0));
    Odrv12 I__2097 (
            .O(N__8973),
            .I(DRA_c_0));
    CascadeMux I__2096 (
            .O(N__8968),
            .I(N__8965));
    InMux I__2095 (
            .O(N__8965),
            .I(N__8962));
    LocalMux I__2094 (
            .O(N__8962),
            .I(N__8959));
    Span12Mux_v I__2093 (
            .O(N__8959),
            .I(N__8956));
    Odrv12 I__2092 (
            .O(N__8956),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    CEMux I__2091 (
            .O(N__8953),
            .I(N__8949));
    CEMux I__2090 (
            .O(N__8952),
            .I(N__8946));
    LocalMux I__2089 (
            .O(N__8949),
            .I(N__8942));
    LocalMux I__2088 (
            .O(N__8946),
            .I(N__8939));
    CEMux I__2087 (
            .O(N__8945),
            .I(N__8936));
    Span4Mux_h I__2086 (
            .O(N__8942),
            .I(N__8927));
    Span4Mux_h I__2085 (
            .O(N__8939),
            .I(N__8927));
    LocalMux I__2084 (
            .O(N__8936),
            .I(N__8927));
    CEMux I__2083 (
            .O(N__8935),
            .I(N__8924));
    CEMux I__2082 (
            .O(N__8934),
            .I(N__8921));
    Span4Mux_v I__2081 (
            .O(N__8927),
            .I(N__8917));
    LocalMux I__2080 (
            .O(N__8924),
            .I(N__8914));
    LocalMux I__2079 (
            .O(N__8921),
            .I(N__8911));
    CEMux I__2078 (
            .O(N__8920),
            .I(N__8908));
    Span4Mux_h I__2077 (
            .O(N__8917),
            .I(N__8905));
    Span4Mux_h I__2076 (
            .O(N__8914),
            .I(N__8902));
    Span4Mux_h I__2075 (
            .O(N__8911),
            .I(N__8899));
    LocalMux I__2074 (
            .O(N__8908),
            .I(N__8896));
    Odrv4 I__2073 (
            .O(N__8905),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    Odrv4 I__2072 (
            .O(N__8902),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    Odrv4 I__2071 (
            .O(N__8899),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    Odrv12 I__2070 (
            .O(N__8896),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    InMux I__2069 (
            .O(N__8887),
            .I(N__8883));
    CascadeMux I__2068 (
            .O(N__8886),
            .I(N__8880));
    LocalMux I__2067 (
            .O(N__8883),
            .I(N__8876));
    InMux I__2066 (
            .O(N__8880),
            .I(N__8873));
    InMux I__2065 (
            .O(N__8879),
            .I(N__8870));
    Span4Mux_v I__2064 (
            .O(N__8876),
            .I(N__8867));
    LocalMux I__2063 (
            .O(N__8873),
            .I(N__8861));
    LocalMux I__2062 (
            .O(N__8870),
            .I(N__8861));
    Span4Mux_v I__2061 (
            .O(N__8867),
            .I(N__8858));
    InMux I__2060 (
            .O(N__8866),
            .I(N__8855));
    Span4Mux_h I__2059 (
            .O(N__8861),
            .I(N__8852));
    Span4Mux_h I__2058 (
            .O(N__8858),
            .I(N__8847));
    LocalMux I__2057 (
            .O(N__8855),
            .I(N__8847));
    Span4Mux_v I__2056 (
            .O(N__8852),
            .I(N__8844));
    Odrv4 I__2055 (
            .O(N__8847),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__2054 (
            .O(N__8844),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__2053 (
            .O(N__8839),
            .I(N__8836));
    LocalMux I__2052 (
            .O(N__8836),
            .I(N__8833));
    Span4Mux_s1_v I__2051 (
            .O(N__8833),
            .I(N__8830));
    Span4Mux_v I__2050 (
            .O(N__8830),
            .I(N__8827));
    Span4Mux_v I__2049 (
            .O(N__8827),
            .I(N__8824));
    Odrv4 I__2048 (
            .O(N__8824),
            .I(CRCSn_c));
    CascadeMux I__2047 (
            .O(N__8821),
            .I(N__8813));
    InMux I__2046 (
            .O(N__8820),
            .I(N__8808));
    InMux I__2045 (
            .O(N__8819),
            .I(N__8805));
    InMux I__2044 (
            .O(N__8818),
            .I(N__8802));
    CascadeMux I__2043 (
            .O(N__8817),
            .I(N__8797));
    InMux I__2042 (
            .O(N__8816),
            .I(N__8794));
    InMux I__2041 (
            .O(N__8813),
            .I(N__8787));
    InMux I__2040 (
            .O(N__8812),
            .I(N__8787));
    InMux I__2039 (
            .O(N__8811),
            .I(N__8787));
    LocalMux I__2038 (
            .O(N__8808),
            .I(N__8782));
    LocalMux I__2037 (
            .O(N__8805),
            .I(N__8782));
    LocalMux I__2036 (
            .O(N__8802),
            .I(N__8778));
    InMux I__2035 (
            .O(N__8801),
            .I(N__8773));
    InMux I__2034 (
            .O(N__8800),
            .I(N__8773));
    InMux I__2033 (
            .O(N__8797),
            .I(N__8770));
    LocalMux I__2032 (
            .O(N__8794),
            .I(N__8761));
    LocalMux I__2031 (
            .O(N__8787),
            .I(N__8761));
    Span4Mux_h I__2030 (
            .O(N__8782),
            .I(N__8761));
    CascadeMux I__2029 (
            .O(N__8781),
            .I(N__8758));
    Span4Mux_v I__2028 (
            .O(N__8778),
            .I(N__8755));
    LocalMux I__2027 (
            .O(N__8773),
            .I(N__8750));
    LocalMux I__2026 (
            .O(N__8770),
            .I(N__8750));
    InMux I__2025 (
            .O(N__8769),
            .I(N__8747));
    InMux I__2024 (
            .O(N__8768),
            .I(N__8744));
    Span4Mux_v I__2023 (
            .O(N__8761),
            .I(N__8741));
    InMux I__2022 (
            .O(N__8758),
            .I(N__8738));
    Span4Mux_h I__2021 (
            .O(N__8755),
            .I(N__8733));
    Span4Mux_v I__2020 (
            .O(N__8750),
            .I(N__8733));
    LocalMux I__2019 (
            .O(N__8747),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__2018 (
            .O(N__8744),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2017 (
            .O(N__8741),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__2016 (
            .O(N__8738),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2015 (
            .O(N__8733),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__2014 (
            .O(N__8722),
            .I(N__8719));
    LocalMux I__2013 (
            .O(N__8719),
            .I(N__8716));
    Span4Mux_s2_v I__2012 (
            .O(N__8716),
            .I(N__8713));
    Span4Mux_v I__2011 (
            .O(N__8713),
            .I(N__8710));
    Span4Mux_v I__2010 (
            .O(N__8710),
            .I(N__8707));
    Odrv4 I__2009 (
            .O(N__8707),
            .I(RASn_c));
    InMux I__2008 (
            .O(N__8704),
            .I(N__8696));
    CascadeMux I__2007 (
            .O(N__8703),
            .I(N__8692));
    CascadeMux I__2006 (
            .O(N__8702),
            .I(N__8687));
    InMux I__2005 (
            .O(N__8701),
            .I(N__8684));
    CascadeMux I__2004 (
            .O(N__8700),
            .I(N__8681));
    CascadeMux I__2003 (
            .O(N__8699),
            .I(N__8677));
    LocalMux I__2002 (
            .O(N__8696),
            .I(N__8673));
    InMux I__2001 (
            .O(N__8695),
            .I(N__8670));
    InMux I__2000 (
            .O(N__8692),
            .I(N__8667));
    InMux I__1999 (
            .O(N__8691),
            .I(N__8664));
    InMux I__1998 (
            .O(N__8690),
            .I(N__8660));
    InMux I__1997 (
            .O(N__8687),
            .I(N__8657));
    LocalMux I__1996 (
            .O(N__8684),
            .I(N__8654));
    InMux I__1995 (
            .O(N__8681),
            .I(N__8651));
    InMux I__1994 (
            .O(N__8680),
            .I(N__8648));
    InMux I__1993 (
            .O(N__8677),
            .I(N__8645));
    InMux I__1992 (
            .O(N__8676),
            .I(N__8641));
    Span4Mux_v I__1991 (
            .O(N__8673),
            .I(N__8638));
    LocalMux I__1990 (
            .O(N__8670),
            .I(N__8633));
    LocalMux I__1989 (
            .O(N__8667),
            .I(N__8633));
    LocalMux I__1988 (
            .O(N__8664),
            .I(N__8630));
    InMux I__1987 (
            .O(N__8663),
            .I(N__8627));
    LocalMux I__1986 (
            .O(N__8660),
            .I(N__8622));
    LocalMux I__1985 (
            .O(N__8657),
            .I(N__8622));
    Span4Mux_v I__1984 (
            .O(N__8654),
            .I(N__8617));
    LocalMux I__1983 (
            .O(N__8651),
            .I(N__8617));
    LocalMux I__1982 (
            .O(N__8648),
            .I(N__8612));
    LocalMux I__1981 (
            .O(N__8645),
            .I(N__8609));
    InMux I__1980 (
            .O(N__8644),
            .I(N__8606));
    LocalMux I__1979 (
            .O(N__8641),
            .I(N__8603));
    Span4Mux_v I__1978 (
            .O(N__8638),
            .I(N__8598));
    Span4Mux_v I__1977 (
            .O(N__8633),
            .I(N__8598));
    Span4Mux_h I__1976 (
            .O(N__8630),
            .I(N__8589));
    LocalMux I__1975 (
            .O(N__8627),
            .I(N__8589));
    Span4Mux_h I__1974 (
            .O(N__8622),
            .I(N__8589));
    Span4Mux_h I__1973 (
            .O(N__8617),
            .I(N__8589));
    InMux I__1972 (
            .O(N__8616),
            .I(N__8584));
    InMux I__1971 (
            .O(N__8615),
            .I(N__8584));
    Span4Mux_v I__1970 (
            .O(N__8612),
            .I(N__8575));
    Span4Mux_h I__1969 (
            .O(N__8609),
            .I(N__8575));
    LocalMux I__1968 (
            .O(N__8606),
            .I(N__8575));
    Span4Mux_v I__1967 (
            .O(N__8603),
            .I(N__8575));
    Odrv4 I__1966 (
            .O(N__8598),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1965 (
            .O(N__8589),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1964 (
            .O(N__8584),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1963 (
            .O(N__8575),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    IoInMux I__1962 (
            .O(N__8566),
            .I(N__8563));
    LocalMux I__1961 (
            .O(N__8563),
            .I(N__8560));
    Span4Mux_s3_v I__1960 (
            .O(N__8560),
            .I(N__8557));
    Sp12to4 I__1959 (
            .O(N__8557),
            .I(N__8554));
    Span12Mux_s10_h I__1958 (
            .O(N__8554),
            .I(N__8551));
    Odrv12 I__1957 (
            .O(N__8551),
            .I(CASn_c));
    InMux I__1956 (
            .O(N__8548),
            .I(N__8545));
    LocalMux I__1955 (
            .O(N__8545),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    InMux I__1954 (
            .O(N__8542),
            .I(N__8535));
    CascadeMux I__1953 (
            .O(N__8541),
            .I(N__8531));
    CascadeMux I__1952 (
            .O(N__8540),
            .I(N__8527));
    CascadeMux I__1951 (
            .O(N__8539),
            .I(N__8524));
    InMux I__1950 (
            .O(N__8538),
            .I(N__8521));
    LocalMux I__1949 (
            .O(N__8535),
            .I(N__8518));
    InMux I__1948 (
            .O(N__8534),
            .I(N__8512));
    InMux I__1947 (
            .O(N__8531),
            .I(N__8507));
    InMux I__1946 (
            .O(N__8530),
            .I(N__8500));
    InMux I__1945 (
            .O(N__8527),
            .I(N__8500));
    InMux I__1944 (
            .O(N__8524),
            .I(N__8500));
    LocalMux I__1943 (
            .O(N__8521),
            .I(N__8497));
    Span4Mux_h I__1942 (
            .O(N__8518),
            .I(N__8494));
    InMux I__1941 (
            .O(N__8517),
            .I(N__8489));
    InMux I__1940 (
            .O(N__8516),
            .I(N__8489));
    InMux I__1939 (
            .O(N__8515),
            .I(N__8486));
    LocalMux I__1938 (
            .O(N__8512),
            .I(N__8483));
    InMux I__1937 (
            .O(N__8511),
            .I(N__8480));
    InMux I__1936 (
            .O(N__8510),
            .I(N__8477));
    LocalMux I__1935 (
            .O(N__8507),
            .I(N__8472));
    LocalMux I__1934 (
            .O(N__8500),
            .I(N__8472));
    Span4Mux_v I__1933 (
            .O(N__8497),
            .I(N__8469));
    Span4Mux_h I__1932 (
            .O(N__8494),
            .I(N__8460));
    LocalMux I__1931 (
            .O(N__8489),
            .I(N__8460));
    LocalMux I__1930 (
            .O(N__8486),
            .I(N__8460));
    Span4Mux_v I__1929 (
            .O(N__8483),
            .I(N__8457));
    LocalMux I__1928 (
            .O(N__8480),
            .I(N__8448));
    LocalMux I__1927 (
            .O(N__8477),
            .I(N__8448));
    Span4Mux_v I__1926 (
            .O(N__8472),
            .I(N__8448));
    Span4Mux_v I__1925 (
            .O(N__8469),
            .I(N__8448));
    InMux I__1924 (
            .O(N__8468),
            .I(N__8443));
    InMux I__1923 (
            .O(N__8467),
            .I(N__8443));
    Span4Mux_v I__1922 (
            .O(N__8460),
            .I(N__8440));
    Odrv4 I__1921 (
            .O(N__8457),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1920 (
            .O(N__8448),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1919 (
            .O(N__8443),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1918 (
            .O(N__8440),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1917 (
            .O(N__8431),
            .I(N__8428));
    LocalMux I__1916 (
            .O(N__8428),
            .I(N__8425));
    IoSpan4Mux I__1915 (
            .O(N__8425),
            .I(N__8422));
    Span4Mux_s1_h I__1914 (
            .O(N__8422),
            .I(N__8419));
    Span4Mux_v I__1913 (
            .O(N__8419),
            .I(N__8416));
    Span4Mux_v I__1912 (
            .O(N__8416),
            .I(N__8413));
    Span4Mux_h I__1911 (
            .O(N__8413),
            .I(N__8410));
    Odrv4 I__1910 (
            .O(N__8410),
            .I(WEn_c));
    InMux I__1909 (
            .O(N__8407),
            .I(N__8404));
    LocalMux I__1908 (
            .O(N__8404),
            .I(N__8400));
    InMux I__1907 (
            .O(N__8403),
            .I(N__8397));
    Span4Mux_v I__1906 (
            .O(N__8400),
            .I(N__8394));
    LocalMux I__1905 (
            .O(N__8397),
            .I(N__8391));
    Span4Mux_h I__1904 (
            .O(N__8394),
            .I(N__8388));
    Sp12to4 I__1903 (
            .O(N__8391),
            .I(N__8385));
    Sp12to4 I__1902 (
            .O(N__8388),
            .I(N__8380));
    Span12Mux_v I__1901 (
            .O(N__8385),
            .I(N__8380));
    Odrv12 I__1900 (
            .O(N__8380),
            .I(RAS0n_c));
    InMux I__1899 (
            .O(N__8377),
            .I(N__8373));
    InMux I__1898 (
            .O(N__8376),
            .I(N__8370));
    LocalMux I__1897 (
            .O(N__8373),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ));
    LocalMux I__1896 (
            .O(N__8370),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ));
    InMux I__1895 (
            .O(N__8365),
            .I(N__8358));
    InMux I__1894 (
            .O(N__8364),
            .I(N__8358));
    InMux I__1893 (
            .O(N__8363),
            .I(N__8355));
    LocalMux I__1892 (
            .O(N__8358),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    LocalMux I__1891 (
            .O(N__8355),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    InMux I__1890 (
            .O(N__8350),
            .I(N__8345));
    InMux I__1889 (
            .O(N__8349),
            .I(N__8342));
    InMux I__1888 (
            .O(N__8348),
            .I(N__8339));
    LocalMux I__1887 (
            .O(N__8345),
            .I(N__8336));
    LocalMux I__1886 (
            .O(N__8342),
            .I(N__8333));
    LocalMux I__1885 (
            .O(N__8339),
            .I(N__8328));
    Span4Mux_v I__1884 (
            .O(N__8336),
            .I(N__8328));
    Odrv12 I__1883 (
            .O(N__8333),
            .I(\U712_CHIP_RAM.N_135 ));
    Odrv4 I__1882 (
            .O(N__8328),
            .I(\U712_CHIP_RAM.N_135 ));
    InMux I__1881 (
            .O(N__8323),
            .I(N__8317));
    InMux I__1880 (
            .O(N__8322),
            .I(N__8314));
    InMux I__1879 (
            .O(N__8321),
            .I(N__8309));
    InMux I__1878 (
            .O(N__8320),
            .I(N__8309));
    LocalMux I__1877 (
            .O(N__8317),
            .I(\U712_CHIP_RAM.N_122 ));
    LocalMux I__1876 (
            .O(N__8314),
            .I(\U712_CHIP_RAM.N_122 ));
    LocalMux I__1875 (
            .O(N__8309),
            .I(\U712_CHIP_RAM.N_122 ));
    CascadeMux I__1874 (
            .O(N__8302),
            .I(\U712_CHIP_RAM.N_135_cascade_ ));
    InMux I__1873 (
            .O(N__8299),
            .I(N__8294));
    InMux I__1872 (
            .O(N__8298),
            .I(N__8291));
    InMux I__1871 (
            .O(N__8297),
            .I(N__8288));
    LocalMux I__1870 (
            .O(N__8294),
            .I(\U712_CHIP_RAM.N_121 ));
    LocalMux I__1869 (
            .O(N__8291),
            .I(\U712_CHIP_RAM.N_121 ));
    LocalMux I__1868 (
            .O(N__8288),
            .I(\U712_CHIP_RAM.N_121 ));
    InMux I__1867 (
            .O(N__8281),
            .I(N__8278));
    LocalMux I__1866 (
            .O(N__8278),
            .I(\U712_CHIP_RAM.N_66 ));
    CascadeMux I__1865 (
            .O(N__8275),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_2_cascade_ ));
    CascadeMux I__1864 (
            .O(N__8272),
            .I(N__8268));
    InMux I__1863 (
            .O(N__8271),
            .I(N__8264));
    InMux I__1862 (
            .O(N__8268),
            .I(N__8261));
    InMux I__1861 (
            .O(N__8267),
            .I(N__8258));
    LocalMux I__1860 (
            .O(N__8264),
            .I(N__8255));
    LocalMux I__1859 (
            .O(N__8261),
            .I(N__8252));
    LocalMux I__1858 (
            .O(N__8258),
            .I(N__8245));
    Span4Mux_h I__1857 (
            .O(N__8255),
            .I(N__8240));
    Span4Mux_h I__1856 (
            .O(N__8252),
            .I(N__8240));
    InMux I__1855 (
            .O(N__8251),
            .I(N__8235));
    InMux I__1854 (
            .O(N__8250),
            .I(N__8235));
    InMux I__1853 (
            .O(N__8249),
            .I(N__8232));
    InMux I__1852 (
            .O(N__8248),
            .I(N__8229));
    Odrv4 I__1851 (
            .O(N__8245),
            .I(\U712_CHIP_RAM.N_61 ));
    Odrv4 I__1850 (
            .O(N__8240),
            .I(\U712_CHIP_RAM.N_61 ));
    LocalMux I__1849 (
            .O(N__8235),
            .I(\U712_CHIP_RAM.N_61 ));
    LocalMux I__1848 (
            .O(N__8232),
            .I(\U712_CHIP_RAM.N_61 ));
    LocalMux I__1847 (
            .O(N__8229),
            .I(\U712_CHIP_RAM.N_61 ));
    InMux I__1846 (
            .O(N__8218),
            .I(N__8215));
    LocalMux I__1845 (
            .O(N__8215),
            .I(N__8211));
    InMux I__1844 (
            .O(N__8214),
            .I(N__8208));
    Span4Mux_h I__1843 (
            .O(N__8211),
            .I(N__8205));
    LocalMux I__1842 (
            .O(N__8208),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__1841 (
            .O(N__8205),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    InMux I__1840 (
            .O(N__8200),
            .I(N__8196));
    InMux I__1839 (
            .O(N__8199),
            .I(N__8193));
    LocalMux I__1838 (
            .O(N__8196),
            .I(N__8190));
    LocalMux I__1837 (
            .O(N__8193),
            .I(N__8186));
    Span4Mux_v I__1836 (
            .O(N__8190),
            .I(N__8183));
    InMux I__1835 (
            .O(N__8189),
            .I(N__8180));
    Span4Mux_v I__1834 (
            .O(N__8186),
            .I(N__8175));
    Span4Mux_h I__1833 (
            .O(N__8183),
            .I(N__8170));
    LocalMux I__1832 (
            .O(N__8180),
            .I(N__8170));
    InMux I__1831 (
            .O(N__8179),
            .I(N__8167));
    CascadeMux I__1830 (
            .O(N__8178),
            .I(N__8164));
    Sp12to4 I__1829 (
            .O(N__8175),
            .I(N__8160));
    Span4Mux_h I__1828 (
            .O(N__8170),
            .I(N__8155));
    LocalMux I__1827 (
            .O(N__8167),
            .I(N__8155));
    InMux I__1826 (
            .O(N__8164),
            .I(N__8150));
    InMux I__1825 (
            .O(N__8163),
            .I(N__8150));
    Span12Mux_h I__1824 (
            .O(N__8160),
            .I(N__8147));
    Sp12to4 I__1823 (
            .O(N__8155),
            .I(N__8142));
    LocalMux I__1822 (
            .O(N__8150),
            .I(N__8142));
    Span12Mux_h I__1821 (
            .O(N__8147),
            .I(N__8139));
    Span12Mux_v I__1820 (
            .O(N__8142),
            .I(N__8136));
    Span12Mux_v I__1819 (
            .O(N__8139),
            .I(N__8131));
    Span12Mux_h I__1818 (
            .O(N__8136),
            .I(N__8131));
    Odrv12 I__1817 (
            .O(N__8131),
            .I(RnW_c));
    CascadeMux I__1816 (
            .O(N__8128),
            .I(N__8124));
    InMux I__1815 (
            .O(N__8127),
            .I(N__8113));
    InMux I__1814 (
            .O(N__8124),
            .I(N__8110));
    InMux I__1813 (
            .O(N__8123),
            .I(N__8106));
    CascadeMux I__1812 (
            .O(N__8122),
            .I(N__8100));
    CascadeMux I__1811 (
            .O(N__8121),
            .I(N__8093));
    InMux I__1810 (
            .O(N__8120),
            .I(N__8079));
    InMux I__1809 (
            .O(N__8119),
            .I(N__8079));
    InMux I__1808 (
            .O(N__8118),
            .I(N__8079));
    InMux I__1807 (
            .O(N__8117),
            .I(N__8079));
    InMux I__1806 (
            .O(N__8116),
            .I(N__8076));
    LocalMux I__1805 (
            .O(N__8113),
            .I(N__8070));
    LocalMux I__1804 (
            .O(N__8110),
            .I(N__8070));
    InMux I__1803 (
            .O(N__8109),
            .I(N__8067));
    LocalMux I__1802 (
            .O(N__8106),
            .I(N__8062));
    InMux I__1801 (
            .O(N__8105),
            .I(N__8057));
    InMux I__1800 (
            .O(N__8104),
            .I(N__8057));
    InMux I__1799 (
            .O(N__8103),
            .I(N__8054));
    InMux I__1798 (
            .O(N__8100),
            .I(N__8051));
    InMux I__1797 (
            .O(N__8099),
            .I(N__8048));
    InMux I__1796 (
            .O(N__8098),
            .I(N__8043));
    InMux I__1795 (
            .O(N__8097),
            .I(N__8043));
    InMux I__1794 (
            .O(N__8096),
            .I(N__8040));
    InMux I__1793 (
            .O(N__8093),
            .I(N__8037));
    InMux I__1792 (
            .O(N__8092),
            .I(N__8028));
    InMux I__1791 (
            .O(N__8091),
            .I(N__8028));
    InMux I__1790 (
            .O(N__8090),
            .I(N__8028));
    InMux I__1789 (
            .O(N__8089),
            .I(N__8028));
    CascadeMux I__1788 (
            .O(N__8088),
            .I(N__8025));
    LocalMux I__1787 (
            .O(N__8079),
            .I(N__8020));
    LocalMux I__1786 (
            .O(N__8076),
            .I(N__8017));
    InMux I__1785 (
            .O(N__8075),
            .I(N__8014));
    Span4Mux_v I__1784 (
            .O(N__8070),
            .I(N__8009));
    LocalMux I__1783 (
            .O(N__8067),
            .I(N__8009));
    InMux I__1782 (
            .O(N__8066),
            .I(N__8004));
    InMux I__1781 (
            .O(N__8065),
            .I(N__8004));
    Span4Mux_v I__1780 (
            .O(N__8062),
            .I(N__8001));
    LocalMux I__1779 (
            .O(N__8057),
            .I(N__7998));
    LocalMux I__1778 (
            .O(N__8054),
            .I(N__7991));
    LocalMux I__1777 (
            .O(N__8051),
            .I(N__7991));
    LocalMux I__1776 (
            .O(N__8048),
            .I(N__7991));
    LocalMux I__1775 (
            .O(N__8043),
            .I(N__7988));
    LocalMux I__1774 (
            .O(N__8040),
            .I(N__7985));
    LocalMux I__1773 (
            .O(N__8037),
            .I(N__7980));
    LocalMux I__1772 (
            .O(N__8028),
            .I(N__7980));
    InMux I__1771 (
            .O(N__8025),
            .I(N__7977));
    InMux I__1770 (
            .O(N__8024),
            .I(N__7974));
    InMux I__1769 (
            .O(N__8023),
            .I(N__7971));
    Span4Mux_h I__1768 (
            .O(N__8020),
            .I(N__7962));
    Span4Mux_h I__1767 (
            .O(N__8017),
            .I(N__7962));
    LocalMux I__1766 (
            .O(N__8014),
            .I(N__7962));
    Span4Mux_h I__1765 (
            .O(N__8009),
            .I(N__7962));
    LocalMux I__1764 (
            .O(N__8004),
            .I(N__7953));
    Span4Mux_h I__1763 (
            .O(N__8001),
            .I(N__7953));
    Span4Mux_h I__1762 (
            .O(N__7998),
            .I(N__7953));
    Span4Mux_h I__1761 (
            .O(N__7991),
            .I(N__7953));
    Span4Mux_h I__1760 (
            .O(N__7988),
            .I(N__7944));
    Span4Mux_h I__1759 (
            .O(N__7985),
            .I(N__7944));
    Span4Mux_h I__1758 (
            .O(N__7980),
            .I(N__7944));
    LocalMux I__1757 (
            .O(N__7977),
            .I(N__7944));
    LocalMux I__1756 (
            .O(N__7974),
            .I(CPU_CYCLEm));
    LocalMux I__1755 (
            .O(N__7971),
            .I(CPU_CYCLEm));
    Odrv4 I__1754 (
            .O(N__7962),
            .I(CPU_CYCLEm));
    Odrv4 I__1753 (
            .O(N__7953),
            .I(CPU_CYCLEm));
    Odrv4 I__1752 (
            .O(N__7944),
            .I(CPU_CYCLEm));
    InMux I__1751 (
            .O(N__7933),
            .I(N__7930));
    LocalMux I__1750 (
            .O(N__7930),
            .I(N__7926));
    InMux I__1749 (
            .O(N__7929),
            .I(N__7923));
    Sp12to4 I__1748 (
            .O(N__7926),
            .I(N__7920));
    LocalMux I__1747 (
            .O(N__7923),
            .I(N__7917));
    Span12Mux_v I__1746 (
            .O(N__7920),
            .I(N__7914));
    Span12Mux_v I__1745 (
            .O(N__7917),
            .I(N__7911));
    Span12Mux_h I__1744 (
            .O(N__7914),
            .I(N__7908));
    Span12Mux_h I__1743 (
            .O(N__7911),
            .I(N__7905));
    Odrv12 I__1742 (
            .O(N__7908),
            .I(AWEn_c));
    Odrv12 I__1741 (
            .O(N__7905),
            .I(AWEn_c));
    InMux I__1740 (
            .O(N__7900),
            .I(N__7897));
    LocalMux I__1739 (
            .O(N__7897),
            .I(\U712_CHIP_RAM.N_47 ));
    CascadeMux I__1738 (
            .O(N__7894),
            .I(N__7891));
    InMux I__1737 (
            .O(N__7891),
            .I(N__7888));
    LocalMux I__1736 (
            .O(N__7888),
            .I(N__7884));
    InMux I__1735 (
            .O(N__7887),
            .I(N__7877));
    Span4Mux_v I__1734 (
            .O(N__7884),
            .I(N__7874));
    InMux I__1733 (
            .O(N__7883),
            .I(N__7867));
    InMux I__1732 (
            .O(N__7882),
            .I(N__7867));
    InMux I__1731 (
            .O(N__7881),
            .I(N__7867));
    InMux I__1730 (
            .O(N__7880),
            .I(N__7864));
    LocalMux I__1729 (
            .O(N__7877),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1728 (
            .O(N__7874),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1727 (
            .O(N__7867),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1726 (
            .O(N__7864),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1725 (
            .O(N__7855),
            .I(N__7850));
    CascadeMux I__1724 (
            .O(N__7854),
            .I(N__7847));
    InMux I__1723 (
            .O(N__7853),
            .I(N__7844));
    LocalMux I__1722 (
            .O(N__7850),
            .I(N__7841));
    InMux I__1721 (
            .O(N__7847),
            .I(N__7836));
    LocalMux I__1720 (
            .O(N__7844),
            .I(N__7833));
    Span4Mux_h I__1719 (
            .O(N__7841),
            .I(N__7830));
    InMux I__1718 (
            .O(N__7840),
            .I(N__7825));
    InMux I__1717 (
            .O(N__7839),
            .I(N__7825));
    LocalMux I__1716 (
            .O(N__7836),
            .I(\U712_CHIP_RAM.N_63 ));
    Odrv4 I__1715 (
            .O(N__7833),
            .I(\U712_CHIP_RAM.N_63 ));
    Odrv4 I__1714 (
            .O(N__7830),
            .I(\U712_CHIP_RAM.N_63 ));
    LocalMux I__1713 (
            .O(N__7825),
            .I(\U712_CHIP_RAM.N_63 ));
    InMux I__1712 (
            .O(N__7816),
            .I(N__7812));
    InMux I__1711 (
            .O(N__7815),
            .I(N__7809));
    LocalMux I__1710 (
            .O(N__7812),
            .I(N__7803));
    LocalMux I__1709 (
            .O(N__7809),
            .I(N__7803));
    InMux I__1708 (
            .O(N__7808),
            .I(N__7800));
    Span4Mux_v I__1707 (
            .O(N__7803),
            .I(N__7792));
    LocalMux I__1706 (
            .O(N__7800),
            .I(N__7789));
    InMux I__1705 (
            .O(N__7799),
            .I(N__7784));
    InMux I__1704 (
            .O(N__7798),
            .I(N__7784));
    InMux I__1703 (
            .O(N__7797),
            .I(N__7781));
    InMux I__1702 (
            .O(N__7796),
            .I(N__7777));
    InMux I__1701 (
            .O(N__7795),
            .I(N__7774));
    Span4Mux_h I__1700 (
            .O(N__7792),
            .I(N__7767));
    Span4Mux_v I__1699 (
            .O(N__7789),
            .I(N__7767));
    LocalMux I__1698 (
            .O(N__7784),
            .I(N__7767));
    LocalMux I__1697 (
            .O(N__7781),
            .I(N__7764));
    InMux I__1696 (
            .O(N__7780),
            .I(N__7761));
    LocalMux I__1695 (
            .O(N__7777),
            .I(N__7758));
    LocalMux I__1694 (
            .O(N__7774),
            .I(N__7755));
    Span4Mux_h I__1693 (
            .O(N__7767),
            .I(N__7747));
    Span4Mux_v I__1692 (
            .O(N__7764),
            .I(N__7747));
    LocalMux I__1691 (
            .O(N__7761),
            .I(N__7744));
    Span4Mux_v I__1690 (
            .O(N__7758),
            .I(N__7739));
    Span4Mux_v I__1689 (
            .O(N__7755),
            .I(N__7739));
    InMux I__1688 (
            .O(N__7754),
            .I(N__7734));
    InMux I__1687 (
            .O(N__7753),
            .I(N__7734));
    InMux I__1686 (
            .O(N__7752),
            .I(N__7731));
    Span4Mux_h I__1685 (
            .O(N__7747),
            .I(N__7728));
    Span12Mux_v I__1684 (
            .O(N__7744),
            .I(N__7719));
    Sp12to4 I__1683 (
            .O(N__7739),
            .I(N__7719));
    LocalMux I__1682 (
            .O(N__7734),
            .I(N__7719));
    LocalMux I__1681 (
            .O(N__7731),
            .I(N__7719));
    Span4Mux_h I__1680 (
            .O(N__7728),
            .I(N__7716));
    Span12Mux_h I__1679 (
            .O(N__7719),
            .I(N__7713));
    Odrv4 I__1678 (
            .O(N__7716),
            .I(RESETn_c));
    Odrv12 I__1677 (
            .O(N__7713),
            .I(RESETn_c));
    CascadeMux I__1676 (
            .O(N__7708),
            .I(N__7703));
    InMux I__1675 (
            .O(N__7707),
            .I(N__7696));
    InMux I__1674 (
            .O(N__7706),
            .I(N__7696));
    InMux I__1673 (
            .O(N__7703),
            .I(N__7693));
    InMux I__1672 (
            .O(N__7702),
            .I(N__7688));
    InMux I__1671 (
            .O(N__7701),
            .I(N__7688));
    LocalMux I__1670 (
            .O(N__7696),
            .I(N__7685));
    LocalMux I__1669 (
            .O(N__7693),
            .I(N__7674));
    LocalMux I__1668 (
            .O(N__7688),
            .I(N__7669));
    Span4Mux_v I__1667 (
            .O(N__7685),
            .I(N__7669));
    InMux I__1666 (
            .O(N__7684),
            .I(N__7664));
    InMux I__1665 (
            .O(N__7683),
            .I(N__7664));
    InMux I__1664 (
            .O(N__7682),
            .I(N__7661));
    InMux I__1663 (
            .O(N__7681),
            .I(N__7654));
    InMux I__1662 (
            .O(N__7680),
            .I(N__7654));
    InMux I__1661 (
            .O(N__7679),
            .I(N__7654));
    InMux I__1660 (
            .O(N__7678),
            .I(N__7649));
    InMux I__1659 (
            .O(N__7677),
            .I(N__7649));
    Span4Mux_v I__1658 (
            .O(N__7674),
            .I(N__7646));
    Odrv4 I__1657 (
            .O(N__7669),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1656 (
            .O(N__7664),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1655 (
            .O(N__7661),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1654 (
            .O(N__7654),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1653 (
            .O(N__7649),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1652 (
            .O(N__7646),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__1651 (
            .O(N__7633),
            .I(\U712_CHIP_RAM.N_63_cascade_ ));
    CascadeMux I__1650 (
            .O(N__7630),
            .I(N__7625));
    CascadeMux I__1649 (
            .O(N__7629),
            .I(N__7621));
    InMux I__1648 (
            .O(N__7628),
            .I(N__7616));
    InMux I__1647 (
            .O(N__7625),
            .I(N__7616));
    CascadeMux I__1646 (
            .O(N__7624),
            .I(N__7612));
    InMux I__1645 (
            .O(N__7621),
            .I(N__7606));
    LocalMux I__1644 (
            .O(N__7616),
            .I(N__7603));
    InMux I__1643 (
            .O(N__7615),
            .I(N__7600));
    InMux I__1642 (
            .O(N__7612),
            .I(N__7597));
    InMux I__1641 (
            .O(N__7611),
            .I(N__7592));
    InMux I__1640 (
            .O(N__7610),
            .I(N__7592));
    InMux I__1639 (
            .O(N__7609),
            .I(N__7589));
    LocalMux I__1638 (
            .O(N__7606),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER46 ));
    Odrv12 I__1637 (
            .O(N__7603),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER46 ));
    LocalMux I__1636 (
            .O(N__7600),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER46 ));
    LocalMux I__1635 (
            .O(N__7597),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER46 ));
    LocalMux I__1634 (
            .O(N__7592),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER46 ));
    LocalMux I__1633 (
            .O(N__7589),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER46 ));
    InMux I__1632 (
            .O(N__7576),
            .I(N__7572));
    InMux I__1631 (
            .O(N__7575),
            .I(N__7566));
    LocalMux I__1630 (
            .O(N__7572),
            .I(N__7563));
    InMux I__1629 (
            .O(N__7571),
            .I(N__7560));
    InMux I__1628 (
            .O(N__7570),
            .I(N__7557));
    InMux I__1627 (
            .O(N__7569),
            .I(N__7554));
    LocalMux I__1626 (
            .O(N__7566),
            .I(\U712_CHIP_RAM.N_127 ));
    Odrv12 I__1625 (
            .O(N__7563),
            .I(\U712_CHIP_RAM.N_127 ));
    LocalMux I__1624 (
            .O(N__7560),
            .I(\U712_CHIP_RAM.N_127 ));
    LocalMux I__1623 (
            .O(N__7557),
            .I(\U712_CHIP_RAM.N_127 ));
    LocalMux I__1622 (
            .O(N__7554),
            .I(\U712_CHIP_RAM.N_127 ));
    InMux I__1621 (
            .O(N__7543),
            .I(N__7537));
    InMux I__1620 (
            .O(N__7542),
            .I(N__7537));
    LocalMux I__1619 (
            .O(N__7537),
            .I(N__7534));
    Span4Mux_v I__1618 (
            .O(N__7534),
            .I(N__7531));
    Odrv4 I__1617 (
            .O(N__7531),
            .I(\U712_CHIP_RAM.N_124 ));
    CascadeMux I__1616 (
            .O(N__7528),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_cascade_ ));
    CascadeMux I__1615 (
            .O(N__7525),
            .I(N__7518));
    CascadeMux I__1614 (
            .O(N__7524),
            .I(N__7515));
    InMux I__1613 (
            .O(N__7523),
            .I(N__7510));
    InMux I__1612 (
            .O(N__7522),
            .I(N__7507));
    InMux I__1611 (
            .O(N__7521),
            .I(N__7502));
    InMux I__1610 (
            .O(N__7518),
            .I(N__7502));
    InMux I__1609 (
            .O(N__7515),
            .I(N__7499));
    InMux I__1608 (
            .O(N__7514),
            .I(N__7494));
    InMux I__1607 (
            .O(N__7513),
            .I(N__7494));
    LocalMux I__1606 (
            .O(N__7510),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1605 (
            .O(N__7507),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1604 (
            .O(N__7502),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1603 (
            .O(N__7499),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1602 (
            .O(N__7494),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__1601 (
            .O(N__7483),
            .I(N__7480));
    LocalMux I__1600 (
            .O(N__7480),
            .I(\U712_CHIP_RAM.N_107 ));
    IoInMux I__1599 (
            .O(N__7477),
            .I(N__7474));
    LocalMux I__1598 (
            .O(N__7474),
            .I(N__7471));
    Span4Mux_s3_v I__1597 (
            .O(N__7471),
            .I(N__7468));
    Span4Mux_h I__1596 (
            .O(N__7468),
            .I(N__7464));
    CascadeMux I__1595 (
            .O(N__7467),
            .I(N__7461));
    Sp12to4 I__1594 (
            .O(N__7464),
            .I(N__7457));
    InMux I__1593 (
            .O(N__7461),
            .I(N__7454));
    CascadeMux I__1592 (
            .O(N__7460),
            .I(N__7451));
    Span12Mux_v I__1591 (
            .O(N__7457),
            .I(N__7448));
    LocalMux I__1590 (
            .O(N__7454),
            .I(N__7445));
    InMux I__1589 (
            .O(N__7451),
            .I(N__7442));
    Odrv12 I__1588 (
            .O(N__7448),
            .I(DBDIR_c));
    Odrv12 I__1587 (
            .O(N__7445),
            .I(DBDIR_c));
    LocalMux I__1586 (
            .O(N__7442),
            .I(DBDIR_c));
    IoInMux I__1585 (
            .O(N__7435),
            .I(N__7432));
    LocalMux I__1584 (
            .O(N__7432),
            .I(N__7429));
    Span4Mux_s1_h I__1583 (
            .O(N__7429),
            .I(N__7426));
    Sp12to4 I__1582 (
            .O(N__7426),
            .I(N__7423));
    Span12Mux_v I__1581 (
            .O(N__7423),
            .I(N__7420));
    Span12Mux_h I__1580 (
            .O(N__7420),
            .I(N__7417));
    Odrv12 I__1579 (
            .O(N__7417),
            .I(DRDDIR_0_i));
    IoInMux I__1578 (
            .O(N__7414),
            .I(N__7411));
    LocalMux I__1577 (
            .O(N__7411),
            .I(N__7408));
    Span4Mux_s2_v I__1576 (
            .O(N__7408),
            .I(N__7405));
    Span4Mux_v I__1575 (
            .O(N__7405),
            .I(N__7402));
    Span4Mux_v I__1574 (
            .O(N__7402),
            .I(N__7399));
    Odrv4 I__1573 (
            .O(N__7399),
            .I(CMA_c_10));
    CEMux I__1572 (
            .O(N__7396),
            .I(N__7389));
    CEMux I__1571 (
            .O(N__7395),
            .I(N__7386));
    CEMux I__1570 (
            .O(N__7394),
            .I(N__7383));
    CEMux I__1569 (
            .O(N__7393),
            .I(N__7380));
    CEMux I__1568 (
            .O(N__7392),
            .I(N__7376));
    LocalMux I__1567 (
            .O(N__7389),
            .I(N__7373));
    LocalMux I__1566 (
            .O(N__7386),
            .I(N__7368));
    LocalMux I__1565 (
            .O(N__7383),
            .I(N__7368));
    LocalMux I__1564 (
            .O(N__7380),
            .I(N__7365));
    CEMux I__1563 (
            .O(N__7379),
            .I(N__7362));
    LocalMux I__1562 (
            .O(N__7376),
            .I(N__7359));
    Span4Mux_h I__1561 (
            .O(N__7373),
            .I(N__7354));
    Span4Mux_v I__1560 (
            .O(N__7368),
            .I(N__7354));
    Span4Mux_v I__1559 (
            .O(N__7365),
            .I(N__7351));
    LocalMux I__1558 (
            .O(N__7362),
            .I(N__7348));
    Span4Mux_h I__1557 (
            .O(N__7359),
            .I(N__7345));
    Span4Mux_h I__1556 (
            .O(N__7354),
            .I(N__7342));
    Span4Mux_v I__1555 (
            .O(N__7351),
            .I(N__7339));
    Odrv12 I__1554 (
            .O(N__7348),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv4 I__1553 (
            .O(N__7345),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv4 I__1552 (
            .O(N__7342),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv4 I__1551 (
            .O(N__7339),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    InMux I__1550 (
            .O(N__7330),
            .I(N__7326));
    InMux I__1549 (
            .O(N__7329),
            .I(N__7323));
    LocalMux I__1548 (
            .O(N__7326),
            .I(N__7320));
    LocalMux I__1547 (
            .O(N__7323),
            .I(N__7317));
    Span4Mux_v I__1546 (
            .O(N__7320),
            .I(N__7314));
    Span12Mux_v I__1545 (
            .O(N__7317),
            .I(N__7309));
    Sp12to4 I__1544 (
            .O(N__7314),
            .I(N__7309));
    Span12Mux_h I__1543 (
            .O(N__7309),
            .I(N__7306));
    Odrv12 I__1542 (
            .O(N__7306),
            .I(DRA_c_7));
    InMux I__1541 (
            .O(N__7303),
            .I(N__7300));
    LocalMux I__1540 (
            .O(N__7300),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__1539 (
            .O(N__7297),
            .I(N__7294));
    LocalMux I__1538 (
            .O(N__7294),
            .I(N__7290));
    InMux I__1537 (
            .O(N__7293),
            .I(N__7287));
    Span4Mux_v I__1536 (
            .O(N__7290),
            .I(N__7284));
    LocalMux I__1535 (
            .O(N__7287),
            .I(N__7281));
    Sp12to4 I__1534 (
            .O(N__7284),
            .I(N__7278));
    Span4Mux_v I__1533 (
            .O(N__7281),
            .I(N__7275));
    Span12Mux_h I__1532 (
            .O(N__7278),
            .I(N__7272));
    Sp12to4 I__1531 (
            .O(N__7275),
            .I(N__7269));
    Odrv12 I__1530 (
            .O(N__7272),
            .I(DRA_c_8));
    Odrv12 I__1529 (
            .O(N__7269),
            .I(DRA_c_8));
    InMux I__1528 (
            .O(N__7264),
            .I(N__7261));
    LocalMux I__1527 (
            .O(N__7261),
            .I(N__7258));
    Odrv4 I__1526 (
            .O(N__7258),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__1525 (
            .O(N__7255),
            .I(N__7252));
    LocalMux I__1524 (
            .O(N__7252),
            .I(N__7248));
    InMux I__1523 (
            .O(N__7251),
            .I(N__7245));
    Odrv4 I__1522 (
            .O(N__7248),
            .I(\U712_CHIP_RAM.N_65 ));
    LocalMux I__1521 (
            .O(N__7245),
            .I(\U712_CHIP_RAM.N_65 ));
    InMux I__1520 (
            .O(N__7240),
            .I(N__7237));
    LocalMux I__1519 (
            .O(N__7237),
            .I(N__7232));
    InMux I__1518 (
            .O(N__7236),
            .I(N__7229));
    InMux I__1517 (
            .O(N__7235),
            .I(N__7226));
    Odrv12 I__1516 (
            .O(N__7232),
            .I(\U712_CHIP_RAM.N_78 ));
    LocalMux I__1515 (
            .O(N__7229),
            .I(\U712_CHIP_RAM.N_78 ));
    LocalMux I__1514 (
            .O(N__7226),
            .I(\U712_CHIP_RAM.N_78 ));
    InMux I__1513 (
            .O(N__7219),
            .I(N__7214));
    InMux I__1512 (
            .O(N__7218),
            .I(N__7211));
    InMux I__1511 (
            .O(N__7217),
            .I(N__7208));
    LocalMux I__1510 (
            .O(N__7214),
            .I(N__7204));
    LocalMux I__1509 (
            .O(N__7211),
            .I(N__7199));
    LocalMux I__1508 (
            .O(N__7208),
            .I(N__7199));
    InMux I__1507 (
            .O(N__7207),
            .I(N__7194));
    Span4Mux_h I__1506 (
            .O(N__7204),
            .I(N__7189));
    Span4Mux_h I__1505 (
            .O(N__7199),
            .I(N__7186));
    InMux I__1504 (
            .O(N__7198),
            .I(N__7181));
    InMux I__1503 (
            .O(N__7197),
            .I(N__7181));
    LocalMux I__1502 (
            .O(N__7194),
            .I(N__7178));
    InMux I__1501 (
            .O(N__7193),
            .I(N__7173));
    InMux I__1500 (
            .O(N__7192),
            .I(N__7173));
    Odrv4 I__1499 (
            .O(N__7189),
            .I(\U712_CHIP_RAM.N_67 ));
    Odrv4 I__1498 (
            .O(N__7186),
            .I(\U712_CHIP_RAM.N_67 ));
    LocalMux I__1497 (
            .O(N__7181),
            .I(\U712_CHIP_RAM.N_67 ));
    Odrv4 I__1496 (
            .O(N__7178),
            .I(\U712_CHIP_RAM.N_67 ));
    LocalMux I__1495 (
            .O(N__7173),
            .I(\U712_CHIP_RAM.N_67 ));
    CascadeMux I__1494 (
            .O(N__7162),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_cascade_ ));
    InMux I__1493 (
            .O(N__7159),
            .I(N__7156));
    LocalMux I__1492 (
            .O(N__7156),
            .I(N__7153));
    Span4Mux_v I__1491 (
            .O(N__7153),
            .I(N__7150));
    Odrv4 I__1490 (
            .O(N__7150),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__1489 (
            .O(N__7147),
            .I(N__7144));
    LocalMux I__1488 (
            .O(N__7144),
            .I(N__7141));
    Span4Mux_v I__1487 (
            .O(N__7141),
            .I(N__7138));
    Odrv4 I__1486 (
            .O(N__7138),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_5 ));
    InMux I__1485 (
            .O(N__7135),
            .I(N__7131));
    InMux I__1484 (
            .O(N__7134),
            .I(N__7128));
    LocalMux I__1483 (
            .O(N__7131),
            .I(\U712_CHIP_RAM.N_77 ));
    LocalMux I__1482 (
            .O(N__7128),
            .I(\U712_CHIP_RAM.N_77 ));
    CascadeMux I__1481 (
            .O(N__7123),
            .I(\U712_CHIP_RAM.N_80_cascade_ ));
    CascadeMux I__1480 (
            .O(N__7120),
            .I(\U712_CHIP_RAM.N_50_cascade_ ));
    InMux I__1479 (
            .O(N__7117),
            .I(N__7113));
    InMux I__1478 (
            .O(N__7116),
            .I(N__7108));
    LocalMux I__1477 (
            .O(N__7113),
            .I(N__7105));
    InMux I__1476 (
            .O(N__7112),
            .I(N__7102));
    InMux I__1475 (
            .O(N__7111),
            .I(N__7099));
    LocalMux I__1474 (
            .O(N__7108),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    Odrv4 I__1473 (
            .O(N__7105),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__1472 (
            .O(N__7102),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__1471 (
            .O(N__7099),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__1470 (
            .O(N__7090),
            .I(N__7085));
    CascadeMux I__1469 (
            .O(N__7089),
            .I(N__7082));
    InMux I__1468 (
            .O(N__7088),
            .I(N__7079));
    LocalMux I__1467 (
            .O(N__7085),
            .I(N__7076));
    InMux I__1466 (
            .O(N__7082),
            .I(N__7073));
    LocalMux I__1465 (
            .O(N__7079),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    Odrv4 I__1464 (
            .O(N__7076),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__1463 (
            .O(N__7073),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    CascadeMux I__1462 (
            .O(N__7066),
            .I(N__7062));
    InMux I__1461 (
            .O(N__7065),
            .I(N__7055));
    InMux I__1460 (
            .O(N__7062),
            .I(N__7055));
    InMux I__1459 (
            .O(N__7061),
            .I(N__7052));
    InMux I__1458 (
            .O(N__7060),
            .I(N__7049));
    LocalMux I__1457 (
            .O(N__7055),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__1456 (
            .O(N__7052),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__1455 (
            .O(N__7049),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__1454 (
            .O(N__7042),
            .I(N__7036));
    InMux I__1453 (
            .O(N__7041),
            .I(N__7036));
    LocalMux I__1452 (
            .O(N__7036),
            .I(\U712_CHIP_RAM.N_60 ));
    InMux I__1451 (
            .O(N__7033),
            .I(N__7030));
    LocalMux I__1450 (
            .O(N__7030),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER39_0 ));
    CascadeMux I__1449 (
            .O(N__7027),
            .I(N__7022));
    CascadeMux I__1448 (
            .O(N__7026),
            .I(N__7019));
    InMux I__1447 (
            .O(N__7025),
            .I(N__7016));
    InMux I__1446 (
            .O(N__7022),
            .I(N__7009));
    InMux I__1445 (
            .O(N__7019),
            .I(N__7009));
    LocalMux I__1444 (
            .O(N__7016),
            .I(N__7006));
    InMux I__1443 (
            .O(N__7015),
            .I(N__7003));
    InMux I__1442 (
            .O(N__7014),
            .I(N__7000));
    LocalMux I__1441 (
            .O(N__7009),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    Odrv4 I__1440 (
            .O(N__7006),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1439 (
            .O(N__7003),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1438 (
            .O(N__7000),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__1437 (
            .O(N__6991),
            .I(N__6985));
    InMux I__1436 (
            .O(N__6990),
            .I(N__6985));
    LocalMux I__1435 (
            .O(N__6985),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER39_2 ));
    InMux I__1434 (
            .O(N__6982),
            .I(N__6978));
    InMux I__1433 (
            .O(N__6981),
            .I(N__6969));
    LocalMux I__1432 (
            .O(N__6978),
            .I(N__6966));
    CascadeMux I__1431 (
            .O(N__6977),
            .I(N__6963));
    CascadeMux I__1430 (
            .O(N__6976),
            .I(N__6960));
    CascadeMux I__1429 (
            .O(N__6975),
            .I(N__6951));
    CascadeMux I__1428 (
            .O(N__6974),
            .I(N__6948));
    InMux I__1427 (
            .O(N__6973),
            .I(N__6944));
    InMux I__1426 (
            .O(N__6972),
            .I(N__6941));
    LocalMux I__1425 (
            .O(N__6969),
            .I(N__6938));
    Span4Mux_h I__1424 (
            .O(N__6966),
            .I(N__6935));
    InMux I__1423 (
            .O(N__6963),
            .I(N__6932));
    InMux I__1422 (
            .O(N__6960),
            .I(N__6929));
    InMux I__1421 (
            .O(N__6959),
            .I(N__6926));
    InMux I__1420 (
            .O(N__6958),
            .I(N__6921));
    InMux I__1419 (
            .O(N__6957),
            .I(N__6921));
    InMux I__1418 (
            .O(N__6956),
            .I(N__6916));
    InMux I__1417 (
            .O(N__6955),
            .I(N__6916));
    InMux I__1416 (
            .O(N__6954),
            .I(N__6907));
    InMux I__1415 (
            .O(N__6951),
            .I(N__6907));
    InMux I__1414 (
            .O(N__6948),
            .I(N__6907));
    InMux I__1413 (
            .O(N__6947),
            .I(N__6907));
    LocalMux I__1412 (
            .O(N__6944),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1411 (
            .O(N__6941),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv12 I__1410 (
            .O(N__6938),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1409 (
            .O(N__6935),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1408 (
            .O(N__6932),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1407 (
            .O(N__6929),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1406 (
            .O(N__6926),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1405 (
            .O(N__6921),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1404 (
            .O(N__6916),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1403 (
            .O(N__6907),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1402 (
            .O(N__6886),
            .I(N__6882));
    InMux I__1401 (
            .O(N__6885),
            .I(N__6879));
    LocalMux I__1400 (
            .O(N__6882),
            .I(\U712_CHIP_RAM.N_50 ));
    LocalMux I__1399 (
            .O(N__6879),
            .I(\U712_CHIP_RAM.N_50 ));
    CascadeMux I__1398 (
            .O(N__6874),
            .I(N__6869));
    CascadeMux I__1397 (
            .O(N__6873),
            .I(N__6865));
    CascadeMux I__1396 (
            .O(N__6872),
            .I(N__6858));
    InMux I__1395 (
            .O(N__6869),
            .I(N__6848));
    InMux I__1394 (
            .O(N__6868),
            .I(N__6848));
    InMux I__1393 (
            .O(N__6865),
            .I(N__6843));
    InMux I__1392 (
            .O(N__6864),
            .I(N__6838));
    InMux I__1391 (
            .O(N__6863),
            .I(N__6838));
    CascadeMux I__1390 (
            .O(N__6862),
            .I(N__6834));
    InMux I__1389 (
            .O(N__6861),
            .I(N__6830));
    InMux I__1388 (
            .O(N__6858),
            .I(N__6827));
    InMux I__1387 (
            .O(N__6857),
            .I(N__6820));
    InMux I__1386 (
            .O(N__6856),
            .I(N__6820));
    InMux I__1385 (
            .O(N__6855),
            .I(N__6820));
    CascadeMux I__1384 (
            .O(N__6854),
            .I(N__6817));
    CascadeMux I__1383 (
            .O(N__6853),
            .I(N__6814));
    LocalMux I__1382 (
            .O(N__6848),
            .I(N__6811));
    InMux I__1381 (
            .O(N__6847),
            .I(N__6808));
    InMux I__1380 (
            .O(N__6846),
            .I(N__6801));
    LocalMux I__1379 (
            .O(N__6843),
            .I(N__6796));
    LocalMux I__1378 (
            .O(N__6838),
            .I(N__6796));
    InMux I__1377 (
            .O(N__6837),
            .I(N__6791));
    InMux I__1376 (
            .O(N__6834),
            .I(N__6791));
    InMux I__1375 (
            .O(N__6833),
            .I(N__6788));
    LocalMux I__1374 (
            .O(N__6830),
            .I(N__6781));
    LocalMux I__1373 (
            .O(N__6827),
            .I(N__6781));
    LocalMux I__1372 (
            .O(N__6820),
            .I(N__6781));
    InMux I__1371 (
            .O(N__6817),
            .I(N__6776));
    InMux I__1370 (
            .O(N__6814),
            .I(N__6776));
    Span12Mux_v I__1369 (
            .O(N__6811),
            .I(N__6771));
    LocalMux I__1368 (
            .O(N__6808),
            .I(N__6771));
    InMux I__1367 (
            .O(N__6807),
            .I(N__6762));
    InMux I__1366 (
            .O(N__6806),
            .I(N__6762));
    InMux I__1365 (
            .O(N__6805),
            .I(N__6762));
    InMux I__1364 (
            .O(N__6804),
            .I(N__6762));
    LocalMux I__1363 (
            .O(N__6801),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv12 I__1362 (
            .O(N__6796),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1361 (
            .O(N__6791),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1360 (
            .O(N__6788),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1359 (
            .O(N__6781),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1358 (
            .O(N__6776),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv12 I__1357 (
            .O(N__6771),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1356 (
            .O(N__6762),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1355 (
            .O(N__6745),
            .I(N__6740));
    InMux I__1354 (
            .O(N__6744),
            .I(N__6735));
    InMux I__1353 (
            .O(N__6743),
            .I(N__6735));
    LocalMux I__1352 (
            .O(N__6740),
            .I(N__6732));
    LocalMux I__1351 (
            .O(N__6735),
            .I(N__6729));
    Span4Mux_v I__1350 (
            .O(N__6732),
            .I(N__6726));
    Sp12to4 I__1349 (
            .O(N__6729),
            .I(N__6723));
    Sp12to4 I__1348 (
            .O(N__6726),
            .I(N__6720));
    Span12Mux_v I__1347 (
            .O(N__6723),
            .I(N__6717));
    Span12Mux_h I__1346 (
            .O(N__6720),
            .I(N__6714));
    Span12Mux_h I__1345 (
            .O(N__6717),
            .I(N__6711));
    Span12Mux_v I__1344 (
            .O(N__6714),
            .I(N__6708));
    Odrv12 I__1343 (
            .O(N__6711),
            .I(CASLn_c));
    Odrv12 I__1342 (
            .O(N__6708),
            .I(CASLn_c));
    InMux I__1341 (
            .O(N__6703),
            .I(N__6697));
    InMux I__1340 (
            .O(N__6702),
            .I(N__6697));
    LocalMux I__1339 (
            .O(N__6697),
            .I(N__6693));
    InMux I__1338 (
            .O(N__6696),
            .I(N__6690));
    Span4Mux_h I__1337 (
            .O(N__6693),
            .I(N__6687));
    LocalMux I__1336 (
            .O(N__6690),
            .I(N__6684));
    Sp12to4 I__1335 (
            .O(N__6687),
            .I(N__6679));
    Sp12to4 I__1334 (
            .O(N__6684),
            .I(N__6679));
    Span12Mux_v I__1333 (
            .O(N__6679),
            .I(N__6676));
    Span12Mux_h I__1332 (
            .O(N__6676),
            .I(N__6673));
    Odrv12 I__1331 (
            .O(N__6673),
            .I(CASUn_c));
    CascadeMux I__1330 (
            .O(N__6670),
            .I(N__6666));
    InMux I__1329 (
            .O(N__6669),
            .I(N__6662));
    InMux I__1328 (
            .O(N__6666),
            .I(N__6657));
    InMux I__1327 (
            .O(N__6665),
            .I(N__6657));
    LocalMux I__1326 (
            .O(N__6662),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    LocalMux I__1325 (
            .O(N__6657),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__1324 (
            .O(N__6652),
            .I(N__6646));
    InMux I__1323 (
            .O(N__6651),
            .I(N__6646));
    LocalMux I__1322 (
            .O(N__6646),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__1321 (
            .O(N__6643),
            .I(N__6640));
    LocalMux I__1320 (
            .O(N__6640),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_2_1 ));
    InMux I__1319 (
            .O(N__6637),
            .I(N__6634));
    LocalMux I__1318 (
            .O(N__6634),
            .I(N__6631));
    Odrv4 I__1317 (
            .O(N__6631),
            .I(\U712_CHIP_RAM.N_108 ));
    CascadeMux I__1316 (
            .O(N__6628),
            .I(\U712_CHIP_RAM.N_77_cascade_ ));
    InMux I__1315 (
            .O(N__6625),
            .I(N__6622));
    LocalMux I__1314 (
            .O(N__6622),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1 ));
    InMux I__1313 (
            .O(N__6619),
            .I(N__6616));
    LocalMux I__1312 (
            .O(N__6616),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_0 ));
    CascadeMux I__1311 (
            .O(N__6613),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_ ));
    InMux I__1310 (
            .O(N__6610),
            .I(N__6607));
    LocalMux I__1309 (
            .O(N__6607),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ));
    CascadeMux I__1308 (
            .O(N__6604),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_ ));
    CEMux I__1307 (
            .O(N__6601),
            .I(N__6598));
    LocalMux I__1306 (
            .O(N__6598),
            .I(N__6595));
    Span4Mux_h I__1305 (
            .O(N__6595),
            .I(N__6592));
    Span4Mux_h I__1304 (
            .O(N__6592),
            .I(N__6589));
    Odrv4 I__1303 (
            .O(N__6589),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0 ));
    InMux I__1302 (
            .O(N__6586),
            .I(N__6579));
    InMux I__1301 (
            .O(N__6585),
            .I(N__6579));
    InMux I__1300 (
            .O(N__6584),
            .I(N__6576));
    LocalMux I__1299 (
            .O(N__6579),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4 ));
    LocalMux I__1298 (
            .O(N__6576),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4 ));
    InMux I__1297 (
            .O(N__6571),
            .I(N__6568));
    LocalMux I__1296 (
            .O(N__6568),
            .I(\U712_CHIP_RAM.N_80 ));
    InMux I__1295 (
            .O(N__6565),
            .I(N__6562));
    LocalMux I__1294 (
            .O(N__6562),
            .I(N__6559));
    Odrv12 I__1293 (
            .O(N__6559),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__1292 (
            .O(N__6556),
            .I(N__6553));
    LocalMux I__1291 (
            .O(N__6553),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    InMux I__1290 (
            .O(N__6550),
            .I(N__6546));
    InMux I__1289 (
            .O(N__6549),
            .I(N__6543));
    LocalMux I__1288 (
            .O(N__6546),
            .I(N__6540));
    LocalMux I__1287 (
            .O(N__6543),
            .I(N__6537));
    Sp12to4 I__1286 (
            .O(N__6540),
            .I(N__6534));
    Span12Mux_v I__1285 (
            .O(N__6537),
            .I(N__6531));
    Span12Mux_v I__1284 (
            .O(N__6534),
            .I(N__6528));
    Span12Mux_h I__1283 (
            .O(N__6531),
            .I(N__6525));
    Span12Mux_h I__1282 (
            .O(N__6528),
            .I(N__6522));
    Odrv12 I__1281 (
            .O(N__6525),
            .I(DRA_c_4));
    Odrv12 I__1280 (
            .O(N__6522),
            .I(DRA_c_4));
    InMux I__1279 (
            .O(N__6517),
            .I(N__6514));
    LocalMux I__1278 (
            .O(N__6514),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__1277 (
            .O(N__6511),
            .I(N__6508));
    LocalMux I__1276 (
            .O(N__6508),
            .I(N__6505));
    Span4Mux_v I__1275 (
            .O(N__6505),
            .I(N__6501));
    InMux I__1274 (
            .O(N__6504),
            .I(N__6498));
    Odrv4 I__1273 (
            .O(N__6501),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_1_a3_0 ));
    LocalMux I__1272 (
            .O(N__6498),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_1_a3_0 ));
    InMux I__1271 (
            .O(N__6493),
            .I(N__6490));
    LocalMux I__1270 (
            .O(N__6490),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i ));
    InMux I__1269 (
            .O(N__6487),
            .I(N__6481));
    InMux I__1268 (
            .O(N__6486),
            .I(N__6481));
    LocalMux I__1267 (
            .O(N__6481),
            .I(N__6478));
    Odrv4 I__1266 (
            .O(N__6478),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6 ));
    InMux I__1265 (
            .O(N__6475),
            .I(N__6472));
    LocalMux I__1264 (
            .O(N__6472),
            .I(N__6469));
    Span4Mux_h I__1263 (
            .O(N__6469),
            .I(N__6466));
    Span4Mux_h I__1262 (
            .O(N__6466),
            .I(N__6463));
    Odrv4 I__1261 (
            .O(N__6463),
            .I(\U712_REG_SM.N_173_0 ));
    InMux I__1260 (
            .O(N__6460),
            .I(N__6457));
    LocalMux I__1259 (
            .O(N__6457),
            .I(N__6454));
    Span4Mux_h I__1258 (
            .O(N__6454),
            .I(N__6451));
    Span4Mux_h I__1257 (
            .O(N__6451),
            .I(N__6447));
    InMux I__1256 (
            .O(N__6450),
            .I(N__6444));
    Odrv4 I__1255 (
            .O(N__6447),
            .I(\U712_REG_SM.N_183_1 ));
    LocalMux I__1254 (
            .O(N__6444),
            .I(\U712_REG_SM.N_183_1 ));
    CascadeMux I__1253 (
            .O(N__6439),
            .I(N__6436));
    InMux I__1252 (
            .O(N__6436),
            .I(N__6433));
    LocalMux I__1251 (
            .O(N__6433),
            .I(N__6430));
    Span4Mux_h I__1250 (
            .O(N__6430),
            .I(N__6427));
    Span4Mux_h I__1249 (
            .O(N__6427),
            .I(N__6423));
    InMux I__1248 (
            .O(N__6426),
            .I(N__6420));
    Odrv4 I__1247 (
            .O(N__6423),
            .I(\U712_REG_SM.N_165_0 ));
    LocalMux I__1246 (
            .O(N__6420),
            .I(\U712_REG_SM.N_165_0 ));
    InMux I__1245 (
            .O(N__6415),
            .I(N__6412));
    LocalMux I__1244 (
            .O(N__6412),
            .I(N__6408));
    InMux I__1243 (
            .O(N__6411),
            .I(N__6405));
    Span4Mux_h I__1242 (
            .O(N__6408),
            .I(N__6399));
    LocalMux I__1241 (
            .O(N__6405),
            .I(N__6399));
    InMux I__1240 (
            .O(N__6404),
            .I(N__6396));
    Span4Mux_h I__1239 (
            .O(N__6399),
            .I(N__6393));
    LocalMux I__1238 (
            .O(N__6396),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    Odrv4 I__1237 (
            .O(N__6393),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    InMux I__1236 (
            .O(N__6388),
            .I(N__6384));
    InMux I__1235 (
            .O(N__6387),
            .I(N__6381));
    LocalMux I__1234 (
            .O(N__6384),
            .I(N__6372));
    LocalMux I__1233 (
            .O(N__6381),
            .I(N__6372));
    InMux I__1232 (
            .O(N__6380),
            .I(N__6369));
    InMux I__1231 (
            .O(N__6379),
            .I(N__6366));
    InMux I__1230 (
            .O(N__6378),
            .I(N__6363));
    InMux I__1229 (
            .O(N__6377),
            .I(N__6360));
    Span4Mux_h I__1228 (
            .O(N__6372),
            .I(N__6355));
    LocalMux I__1227 (
            .O(N__6369),
            .I(N__6355));
    LocalMux I__1226 (
            .O(N__6366),
            .I(N__6352));
    LocalMux I__1225 (
            .O(N__6363),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1224 (
            .O(N__6360),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1223 (
            .O(N__6355),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1222 (
            .O(N__6352),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    CascadeMux I__1221 (
            .O(N__6343),
            .I(N__6340));
    InMux I__1220 (
            .O(N__6340),
            .I(N__6337));
    LocalMux I__1219 (
            .O(N__6337),
            .I(N__6333));
    InMux I__1218 (
            .O(N__6336),
            .I(N__6330));
    Span4Mux_h I__1217 (
            .O(N__6333),
            .I(N__6327));
    LocalMux I__1216 (
            .O(N__6330),
            .I(\U712_CHIP_RAM.un1_DBR_SYNC ));
    Odrv4 I__1215 (
            .O(N__6327),
            .I(\U712_CHIP_RAM.un1_DBR_SYNC ));
    CEMux I__1214 (
            .O(N__6322),
            .I(N__6319));
    LocalMux I__1213 (
            .O(N__6319),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0 ));
    InMux I__1212 (
            .O(N__6316),
            .I(N__6313));
    LocalMux I__1211 (
            .O(N__6313),
            .I(N__6309));
    InMux I__1210 (
            .O(N__6312),
            .I(N__6306));
    Span4Mux_h I__1209 (
            .O(N__6309),
            .I(N__6300));
    LocalMux I__1208 (
            .O(N__6306),
            .I(N__6300));
    InMux I__1207 (
            .O(N__6305),
            .I(N__6297));
    Odrv4 I__1206 (
            .O(N__6300),
            .I(\U712_REG_SM.DS_ENZ0 ));
    LocalMux I__1205 (
            .O(N__6297),
            .I(\U712_REG_SM.DS_ENZ0 ));
    InMux I__1204 (
            .O(N__6292),
            .I(N__6289));
    LocalMux I__1203 (
            .O(N__6289),
            .I(N__6285));
    CascadeMux I__1202 (
            .O(N__6288),
            .I(N__6282));
    Span4Mux_v I__1201 (
            .O(N__6285),
            .I(N__6279));
    InMux I__1200 (
            .O(N__6282),
            .I(N__6276));
    Odrv4 I__1199 (
            .O(N__6279),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    LocalMux I__1198 (
            .O(N__6276),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    IoInMux I__1197 (
            .O(N__6271),
            .I(N__6268));
    LocalMux I__1196 (
            .O(N__6268),
            .I(N__6265));
    IoSpan4Mux I__1195 (
            .O(N__6265),
            .I(N__6262));
    Span4Mux_s3_v I__1194 (
            .O(N__6262),
            .I(N__6259));
    Sp12to4 I__1193 (
            .O(N__6259),
            .I(N__6256));
    Span12Mux_s11_v I__1192 (
            .O(N__6256),
            .I(N__6253));
    Odrv12 I__1191 (
            .O(N__6253),
            .I(U712_REG_SM_un1_LDSn_i));
    InMux I__1190 (
            .O(N__6250),
            .I(N__6247));
    LocalMux I__1189 (
            .O(N__6247),
            .I(N__6244));
    Odrv4 I__1188 (
            .O(N__6244),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ));
    InMux I__1187 (
            .O(N__6241),
            .I(N__6237));
    InMux I__1186 (
            .O(N__6240),
            .I(N__6234));
    LocalMux I__1185 (
            .O(N__6237),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__1184 (
            .O(N__6234),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    CascadeMux I__1183 (
            .O(N__6229),
            .I(N__6225));
    InMux I__1182 (
            .O(N__6228),
            .I(N__6222));
    InMux I__1181 (
            .O(N__6225),
            .I(N__6219));
    LocalMux I__1180 (
            .O(N__6222),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__1179 (
            .O(N__6219),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__1178 (
            .O(N__6214),
            .I(N__6211));
    LocalMux I__1177 (
            .O(N__6211),
            .I(N__6208));
    Odrv4 I__1176 (
            .O(N__6208),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    IoInMux I__1175 (
            .O(N__6205),
            .I(N__6202));
    LocalMux I__1174 (
            .O(N__6202),
            .I(N__6199));
    IoSpan4Mux I__1173 (
            .O(N__6199),
            .I(N__6196));
    IoSpan4Mux I__1172 (
            .O(N__6196),
            .I(N__6193));
    Span4Mux_s2_h I__1171 (
            .O(N__6193),
            .I(N__6190));
    Sp12to4 I__1170 (
            .O(N__6190),
            .I(N__6187));
    Odrv12 I__1169 (
            .O(N__6187),
            .I(CMA_c_7));
    InMux I__1168 (
            .O(N__6184),
            .I(N__6181));
    LocalMux I__1167 (
            .O(N__6181),
            .I(N__6178));
    Span4Mux_v I__1166 (
            .O(N__6178),
            .I(N__6175));
    Span4Mux_v I__1165 (
            .O(N__6175),
            .I(N__6172));
    Sp12to4 I__1164 (
            .O(N__6172),
            .I(N__6169));
    Span12Mux_h I__1163 (
            .O(N__6169),
            .I(N__6166));
    Odrv12 I__1162 (
            .O(N__6166),
            .I(A_c_18));
    CascadeMux I__1161 (
            .O(N__6163),
            .I(N__6160));
    InMux I__1160 (
            .O(N__6160),
            .I(N__6157));
    LocalMux I__1159 (
            .O(N__6157),
            .I(N__6154));
    Span4Mux_v I__1158 (
            .O(N__6154),
            .I(N__6151));
    Span4Mux_v I__1157 (
            .O(N__6151),
            .I(N__6148));
    Sp12to4 I__1156 (
            .O(N__6148),
            .I(N__6145));
    Span12Mux_h I__1155 (
            .O(N__6145),
            .I(N__6142));
    Odrv12 I__1154 (
            .O(N__6142),
            .I(A_c_16));
    InMux I__1153 (
            .O(N__6139),
            .I(N__6136));
    LocalMux I__1152 (
            .O(N__6136),
            .I(\U712_CHIP_RAM.N_39 ));
    InMux I__1151 (
            .O(N__6133),
            .I(N__6130));
    LocalMux I__1150 (
            .O(N__6130),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_7 ));
    CascadeMux I__1149 (
            .O(N__6127),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_0_cascade_ ));
    CEMux I__1148 (
            .O(N__6124),
            .I(N__6120));
    CEMux I__1147 (
            .O(N__6123),
            .I(N__6117));
    LocalMux I__1146 (
            .O(N__6120),
            .I(N__6114));
    LocalMux I__1145 (
            .O(N__6117),
            .I(N__6111));
    Odrv4 I__1144 (
            .O(N__6114),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_i ));
    Odrv4 I__1143 (
            .O(N__6111),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_i ));
    CascadeMux I__1142 (
            .O(N__6106),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_5_cascade_ ));
    InMux I__1141 (
            .O(N__6103),
            .I(N__6100));
    LocalMux I__1140 (
            .O(N__6100),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER18_0 ));
    CascadeMux I__1139 (
            .O(N__6097),
            .I(N__6094));
    InMux I__1138 (
            .O(N__6094),
            .I(N__6091));
    LocalMux I__1137 (
            .O(N__6091),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__1136 (
            .O(N__6088),
            .I(N__6085));
    LocalMux I__1135 (
            .O(N__6085),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_4 ));
    InMux I__1134 (
            .O(N__6082),
            .I(N__6078));
    InMux I__1133 (
            .O(N__6081),
            .I(N__6075));
    LocalMux I__1132 (
            .O(N__6078),
            .I(\U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa ));
    LocalMux I__1131 (
            .O(N__6075),
            .I(\U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa ));
    InMux I__1130 (
            .O(N__6070),
            .I(N__6066));
    InMux I__1129 (
            .O(N__6069),
            .I(N__6063));
    LocalMux I__1128 (
            .O(N__6066),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER18_0 ));
    LocalMux I__1127 (
            .O(N__6063),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER18_0 ));
    CascadeMux I__1126 (
            .O(N__6058),
            .I(\U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa_cascade_ ));
    CascadeMux I__1125 (
            .O(N__6055),
            .I(N__6050));
    CascadeMux I__1124 (
            .O(N__6054),
            .I(N__6046));
    InMux I__1123 (
            .O(N__6053),
            .I(N__6043));
    InMux I__1122 (
            .O(N__6050),
            .I(N__6040));
    InMux I__1121 (
            .O(N__6049),
            .I(N__6037));
    InMux I__1120 (
            .O(N__6046),
            .I(N__6034));
    LocalMux I__1119 (
            .O(N__6043),
            .I(\U712_CHIP_RAM.N_158_0 ));
    LocalMux I__1118 (
            .O(N__6040),
            .I(\U712_CHIP_RAM.N_158_0 ));
    LocalMux I__1117 (
            .O(N__6037),
            .I(\U712_CHIP_RAM.N_158_0 ));
    LocalMux I__1116 (
            .O(N__6034),
            .I(\U712_CHIP_RAM.N_158_0 ));
    InMux I__1115 (
            .O(N__6025),
            .I(N__6022));
    LocalMux I__1114 (
            .O(N__6022),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_ns_1_1 ));
    CascadeMux I__1113 (
            .O(N__6019),
            .I(N__6016));
    InMux I__1112 (
            .O(N__6016),
            .I(N__6013));
    LocalMux I__1111 (
            .O(N__6013),
            .I(\U712_CHIP_RAM.N_132 ));
    SRMux I__1110 (
            .O(N__6010),
            .I(N__6007));
    LocalMux I__1109 (
            .O(N__6007),
            .I(N__6004));
    Odrv4 I__1108 (
            .O(N__6004),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__1107 (
            .O(N__6001),
            .I(N__5998));
    LocalMux I__1106 (
            .O(N__5998),
            .I(N__5995));
    Odrv12 I__1105 (
            .O(N__5995),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__1104 (
            .O(N__5992),
            .I(N__5989));
    LocalMux I__1103 (
            .O(N__5989),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__1102 (
            .O(N__5986),
            .I(N__5983));
    LocalMux I__1101 (
            .O(N__5983),
            .I(N__5980));
    Span4Mux_v I__1100 (
            .O(N__5980),
            .I(N__5977));
    Sp12to4 I__1099 (
            .O(N__5977),
            .I(N__5974));
    Span12Mux_h I__1098 (
            .O(N__5974),
            .I(N__5971));
    Span12Mux_v I__1097 (
            .O(N__5971),
            .I(N__5968));
    Odrv12 I__1096 (
            .O(N__5968),
            .I(A_c_17));
    CascadeMux I__1095 (
            .O(N__5965),
            .I(\U712_CHIP_RAM.CMA_5_0_8_cascade_ ));
    IoInMux I__1094 (
            .O(N__5962),
            .I(N__5959));
    LocalMux I__1093 (
            .O(N__5959),
            .I(N__5956));
    IoSpan4Mux I__1092 (
            .O(N__5956),
            .I(N__5953));
    Span4Mux_s3_h I__1091 (
            .O(N__5953),
            .I(N__5950));
    Sp12to4 I__1090 (
            .O(N__5950),
            .I(N__5947));
    Span12Mux_h I__1089 (
            .O(N__5947),
            .I(N__5944));
    Odrv12 I__1088 (
            .O(N__5944),
            .I(CMA_c_8));
    InMux I__1087 (
            .O(N__5941),
            .I(N__5938));
    LocalMux I__1086 (
            .O(N__5938),
            .I(N__5935));
    Odrv4 I__1085 (
            .O(N__5935),
            .I(\U712_CHIP_RAM.N_38 ));
    IoInMux I__1084 (
            .O(N__5932),
            .I(N__5929));
    LocalMux I__1083 (
            .O(N__5929),
            .I(N__5926));
    Span4Mux_s2_h I__1082 (
            .O(N__5926),
            .I(N__5923));
    Sp12to4 I__1081 (
            .O(N__5923),
            .I(N__5920));
    Span12Mux_s6_v I__1080 (
            .O(N__5920),
            .I(N__5917));
    Span12Mux_h I__1079 (
            .O(N__5917),
            .I(N__5914));
    Odrv12 I__1078 (
            .O(N__5914),
            .I(CMA_c_6));
    InMux I__1077 (
            .O(N__5911),
            .I(N__5908));
    LocalMux I__1076 (
            .O(N__5908),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    CascadeMux I__1075 (
            .O(N__5905),
            .I(N__5902));
    InMux I__1074 (
            .O(N__5902),
            .I(N__5899));
    LocalMux I__1073 (
            .O(N__5899),
            .I(N__5896));
    Span4Mux_h I__1072 (
            .O(N__5896),
            .I(N__5893));
    Sp12to4 I__1071 (
            .O(N__5893),
            .I(N__5890));
    Span12Mux_v I__1070 (
            .O(N__5890),
            .I(N__5887));
    Span12Mux_h I__1069 (
            .O(N__5887),
            .I(N__5884));
    Odrv12 I__1068 (
            .O(N__5884),
            .I(A_c_19));
    IoInMux I__1067 (
            .O(N__5881),
            .I(N__5878));
    LocalMux I__1066 (
            .O(N__5878),
            .I(N__5875));
    Span4Mux_s3_h I__1065 (
            .O(N__5875),
            .I(N__5872));
    Span4Mux_v I__1064 (
            .O(N__5872),
            .I(N__5869));
    Span4Mux_v I__1063 (
            .O(N__5869),
            .I(N__5866));
    Sp12to4 I__1062 (
            .O(N__5866),
            .I(N__5863));
    Odrv12 I__1061 (
            .O(N__5863),
            .I(CMA_c_9));
    InMux I__1060 (
            .O(N__5860),
            .I(N__5857));
    LocalMux I__1059 (
            .O(N__5857),
            .I(N__5853));
    InMux I__1058 (
            .O(N__5856),
            .I(N__5850));
    Span12Mux_v I__1057 (
            .O(N__5853),
            .I(N__5847));
    LocalMux I__1056 (
            .O(N__5850),
            .I(N__5844));
    Span12Mux_v I__1055 (
            .O(N__5847),
            .I(N__5841));
    Span12Mux_h I__1054 (
            .O(N__5844),
            .I(N__5838));
    Span12Mux_h I__1053 (
            .O(N__5841),
            .I(N__5835));
    Span12Mux_v I__1052 (
            .O(N__5838),
            .I(N__5832));
    Odrv12 I__1051 (
            .O(N__5835),
            .I(DRA_c_1));
    Odrv12 I__1050 (
            .O(N__5832),
            .I(DRA_c_1));
    InMux I__1049 (
            .O(N__5827),
            .I(N__5824));
    LocalMux I__1048 (
            .O(N__5824),
            .I(N__5821));
    Odrv4 I__1047 (
            .O(N__5821),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1046 (
            .O(N__5818),
            .I(N__5815));
    LocalMux I__1045 (
            .O(N__5815),
            .I(N__5811));
    InMux I__1044 (
            .O(N__5814),
            .I(N__5808));
    Sp12to4 I__1043 (
            .O(N__5811),
            .I(N__5803));
    LocalMux I__1042 (
            .O(N__5808),
            .I(N__5803));
    Span12Mux_v I__1041 (
            .O(N__5803),
            .I(N__5800));
    Span12Mux_h I__1040 (
            .O(N__5800),
            .I(N__5797));
    Odrv12 I__1039 (
            .O(N__5797),
            .I(DRA_c_6));
    InMux I__1038 (
            .O(N__5794),
            .I(N__5791));
    LocalMux I__1037 (
            .O(N__5791),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    IoInMux I__1036 (
            .O(N__5788),
            .I(N__5785));
    LocalMux I__1035 (
            .O(N__5785),
            .I(N__5782));
    Span4Mux_s0_v I__1034 (
            .O(N__5782),
            .I(N__5779));
    Sp12to4 I__1033 (
            .O(N__5779),
            .I(N__5776));
    Span12Mux_h I__1032 (
            .O(N__5776),
            .I(N__5773));
    Span12Mux_v I__1031 (
            .O(N__5773),
            .I(N__5765));
    InMux I__1030 (
            .O(N__5772),
            .I(N__5756));
    InMux I__1029 (
            .O(N__5771),
            .I(N__5756));
    InMux I__1028 (
            .O(N__5770),
            .I(N__5756));
    InMux I__1027 (
            .O(N__5769),
            .I(N__5756));
    InMux I__1026 (
            .O(N__5768),
            .I(N__5753));
    Odrv12 I__1025 (
            .O(N__5765),
            .I(DBENn_c));
    LocalMux I__1024 (
            .O(N__5756),
            .I(DBENn_c));
    LocalMux I__1023 (
            .O(N__5753),
            .I(DBENn_c));
    IoInMux I__1022 (
            .O(N__5746),
            .I(N__5743));
    LocalMux I__1021 (
            .O(N__5743),
            .I(N__5740));
    Span4Mux_s3_h I__1020 (
            .O(N__5740),
            .I(N__5737));
    Sp12to4 I__1019 (
            .O(N__5737),
            .I(N__5734));
    Span12Mux_v I__1018 (
            .O(N__5734),
            .I(N__5731));
    Span12Mux_h I__1017 (
            .O(N__5731),
            .I(N__5728));
    Odrv12 I__1016 (
            .O(N__5728),
            .I(CUUBEn_c));
    InMux I__1015 (
            .O(N__5725),
            .I(N__5721));
    InMux I__1014 (
            .O(N__5724),
            .I(N__5718));
    LocalMux I__1013 (
            .O(N__5721),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ));
    LocalMux I__1012 (
            .O(N__5718),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ));
    InMux I__1011 (
            .O(N__5713),
            .I(bfn_14_4_0_));
    InMux I__1010 (
            .O(N__5710),
            .I(N__5706));
    InMux I__1009 (
            .O(N__5709),
            .I(N__5703));
    LocalMux I__1008 (
            .O(N__5706),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__1007 (
            .O(N__5703),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__1006 (
            .O(N__5698),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__1005 (
            .O(N__5695),
            .I(N__5691));
    InMux I__1004 (
            .O(N__5694),
            .I(N__5688));
    LocalMux I__1003 (
            .O(N__5691),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__1002 (
            .O(N__5688),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    InMux I__1001 (
            .O(N__5683),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__1000 (
            .O(N__5680),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    CascadeMux I__999 (
            .O(N__5677),
            .I(N__5673));
    InMux I__998 (
            .O(N__5676),
            .I(N__5670));
    InMux I__997 (
            .O(N__5673),
            .I(N__5667));
    LocalMux I__996 (
            .O(N__5670),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__995 (
            .O(N__5667),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__994 (
            .O(N__5662),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__993 (
            .O(N__5659),
            .I(N__5655));
    InMux I__992 (
            .O(N__5658),
            .I(N__5652));
    LocalMux I__991 (
            .O(N__5655),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__990 (
            .O(N__5652),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__989 (
            .O(N__5647),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__988 (
            .O(N__5644),
            .I(N__5640));
    InMux I__987 (
            .O(N__5643),
            .I(N__5637));
    LocalMux I__986 (
            .O(N__5640),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__985 (
            .O(N__5637),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__984 (
            .O(N__5632),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__983 (
            .O(N__5629),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__982 (
            .O(N__5626),
            .I(N__5623));
    GlobalMux I__981 (
            .O(N__5623),
            .I(N__5620));
    gio2CtrlBuf I__980 (
            .O(N__5620),
            .I(C1_c_g));
    InMux I__979 (
            .O(N__5617),
            .I(N__5613));
    InMux I__978 (
            .O(N__5616),
            .I(N__5610));
    LocalMux I__977 (
            .O(N__5613),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0 ));
    LocalMux I__976 (
            .O(N__5610),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0 ));
    InMux I__975 (
            .O(N__5605),
            .I(N__5602));
    LocalMux I__974 (
            .O(N__5602),
            .I(N__5599));
    Span4Mux_h I__973 (
            .O(N__5599),
            .I(N__5596));
    Odrv4 I__972 (
            .O(N__5596),
            .I(\U712_CHIP_RAM.DMA_CYCLE_7 ));
    CascadeMux I__971 (
            .O(N__5593),
            .I(\U712_BYTE_ENABLE.un2_CUMBEnZ0_cascade_ ));
    IoInMux I__970 (
            .O(N__5590),
            .I(N__5587));
    LocalMux I__969 (
            .O(N__5587),
            .I(N__5584));
    Span4Mux_s3_h I__968 (
            .O(N__5584),
            .I(N__5581));
    Span4Mux_v I__967 (
            .O(N__5581),
            .I(N__5578));
    Sp12to4 I__966 (
            .O(N__5578),
            .I(N__5575));
    Span12Mux_h I__965 (
            .O(N__5575),
            .I(N__5572));
    Span12Mux_v I__964 (
            .O(N__5572),
            .I(N__5569));
    Odrv12 I__963 (
            .O(N__5569),
            .I(CUMBEn_c));
    InMux I__962 (
            .O(N__5566),
            .I(N__5560));
    InMux I__961 (
            .O(N__5565),
            .I(N__5560));
    LocalMux I__960 (
            .O(N__5560),
            .I(\U712_BYTE_ENABLE.LLBE_0_0_tz ));
    CascadeMux I__959 (
            .O(N__5557),
            .I(\U712_BYTE_ENABLE.un2_CLLBEnZ0_cascade_ ));
    IoInMux I__958 (
            .O(N__5554),
            .I(N__5551));
    LocalMux I__957 (
            .O(N__5551),
            .I(N__5548));
    IoSpan4Mux I__956 (
            .O(N__5548),
            .I(N__5545));
    Sp12to4 I__955 (
            .O(N__5545),
            .I(N__5542));
    Span12Mux_s7_v I__954 (
            .O(N__5542),
            .I(N__5539));
    Span12Mux_v I__953 (
            .O(N__5539),
            .I(N__5536));
    Odrv12 I__952 (
            .O(N__5536),
            .I(CLLBEn_c));
    CascadeMux I__951 (
            .O(N__5533),
            .I(\U712_BYTE_ENABLE.un2_CLMBEnZ0_cascade_ ));
    IoInMux I__950 (
            .O(N__5530),
            .I(N__5527));
    LocalMux I__949 (
            .O(N__5527),
            .I(N__5524));
    Span4Mux_s3_h I__948 (
            .O(N__5524),
            .I(N__5521));
    Sp12to4 I__947 (
            .O(N__5521),
            .I(N__5518));
    Span12Mux_v I__946 (
            .O(N__5518),
            .I(N__5515));
    Span12Mux_h I__945 (
            .O(N__5515),
            .I(N__5512));
    Odrv12 I__944 (
            .O(N__5512),
            .I(CLMBEn_c));
    InMux I__943 (
            .O(N__5509),
            .I(N__5497));
    InMux I__942 (
            .O(N__5508),
            .I(N__5497));
    InMux I__941 (
            .O(N__5507),
            .I(N__5497));
    InMux I__940 (
            .O(N__5506),
            .I(N__5497));
    LocalMux I__939 (
            .O(N__5497),
            .I(N__5494));
    Span4Mux_v I__938 (
            .O(N__5494),
            .I(N__5491));
    Span4Mux_v I__937 (
            .O(N__5491),
            .I(N__5488));
    Sp12to4 I__936 (
            .O(N__5488),
            .I(N__5485));
    Span12Mux_h I__935 (
            .O(N__5485),
            .I(N__5482));
    Odrv12 I__934 (
            .O(N__5482),
            .I(A_c_1));
    InMux I__933 (
            .O(N__5479),
            .I(N__5470));
    InMux I__932 (
            .O(N__5478),
            .I(N__5470));
    InMux I__931 (
            .O(N__5477),
            .I(N__5467));
    InMux I__930 (
            .O(N__5476),
            .I(N__5462));
    InMux I__929 (
            .O(N__5475),
            .I(N__5462));
    LocalMux I__928 (
            .O(N__5470),
            .I(N__5457));
    LocalMux I__927 (
            .O(N__5467),
            .I(N__5457));
    LocalMux I__926 (
            .O(N__5462),
            .I(N__5454));
    Span4Mux_v I__925 (
            .O(N__5457),
            .I(N__5451));
    Span4Mux_v I__924 (
            .O(N__5454),
            .I(N__5448));
    Sp12to4 I__923 (
            .O(N__5451),
            .I(N__5443));
    Sp12to4 I__922 (
            .O(N__5448),
            .I(N__5443));
    Span12Mux_h I__921 (
            .O(N__5443),
            .I(N__5440));
    Odrv12 I__920 (
            .O(N__5440),
            .I(A_c_0));
    CascadeMux I__919 (
            .O(N__5437),
            .I(N__5431));
    CascadeMux I__918 (
            .O(N__5436),
            .I(N__5428));
    CascadeMux I__917 (
            .O(N__5435),
            .I(N__5425));
    CascadeMux I__916 (
            .O(N__5434),
            .I(N__5422));
    InMux I__915 (
            .O(N__5431),
            .I(N__5413));
    InMux I__914 (
            .O(N__5428),
            .I(N__5413));
    InMux I__913 (
            .O(N__5425),
            .I(N__5413));
    InMux I__912 (
            .O(N__5422),
            .I(N__5413));
    LocalMux I__911 (
            .O(N__5413),
            .I(N__5410));
    Odrv4 I__910 (
            .O(N__5410),
            .I(\U712_BYTE_ENABLE.LW_TRANS_0 ));
    CascadeMux I__909 (
            .O(N__5407),
            .I(\U712_BYTE_ENABLE.un2_CUUBEnZ0_cascade_ ));
    InMux I__908 (
            .O(N__5404),
            .I(N__5398));
    InMux I__907 (
            .O(N__5403),
            .I(N__5398));
    LocalMux I__906 (
            .O(N__5398),
            .I(N__5395));
    Odrv4 I__905 (
            .O(N__5395),
            .I(\U712_CHIP_RAM.N_51 ));
    CascadeMux I__904 (
            .O(N__5392),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER16_2_0_cascade_ ));
    CascadeMux I__903 (
            .O(N__5389),
            .I(\U712_CHIP_RAM.N_99_cascade_ ));
    CascadeMux I__902 (
            .O(N__5386),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_cascade_ ));
    CascadeMux I__901 (
            .O(N__5383),
            .I(\U712_CHIP_RAM.N_67_cascade_ ));
    CascadeMux I__900 (
            .O(N__5380),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER18_0_cascade_ ));
    CascadeMux I__899 (
            .O(N__5377),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_m2_3_cascade_ ));
    InMux I__898 (
            .O(N__5374),
            .I(N__5371));
    LocalMux I__897 (
            .O(N__5371),
            .I(\U712_CHIP_RAM.N_35 ));
    IoInMux I__896 (
            .O(N__5368),
            .I(N__5365));
    LocalMux I__895 (
            .O(N__5365),
            .I(N__5362));
    Span4Mux_s3_h I__894 (
            .O(N__5362),
            .I(N__5359));
    Sp12to4 I__893 (
            .O(N__5359),
            .I(N__5356));
    Span12Mux_s6_v I__892 (
            .O(N__5356),
            .I(N__5353));
    Span12Mux_h I__891 (
            .O(N__5353),
            .I(N__5350));
    Odrv12 I__890 (
            .O(N__5350),
            .I(CMA_c_3));
    InMux I__889 (
            .O(N__5347),
            .I(N__5344));
    LocalMux I__888 (
            .O(N__5344),
            .I(N__5341));
    Span4Mux_v I__887 (
            .O(N__5341),
            .I(N__5338));
    Sp12to4 I__886 (
            .O(N__5338),
            .I(N__5335));
    Span12Mux_h I__885 (
            .O(N__5335),
            .I(N__5332));
    Odrv12 I__884 (
            .O(N__5332),
            .I(A_c_6));
    CascadeMux I__883 (
            .O(N__5329),
            .I(N__5326));
    InMux I__882 (
            .O(N__5326),
            .I(N__5323));
    LocalMux I__881 (
            .O(N__5323),
            .I(N__5320));
    Span4Mux_v I__880 (
            .O(N__5320),
            .I(N__5317));
    Span4Mux_v I__879 (
            .O(N__5317),
            .I(N__5314));
    Sp12to4 I__878 (
            .O(N__5314),
            .I(N__5311));
    Span12Mux_h I__877 (
            .O(N__5311),
            .I(N__5308));
    Odrv12 I__876 (
            .O(N__5308),
            .I(A_c_13));
    CascadeMux I__875 (
            .O(N__5305),
            .I(\U712_CHIP_RAM.N_36_cascade_ ));
    IoInMux I__874 (
            .O(N__5302),
            .I(N__5299));
    LocalMux I__873 (
            .O(N__5299),
            .I(N__5296));
    IoSpan4Mux I__872 (
            .O(N__5296),
            .I(N__5293));
    Sp12to4 I__871 (
            .O(N__5293),
            .I(N__5290));
    Span12Mux_s9_v I__870 (
            .O(N__5290),
            .I(N__5287));
    Span12Mux_h I__869 (
            .O(N__5287),
            .I(N__5284));
    Odrv12 I__868 (
            .O(N__5284),
            .I(CMA_c_4));
    InMux I__867 (
            .O(N__5281),
            .I(N__5278));
    LocalMux I__866 (
            .O(N__5278),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_ns_1_2 ));
    CascadeMux I__865 (
            .O(N__5275),
            .I(\U712_CHIP_RAM.N_61_cascade_ ));
    CascadeMux I__864 (
            .O(N__5272),
            .I(\U712_CHIP_RAM.N_65_cascade_ ));
    InMux I__863 (
            .O(N__5269),
            .I(N__5266));
    LocalMux I__862 (
            .O(N__5266),
            .I(\U712_CHIP_RAM.N_104_1 ));
    InMux I__861 (
            .O(N__5263),
            .I(N__5260));
    LocalMux I__860 (
            .O(N__5260),
            .I(N__5257));
    Span4Mux_v I__859 (
            .O(N__5257),
            .I(N__5254));
    Sp12to4 I__858 (
            .O(N__5254),
            .I(N__5251));
    Span12Mux_h I__857 (
            .O(N__5251),
            .I(N__5248));
    Odrv12 I__856 (
            .O(N__5248),
            .I(A_c_9));
    CascadeMux I__855 (
            .O(N__5245),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_ ));
    InMux I__854 (
            .O(N__5242),
            .I(N__5239));
    LocalMux I__853 (
            .O(N__5239),
            .I(N__5236));
    Span4Mux_v I__852 (
            .O(N__5236),
            .I(N__5233));
    Sp12to4 I__851 (
            .O(N__5233),
            .I(N__5230));
    Span12Mux_h I__850 (
            .O(N__5230),
            .I(N__5227));
    Span12Mux_v I__849 (
            .O(N__5227),
            .I(N__5224));
    Odrv12 I__848 (
            .O(N__5224),
            .I(A_c_2));
    InMux I__847 (
            .O(N__5221),
            .I(N__5218));
    LocalMux I__846 (
            .O(N__5218),
            .I(\U712_CHIP_RAM.N_32 ));
    InMux I__845 (
            .O(N__5215),
            .I(N__5212));
    LocalMux I__844 (
            .O(N__5212),
            .I(N__5209));
    Odrv4 I__843 (
            .O(N__5209),
            .I(\U712_CHIP_RAM.N_37 ));
    IoInMux I__842 (
            .O(N__5206),
            .I(N__5203));
    LocalMux I__841 (
            .O(N__5203),
            .I(N__5200));
    Span4Mux_s3_h I__840 (
            .O(N__5200),
            .I(N__5197));
    Span4Mux_v I__839 (
            .O(N__5197),
            .I(N__5194));
    Sp12to4 I__838 (
            .O(N__5194),
            .I(N__5191));
    Span12Mux_h I__837 (
            .O(N__5191),
            .I(N__5188));
    Odrv12 I__836 (
            .O(N__5188),
            .I(CMA_c_5));
    InMux I__835 (
            .O(N__5185),
            .I(N__5181));
    InMux I__834 (
            .O(N__5184),
            .I(N__5178));
    LocalMux I__833 (
            .O(N__5181),
            .I(N__5173));
    LocalMux I__832 (
            .O(N__5178),
            .I(N__5173));
    Span4Mux_v I__831 (
            .O(N__5173),
            .I(N__5170));
    Span4Mux_v I__830 (
            .O(N__5170),
            .I(N__5167));
    Sp12to4 I__829 (
            .O(N__5167),
            .I(N__5164));
    Span12Mux_h I__828 (
            .O(N__5164),
            .I(N__5161));
    Odrv12 I__827 (
            .O(N__5161),
            .I(DRA_c_3));
    InMux I__826 (
            .O(N__5158),
            .I(N__5155));
    LocalMux I__825 (
            .O(N__5155),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__824 (
            .O(N__5152),
            .I(N__5149));
    LocalMux I__823 (
            .O(N__5149),
            .I(N__5145));
    InMux I__822 (
            .O(N__5148),
            .I(N__5142));
    Span4Mux_v I__821 (
            .O(N__5145),
            .I(N__5139));
    LocalMux I__820 (
            .O(N__5142),
            .I(N__5136));
    Sp12to4 I__819 (
            .O(N__5139),
            .I(N__5133));
    Sp12to4 I__818 (
            .O(N__5136),
            .I(N__5130));
    Span12Mux_h I__817 (
            .O(N__5133),
            .I(N__5127));
    Span12Mux_v I__816 (
            .O(N__5130),
            .I(N__5124));
    Span12Mux_v I__815 (
            .O(N__5127),
            .I(N__5121));
    Span12Mux_h I__814 (
            .O(N__5124),
            .I(N__5118));
    Odrv12 I__813 (
            .O(N__5121),
            .I(DRA_c_2));
    Odrv12 I__812 (
            .O(N__5118),
            .I(DRA_c_2));
    InMux I__811 (
            .O(N__5113),
            .I(N__5110));
    LocalMux I__810 (
            .O(N__5110),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__809 (
            .O(N__5107),
            .I(N__5104));
    LocalMux I__808 (
            .O(N__5104),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__807 (
            .O(N__5101),
            .I(N__5098));
    LocalMux I__806 (
            .O(N__5098),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__805 (
            .O(N__5095),
            .I(N__5092));
    LocalMux I__804 (
            .O(N__5092),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_5 ));
    InMux I__803 (
            .O(N__5089),
            .I(N__5085));
    InMux I__802 (
            .O(N__5088),
            .I(N__5082));
    LocalMux I__801 (
            .O(N__5085),
            .I(N__5077));
    LocalMux I__800 (
            .O(N__5082),
            .I(N__5077));
    Span4Mux_v I__799 (
            .O(N__5077),
            .I(N__5074));
    Span4Mux_v I__798 (
            .O(N__5074),
            .I(N__5071));
    Sp12to4 I__797 (
            .O(N__5071),
            .I(N__5068));
    Span12Mux_h I__796 (
            .O(N__5068),
            .I(N__5065));
    Odrv12 I__795 (
            .O(N__5065),
            .I(DRA_c_5));
    CascadeMux I__794 (
            .O(N__5062),
            .I(N__5059));
    InMux I__793 (
            .O(N__5059),
            .I(N__5056));
    LocalMux I__792 (
            .O(N__5056),
            .I(N__5052));
    InMux I__791 (
            .O(N__5055),
            .I(N__5049));
    Odrv4 I__790 (
            .O(N__5052),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__789 (
            .O(N__5049),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__788 (
            .O(N__5044),
            .I(N__5040));
    CascadeMux I__787 (
            .O(N__5043),
            .I(N__5033));
    LocalMux I__786 (
            .O(N__5040),
            .I(N__5030));
    InMux I__785 (
            .O(N__5039),
            .I(N__5027));
    InMux I__784 (
            .O(N__5038),
            .I(N__5024));
    InMux I__783 (
            .O(N__5037),
            .I(N__5017));
    InMux I__782 (
            .O(N__5036),
            .I(N__5017));
    InMux I__781 (
            .O(N__5033),
            .I(N__5017));
    Span4Mux_h I__780 (
            .O(N__5030),
            .I(N__5014));
    LocalMux I__779 (
            .O(N__5027),
            .I(N__5007));
    LocalMux I__778 (
            .O(N__5024),
            .I(N__5007));
    LocalMux I__777 (
            .O(N__5017),
            .I(N__5007));
    Odrv4 I__776 (
            .O(N__5014),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    Odrv12 I__775 (
            .O(N__5007),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    CascadeMux I__774 (
            .O(N__5002),
            .I(N__4999));
    InMux I__773 (
            .O(N__4999),
            .I(N__4996));
    LocalMux I__772 (
            .O(N__4996),
            .I(N__4993));
    Odrv4 I__771 (
            .O(N__4993),
            .I(\U712_REG_SM.RnW_m ));
    InMux I__770 (
            .O(N__4990),
            .I(N__4987));
    LocalMux I__769 (
            .O(N__4987),
            .I(\U712_REG_SM.un1_LDS_OUT_0_sqmuxa_1_0 ));
    InMux I__768 (
            .O(N__4984),
            .I(N__4981));
    LocalMux I__767 (
            .O(N__4981),
            .I(N__4978));
    Span12Mux_h I__766 (
            .O(N__4978),
            .I(N__4975));
    Span12Mux_v I__765 (
            .O(N__4975),
            .I(N__4972));
    Odrv12 I__764 (
            .O(N__4972),
            .I(DBRn_c));
    InMux I__763 (
            .O(N__4969),
            .I(N__4965));
    CascadeMux I__762 (
            .O(N__4968),
            .I(N__4962));
    LocalMux I__761 (
            .O(N__4965),
            .I(N__4959));
    InMux I__760 (
            .O(N__4962),
            .I(N__4956));
    Span4Mux_v I__759 (
            .O(N__4959),
            .I(N__4952));
    LocalMux I__758 (
            .O(N__4956),
            .I(N__4949));
    InMux I__757 (
            .O(N__4955),
            .I(N__4945));
    Sp12to4 I__756 (
            .O(N__4952),
            .I(N__4940));
    Span12Mux_v I__755 (
            .O(N__4949),
            .I(N__4940));
    InMux I__754 (
            .O(N__4948),
            .I(N__4937));
    LocalMux I__753 (
            .O(N__4945),
            .I(U712_REG_SM_DBR_SYNC_0));
    Odrv12 I__752 (
            .O(N__4940),
            .I(U712_REG_SM_DBR_SYNC_0));
    LocalMux I__751 (
            .O(N__4937),
            .I(U712_REG_SM_DBR_SYNC_0));
    InMux I__750 (
            .O(N__4930),
            .I(N__4926));
    InMux I__749 (
            .O(N__4929),
            .I(N__4923));
    LocalMux I__748 (
            .O(N__4926),
            .I(N__4918));
    LocalMux I__747 (
            .O(N__4923),
            .I(N__4918));
    Span4Mux_h I__746 (
            .O(N__4918),
            .I(N__4914));
    InMux I__745 (
            .O(N__4917),
            .I(N__4911));
    Odrv4 I__744 (
            .O(N__4914),
            .I(U712_REG_SM_DBR_SYNC_1));
    LocalMux I__743 (
            .O(N__4911),
            .I(U712_REG_SM_DBR_SYNC_1));
    InMux I__742 (
            .O(N__4906),
            .I(N__4903));
    LocalMux I__741 (
            .O(N__4903),
            .I(N__4899));
    InMux I__740 (
            .O(N__4902),
            .I(N__4896));
    Span4Mux_v I__739 (
            .O(N__4899),
            .I(N__4893));
    LocalMux I__738 (
            .O(N__4896),
            .I(N__4890));
    Span4Mux_h I__737 (
            .O(N__4893),
            .I(N__4887));
    Span4Mux_v I__736 (
            .O(N__4890),
            .I(N__4884));
    Sp12to4 I__735 (
            .O(N__4887),
            .I(N__4879));
    Sp12to4 I__734 (
            .O(N__4884),
            .I(N__4879));
    Span12Mux_h I__733 (
            .O(N__4879),
            .I(N__4876));
    Span12Mux_v I__732 (
            .O(N__4876),
            .I(N__4873));
    Odrv12 I__731 (
            .O(N__4873),
            .I(SIZ_c_1));
    InMux I__730 (
            .O(N__4870),
            .I(N__4866));
    CascadeMux I__729 (
            .O(N__4869),
            .I(N__4863));
    LocalMux I__728 (
            .O(N__4866),
            .I(N__4860));
    InMux I__727 (
            .O(N__4863),
            .I(N__4857));
    Odrv4 I__726 (
            .O(N__4860),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    LocalMux I__725 (
            .O(N__4857),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    IoInMux I__724 (
            .O(N__4852),
            .I(N__4849));
    LocalMux I__723 (
            .O(N__4849),
            .I(N__4846));
    Span4Mux_s3_v I__722 (
            .O(N__4846),
            .I(N__4843));
    Span4Mux_v I__721 (
            .O(N__4843),
            .I(N__4840));
    Span4Mux_v I__720 (
            .O(N__4840),
            .I(N__4837));
    Sp12to4 I__719 (
            .O(N__4837),
            .I(N__4834));
    Odrv12 I__718 (
            .O(N__4834),
            .I(U712_REG_SM_un1_UDSn_i));
    IoInMux I__717 (
            .O(N__4831),
            .I(N__4828));
    LocalMux I__716 (
            .O(N__4828),
            .I(N__4825));
    Odrv12 I__715 (
            .O(N__4825),
            .I(RESETn_c_i));
    InMux I__714 (
            .O(N__4822),
            .I(N__4819));
    LocalMux I__713 (
            .O(N__4819),
            .I(N__4816));
    Span12Mux_v I__712 (
            .O(N__4816),
            .I(N__4813));
    Span12Mux_h I__711 (
            .O(N__4813),
            .I(N__4810));
    Odrv12 I__710 (
            .O(N__4810),
            .I(A_c_15));
    InMux I__709 (
            .O(N__4807),
            .I(N__4804));
    LocalMux I__708 (
            .O(N__4804),
            .I(N__4801));
    Span4Mux_v I__707 (
            .O(N__4801),
            .I(N__4798));
    Sp12to4 I__706 (
            .O(N__4798),
            .I(N__4795));
    Span12Mux_h I__705 (
            .O(N__4795),
            .I(N__4792));
    Odrv12 I__704 (
            .O(N__4792),
            .I(A_c_8));
    CascadeMux I__703 (
            .O(N__4789),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_6_cascade_ ));
    InMux I__702 (
            .O(N__4786),
            .I(N__4783));
    LocalMux I__701 (
            .O(N__4783),
            .I(N__4780));
    Span12Mux_v I__700 (
            .O(N__4780),
            .I(N__4777));
    Span12Mux_h I__699 (
            .O(N__4777),
            .I(N__4774));
    Odrv12 I__698 (
            .O(N__4774),
            .I(A_c_5));
    CascadeMux I__697 (
            .O(N__4771),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_ ));
    InMux I__696 (
            .O(N__4768),
            .I(N__4765));
    LocalMux I__695 (
            .O(N__4765),
            .I(N__4762));
    Span4Mux_v I__694 (
            .O(N__4762),
            .I(N__4759));
    Sp12to4 I__693 (
            .O(N__4759),
            .I(N__4756));
    Span12Mux_h I__692 (
            .O(N__4756),
            .I(N__4753));
    Odrv12 I__691 (
            .O(N__4753),
            .I(A_c_12));
    InMux I__690 (
            .O(N__4750),
            .I(N__4747));
    LocalMux I__689 (
            .O(N__4747),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__688 (
            .O(N__4744),
            .I(N__4741));
    LocalMux I__687 (
            .O(N__4741),
            .I(N__4738));
    Odrv4 I__686 (
            .O(N__4738),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__685 (
            .O(N__4735),
            .I(N__4730));
    InMux I__684 (
            .O(N__4734),
            .I(N__4727));
    InMux I__683 (
            .O(N__4733),
            .I(N__4724));
    LocalMux I__682 (
            .O(N__4730),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__681 (
            .O(N__4727),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__680 (
            .O(N__4724),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    InMux I__679 (
            .O(N__4717),
            .I(N__4714));
    LocalMux I__678 (
            .O(N__4714),
            .I(N__4709));
    InMux I__677 (
            .O(N__4713),
            .I(N__4706));
    InMux I__676 (
            .O(N__4712),
            .I(N__4703));
    Odrv4 I__675 (
            .O(N__4709),
            .I(\U712_REG_SM.N_167_0 ));
    LocalMux I__674 (
            .O(N__4706),
            .I(\U712_REG_SM.N_167_0 ));
    LocalMux I__673 (
            .O(N__4703),
            .I(\U712_REG_SM.N_167_0 ));
    InMux I__672 (
            .O(N__4696),
            .I(N__4693));
    LocalMux I__671 (
            .O(N__4693),
            .I(N__4690));
    Span4Mux_h I__670 (
            .O(N__4690),
            .I(N__4687));
    Odrv4 I__669 (
            .O(N__4687),
            .I(\U712_REG_SM.N_117 ));
    InMux I__668 (
            .O(N__4684),
            .I(N__4681));
    LocalMux I__667 (
            .O(N__4681),
            .I(N__4677));
    CascadeMux I__666 (
            .O(N__4680),
            .I(N__4673));
    Span4Mux_v I__665 (
            .O(N__4677),
            .I(N__4670));
    InMux I__664 (
            .O(N__4676),
            .I(N__4667));
    InMux I__663 (
            .O(N__4673),
            .I(N__4664));
    Sp12to4 I__662 (
            .O(N__4670),
            .I(N__4659));
    LocalMux I__661 (
            .O(N__4667),
            .I(N__4659));
    LocalMux I__660 (
            .O(N__4664),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv12 I__659 (
            .O(N__4659),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    InMux I__658 (
            .O(N__4654),
            .I(N__4647));
    InMux I__657 (
            .O(N__4653),
            .I(N__4647));
    InMux I__656 (
            .O(N__4652),
            .I(N__4644));
    LocalMux I__655 (
            .O(N__4647),
            .I(N__4639));
    LocalMux I__654 (
            .O(N__4644),
            .I(N__4639));
    Sp12to4 I__653 (
            .O(N__4639),
            .I(N__4636));
    Span12Mux_v I__652 (
            .O(N__4636),
            .I(N__4633));
    Span12Mux_h I__651 (
            .O(N__4633),
            .I(N__4630));
    Odrv12 I__650 (
            .O(N__4630),
            .I(SIZ_c_0));
    InMux I__649 (
            .O(N__4627),
            .I(N__4624));
    LocalMux I__648 (
            .O(N__4624),
            .I(\U712_REG_SM.LDS_OUT_2_0_0 ));
    InMux I__647 (
            .O(N__4621),
            .I(N__4618));
    LocalMux I__646 (
            .O(N__4618),
            .I(\U712_REG_SM.UDS_OUT_2_0_0 ));
    IoInMux I__645 (
            .O(N__4615),
            .I(N__4612));
    LocalMux I__644 (
            .O(N__4612),
            .I(N__4609));
    Span12Mux_s0_v I__643 (
            .O(N__4609),
            .I(N__4606));
    Span12Mux_v I__642 (
            .O(N__4606),
            .I(N__4603));
    Odrv12 I__641 (
            .O(N__4603),
            .I(CMA_c_0));
    InMux I__640 (
            .O(N__4600),
            .I(N__4597));
    LocalMux I__639 (
            .O(N__4597),
            .I(\U712_CHIP_RAM.N_33 ));
    IoInMux I__638 (
            .O(N__4594),
            .I(N__4591));
    LocalMux I__637 (
            .O(N__4591),
            .I(N__4588));
    Span12Mux_s11_v I__636 (
            .O(N__4588),
            .I(N__4585));
    Odrv12 I__635 (
            .O(N__4585),
            .I(CMA_c_1));
    IoInMux I__634 (
            .O(N__4582),
            .I(N__4579));
    LocalMux I__633 (
            .O(N__4579),
            .I(N__4576));
    IoSpan4Mux I__632 (
            .O(N__4576),
            .I(N__4573));
    Sp12to4 I__631 (
            .O(N__4573),
            .I(N__4570));
    Span12Mux_s7_v I__630 (
            .O(N__4570),
            .I(N__4567));
    Odrv12 I__629 (
            .O(N__4567),
            .I(CMA_c_2));
    InMux I__628 (
            .O(N__4564),
            .I(N__4561));
    LocalMux I__627 (
            .O(N__4561),
            .I(N__4558));
    Span4Mux_v I__626 (
            .O(N__4558),
            .I(N__4555));
    Span4Mux_v I__625 (
            .O(N__4555),
            .I(N__4552));
    Sp12to4 I__624 (
            .O(N__4552),
            .I(N__4549));
    Span12Mux_h I__623 (
            .O(N__4549),
            .I(N__4546));
    Odrv12 I__622 (
            .O(N__4546),
            .I(A_c_4));
    CascadeMux I__621 (
            .O(N__4543),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_ ));
    InMux I__620 (
            .O(N__4540),
            .I(N__4537));
    LocalMux I__619 (
            .O(N__4537),
            .I(N__4534));
    Span12Mux_v I__618 (
            .O(N__4534),
            .I(N__4531));
    Span12Mux_h I__617 (
            .O(N__4531),
            .I(N__4528));
    Odrv12 I__616 (
            .O(N__4528),
            .I(A_c_11));
    InMux I__615 (
            .O(N__4525),
            .I(N__4522));
    LocalMux I__614 (
            .O(N__4522),
            .I(\U712_CHIP_RAM.N_34 ));
    InMux I__613 (
            .O(N__4519),
            .I(N__4516));
    LocalMux I__612 (
            .O(N__4516),
            .I(N__4513));
    Span4Mux_h I__611 (
            .O(N__4513),
            .I(N__4510));
    Span4Mux_v I__610 (
            .O(N__4510),
            .I(N__4507));
    Sp12to4 I__609 (
            .O(N__4507),
            .I(N__4504));
    Odrv12 I__608 (
            .O(N__4504),
            .I(A_c_7));
    CascadeMux I__607 (
            .O(N__4501),
            .I(N__4498));
    InMux I__606 (
            .O(N__4498),
            .I(N__4495));
    LocalMux I__605 (
            .O(N__4495),
            .I(N__4492));
    Span4Mux_v I__604 (
            .O(N__4492),
            .I(N__4489));
    Span4Mux_v I__603 (
            .O(N__4489),
            .I(N__4486));
    Sp12to4 I__602 (
            .O(N__4486),
            .I(N__4483));
    Span12Mux_h I__601 (
            .O(N__4483),
            .I(N__4480));
    Odrv12 I__600 (
            .O(N__4480),
            .I(A_c_14));
    CascadeMux I__599 (
            .O(N__4477),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa_1_cascade_ ));
    InMux I__598 (
            .O(N__4474),
            .I(N__4471));
    LocalMux I__597 (
            .O(N__4471),
            .I(N__4467));
    InMux I__596 (
            .O(N__4470),
            .I(N__4464));
    Odrv4 I__595 (
            .O(N__4467),
            .I(\U712_REG_SM.N_68 ));
    LocalMux I__594 (
            .O(N__4464),
            .I(\U712_REG_SM.N_68 ));
    CascadeMux I__593 (
            .O(N__4459),
            .I(\U712_REG_SM.N_188_cascade_ ));
    InMux I__592 (
            .O(N__4456),
            .I(N__4451));
    InMux I__591 (
            .O(N__4455),
            .I(N__4446));
    InMux I__590 (
            .O(N__4454),
            .I(N__4446));
    LocalMux I__589 (
            .O(N__4451),
            .I(\U712_REG_SM.N_162_0 ));
    LocalMux I__588 (
            .O(N__4446),
            .I(\U712_REG_SM.N_162_0 ));
    InMux I__587 (
            .O(N__4441),
            .I(N__4437));
    InMux I__586 (
            .O(N__4440),
            .I(N__4434));
    LocalMux I__585 (
            .O(N__4437),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__584 (
            .O(N__4434),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    IoInMux I__583 (
            .O(N__4429),
            .I(N__4425));
    IoInMux I__582 (
            .O(N__4428),
            .I(N__4422));
    LocalMux I__581 (
            .O(N__4425),
            .I(N__4419));
    LocalMux I__580 (
            .O(N__4422),
            .I(N__4416));
    IoSpan4Mux I__579 (
            .O(N__4419),
            .I(N__4413));
    IoSpan4Mux I__578 (
            .O(N__4416),
            .I(N__4410));
    Span4Mux_s1_v I__577 (
            .O(N__4413),
            .I(N__4407));
    Span4Mux_s1_v I__576 (
            .O(N__4410),
            .I(N__4404));
    Sp12to4 I__575 (
            .O(N__4407),
            .I(N__4401));
    Sp12to4 I__574 (
            .O(N__4404),
            .I(N__4398));
    Span12Mux_v I__573 (
            .O(N__4401),
            .I(N__4394));
    Span12Mux_v I__572 (
            .O(N__4398),
            .I(N__4391));
    InMux I__571 (
            .O(N__4397),
            .I(N__4388));
    Odrv12 I__570 (
            .O(N__4394),
            .I(ASn_c));
    Odrv12 I__569 (
            .O(N__4391),
            .I(ASn_c));
    LocalMux I__568 (
            .O(N__4388),
            .I(ASn_c));
    CascadeMux I__567 (
            .O(N__4381),
            .I(N__4378));
    InMux I__566 (
            .O(N__4378),
            .I(N__4372));
    InMux I__565 (
            .O(N__4377),
            .I(N__4372));
    LocalMux I__564 (
            .O(N__4372),
            .I(N__4369));
    Span4Mux_v I__563 (
            .O(N__4369),
            .I(N__4366));
    Span4Mux_v I__562 (
            .O(N__4366),
            .I(N__4363));
    Sp12to4 I__561 (
            .O(N__4363),
            .I(N__4360));
    Span12Mux_h I__560 (
            .O(N__4360),
            .I(N__4357));
    Odrv12 I__559 (
            .O(N__4357),
            .I(REGSPACEn_c));
    InMux I__558 (
            .O(N__4354),
            .I(N__4348));
    InMux I__557 (
            .O(N__4353),
            .I(N__4348));
    LocalMux I__556 (
            .O(N__4348),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa_1 ));
    InMux I__555 (
            .O(N__4345),
            .I(N__4336));
    InMux I__554 (
            .O(N__4344),
            .I(N__4336));
    InMux I__553 (
            .O(N__4343),
            .I(N__4336));
    LocalMux I__552 (
            .O(N__4336),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    CascadeMux I__551 (
            .O(N__4333),
            .I(N__4329));
    InMux I__550 (
            .O(N__4332),
            .I(N__4326));
    InMux I__549 (
            .O(N__4329),
            .I(N__4323));
    LocalMux I__548 (
            .O(N__4326),
            .I(N__4320));
    LocalMux I__547 (
            .O(N__4323),
            .I(N__4317));
    Span4Mux_v I__546 (
            .O(N__4320),
            .I(N__4311));
    Span4Mux_v I__545 (
            .O(N__4317),
            .I(N__4311));
    InMux I__544 (
            .O(N__4316),
            .I(N__4308));
    Sp12to4 I__543 (
            .O(N__4311),
            .I(N__4303));
    LocalMux I__542 (
            .O(N__4308),
            .I(N__4303));
    Span12Mux_h I__541 (
            .O(N__4303),
            .I(N__4300));
    Span12Mux_v I__540 (
            .O(N__4300),
            .I(N__4297));
    Odrv12 I__539 (
            .O(N__4297),
            .I(TSn_c));
    InMux I__538 (
            .O(N__4294),
            .I(N__4291));
    LocalMux I__537 (
            .O(N__4291),
            .I(N__4287));
    IoInMux I__536 (
            .O(N__4290),
            .I(N__4284));
    Span12Mux_h I__535 (
            .O(N__4287),
            .I(N__4281));
    LocalMux I__534 (
            .O(N__4284),
            .I(N__4278));
    Span12Mux_v I__533 (
            .O(N__4281),
            .I(N__4275));
    IoSpan4Mux I__532 (
            .O(N__4278),
            .I(N__4272));
    Odrv12 I__531 (
            .O(N__4275),
            .I(RAMENn_c));
    Odrv4 I__530 (
            .O(N__4272),
            .I(RAMENn_c));
    InMux I__529 (
            .O(N__4267),
            .I(N__4258));
    InMux I__528 (
            .O(N__4266),
            .I(N__4258));
    InMux I__527 (
            .O(N__4265),
            .I(N__4253));
    InMux I__526 (
            .O(N__4264),
            .I(N__4253));
    InMux I__525 (
            .O(N__4263),
            .I(N__4250));
    LocalMux I__524 (
            .O(N__4258),
            .I(\U712_REG_SM.N_171_0 ));
    LocalMux I__523 (
            .O(N__4253),
            .I(\U712_REG_SM.N_171_0 ));
    LocalMux I__522 (
            .O(N__4250),
            .I(\U712_REG_SM.N_171_0 ));
    InMux I__521 (
            .O(N__4243),
            .I(N__4236));
    InMux I__520 (
            .O(N__4242),
            .I(N__4229));
    InMux I__519 (
            .O(N__4241),
            .I(N__4229));
    InMux I__518 (
            .O(N__4240),
            .I(N__4229));
    InMux I__517 (
            .O(N__4239),
            .I(N__4226));
    LocalMux I__516 (
            .O(N__4236),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__515 (
            .O(N__4229),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__514 (
            .O(N__4226),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    CascadeMux I__513 (
            .O(N__4219),
            .I(\U712_REG_SM.N_165_0_cascade_ ));
    InMux I__512 (
            .O(N__4216),
            .I(N__4210));
    InMux I__511 (
            .O(N__4215),
            .I(N__4205));
    InMux I__510 (
            .O(N__4214),
            .I(N__4205));
    InMux I__509 (
            .O(N__4213),
            .I(N__4202));
    LocalMux I__508 (
            .O(N__4210),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    LocalMux I__507 (
            .O(N__4205),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    LocalMux I__506 (
            .O(N__4202),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    InMux I__505 (
            .O(N__4195),
            .I(N__4192));
    LocalMux I__504 (
            .O(N__4192),
            .I(\U712_CHIP_RAM.CPU_TACK_6 ));
    CascadeMux I__503 (
            .O(N__4189),
            .I(N__4185));
    InMux I__502 (
            .O(N__4188),
            .I(N__4179));
    InMux I__501 (
            .O(N__4185),
            .I(N__4179));
    InMux I__500 (
            .O(N__4184),
            .I(N__4176));
    LocalMux I__499 (
            .O(N__4179),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__498 (
            .O(N__4176),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__497 (
            .O(N__4171),
            .I(N__4167));
    InMux I__496 (
            .O(N__4170),
            .I(N__4164));
    LocalMux I__495 (
            .O(N__4167),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    LocalMux I__494 (
            .O(N__4164),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__493 (
            .O(N__4159),
            .I(N__4156));
    LocalMux I__492 (
            .O(N__4156),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0 ));
    InMux I__491 (
            .O(N__4153),
            .I(N__4150));
    LocalMux I__490 (
            .O(N__4150),
            .I(N__4147));
    Span12Mux_h I__489 (
            .O(N__4147),
            .I(N__4144));
    Span12Mux_v I__488 (
            .O(N__4144),
            .I(N__4141));
    Odrv12 I__487 (
            .O(N__4141),
            .I(A_c_3));
    CascadeMux I__486 (
            .O(N__4138),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_ ));
    InMux I__485 (
            .O(N__4135),
            .I(N__4132));
    LocalMux I__484 (
            .O(N__4132),
            .I(N__4129));
    Span4Mux_v I__483 (
            .O(N__4129),
            .I(N__4126));
    Sp12to4 I__482 (
            .O(N__4126),
            .I(N__4123));
    Span12Mux_h I__481 (
            .O(N__4123),
            .I(N__4120));
    Odrv12 I__480 (
            .O(N__4120),
            .I(A_c_10));
    InMux I__479 (
            .O(N__4117),
            .I(N__4114));
    LocalMux I__478 (
            .O(N__4114),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__477 (
            .O(N__4111),
            .I(N__4108));
    LocalMux I__476 (
            .O(N__4108),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_a3_0 ));
    CascadeMux I__475 (
            .O(N__4105),
            .I(N__4102));
    InMux I__474 (
            .O(N__4102),
            .I(N__4098));
    InMux I__473 (
            .O(N__4101),
            .I(N__4095));
    LocalMux I__472 (
            .O(N__4098),
            .I(CPU_TACKm));
    LocalMux I__471 (
            .O(N__4095),
            .I(CPU_TACKm));
    CascadeMux I__470 (
            .O(N__4090),
            .I(N__4087));
    InMux I__469 (
            .O(N__4087),
            .I(N__4084));
    LocalMux I__468 (
            .O(N__4084),
            .I(N__4079));
    InMux I__467 (
            .O(N__4083),
            .I(N__4074));
    InMux I__466 (
            .O(N__4082),
            .I(N__4074));
    Odrv12 I__465 (
            .O(N__4079),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    LocalMux I__464 (
            .O(N__4074),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    CascadeMux I__463 (
            .O(N__4069),
            .I(\U712_REG_SM.N_173_0_cascade_ ));
    InMux I__462 (
            .O(N__4066),
            .I(N__4061));
    InMux I__461 (
            .O(N__4065),
            .I(N__4056));
    InMux I__460 (
            .O(N__4064),
            .I(N__4056));
    LocalMux I__459 (
            .O(N__4061),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__458 (
            .O(N__4056),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    CascadeMux I__457 (
            .O(N__4051),
            .I(\U712_REG_SM.N_54_cascade_ ));
    InMux I__456 (
            .O(N__4048),
            .I(N__4045));
    LocalMux I__455 (
            .O(N__4045),
            .I(\U712_REG_SM.un1_STATE_COUNT_5_0_1 ));
    InMux I__454 (
            .O(N__4042),
            .I(N__4038));
    InMux I__453 (
            .O(N__4041),
            .I(N__4035));
    LocalMux I__452 (
            .O(N__4038),
            .I(REG_TACK));
    LocalMux I__451 (
            .O(N__4035),
            .I(REG_TACK));
    CascadeMux I__450 (
            .O(N__4030),
            .I(\U712_REG_SM.N_162_0_cascade_ ));
    InMux I__449 (
            .O(N__4027),
            .I(N__4024));
    LocalMux I__448 (
            .O(N__4024),
            .I(N__4014));
    InMux I__447 (
            .O(N__4023),
            .I(N__4009));
    InMux I__446 (
            .O(N__4022),
            .I(N__4009));
    InMux I__445 (
            .O(N__4021),
            .I(N__4006));
    InMux I__444 (
            .O(N__4020),
            .I(N__3999));
    InMux I__443 (
            .O(N__4019),
            .I(N__3999));
    InMux I__442 (
            .O(N__4018),
            .I(N__3999));
    InMux I__441 (
            .O(N__4017),
            .I(N__3996));
    Span4Mux_v I__440 (
            .O(N__4014),
            .I(N__3993));
    LocalMux I__439 (
            .O(N__4009),
            .I(N__3986));
    LocalMux I__438 (
            .O(N__4006),
            .I(N__3986));
    LocalMux I__437 (
            .O(N__3999),
            .I(N__3986));
    LocalMux I__436 (
            .O(N__3996),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    Odrv4 I__435 (
            .O(N__3993),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    Odrv4 I__434 (
            .O(N__3986),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__433 (
            .O(N__3979),
            .I(N__3971));
    InMux I__432 (
            .O(N__3978),
            .I(N__3971));
    InMux I__431 (
            .O(N__3977),
            .I(N__3968));
    InMux I__430 (
            .O(N__3976),
            .I(N__3965));
    LocalMux I__429 (
            .O(N__3971),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__428 (
            .O(N__3968),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__427 (
            .O(N__3965),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    CascadeMux I__426 (
            .O(N__3958),
            .I(N__3953));
    InMux I__425 (
            .O(N__3957),
            .I(N__3948));
    InMux I__424 (
            .O(N__3956),
            .I(N__3943));
    InMux I__423 (
            .O(N__3953),
            .I(N__3943));
    InMux I__422 (
            .O(N__3952),
            .I(N__3940));
    InMux I__421 (
            .O(N__3951),
            .I(N__3937));
    LocalMux I__420 (
            .O(N__3948),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__419 (
            .O(N__3943),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__418 (
            .O(N__3940),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__417 (
            .O(N__3937),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__416 (
            .O(N__3928),
            .I(N__3925));
    LocalMux I__415 (
            .O(N__3925),
            .I(N__3919));
    InMux I__414 (
            .O(N__3924),
            .I(N__3912));
    InMux I__413 (
            .O(N__3923),
            .I(N__3912));
    InMux I__412 (
            .O(N__3922),
            .I(N__3912));
    Span4Mux_v I__411 (
            .O(N__3919),
            .I(N__3909));
    LocalMux I__410 (
            .O(N__3912),
            .I(N__3906));
    Span4Mux_v I__409 (
            .O(N__3909),
            .I(N__3903));
    Span4Mux_h I__408 (
            .O(N__3906),
            .I(N__3900));
    Sp12to4 I__407 (
            .O(N__3903),
            .I(N__3897));
    Sp12to4 I__406 (
            .O(N__3900),
            .I(N__3894));
    Span12Mux_h I__405 (
            .O(N__3897),
            .I(N__3889));
    Span12Mux_v I__404 (
            .O(N__3894),
            .I(N__3889));
    Odrv12 I__403 (
            .O(N__3889),
            .I(CLK40_OUT_i));
    InMux I__402 (
            .O(N__3886),
            .I(N__3874));
    InMux I__401 (
            .O(N__3885),
            .I(N__3874));
    InMux I__400 (
            .O(N__3884),
            .I(N__3874));
    InMux I__399 (
            .O(N__3883),
            .I(N__3874));
    LocalMux I__398 (
            .O(N__3874),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__397 (
            .O(N__3871),
            .I(N__3866));
    InMux I__396 (
            .O(N__3870),
            .I(N__3863));
    InMux I__395 (
            .O(N__3869),
            .I(N__3860));
    LocalMux I__394 (
            .O(N__3866),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__393 (
            .O(N__3863),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__392 (
            .O(N__3860),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__391 (
            .O(N__3853),
            .I(N__3849));
    CascadeMux I__390 (
            .O(N__3852),
            .I(N__3846));
    InMux I__389 (
            .O(N__3849),
            .I(N__3843));
    InMux I__388 (
            .O(N__3846),
            .I(N__3840));
    LocalMux I__387 (
            .O(N__3843),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__386 (
            .O(N__3840),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__385 (
            .O(N__3835),
            .I(N__3829));
    InMux I__384 (
            .O(N__3834),
            .I(N__3826));
    InMux I__383 (
            .O(N__3833),
            .I(N__3823));
    InMux I__382 (
            .O(N__3832),
            .I(N__3818));
    InMux I__381 (
            .O(N__3829),
            .I(N__3818));
    LocalMux I__380 (
            .O(N__3826),
            .I(N__3813));
    LocalMux I__379 (
            .O(N__3823),
            .I(N__3813));
    LocalMux I__378 (
            .O(N__3818),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    Odrv4 I__377 (
            .O(N__3813),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CascadeMux I__376 (
            .O(N__3808),
            .I(\U712_CYCLE_TERM.N_45_0_0_en_cascade_ ));
    CEMux I__375 (
            .O(N__3805),
            .I(N__3802));
    LocalMux I__374 (
            .O(N__3802),
            .I(\U712_CYCLE_TERM.N_45_0_0_en_0 ));
    IoInMux I__373 (
            .O(N__3799),
            .I(N__3796));
    LocalMux I__372 (
            .O(N__3796),
            .I(N__3793));
    IoSpan4Mux I__371 (
            .O(N__3793),
            .I(N__3790));
    Span4Mux_s3_v I__370 (
            .O(N__3790),
            .I(N__3787));
    Sp12to4 I__369 (
            .O(N__3787),
            .I(N__3784));
    Odrv12 I__368 (
            .O(N__3784),
            .I(VBENn_c));
    CascadeMux I__367 (
            .O(N__3781),
            .I(N__3777));
    CascadeMux I__366 (
            .O(N__3780),
            .I(N__3774));
    InMux I__365 (
            .O(N__3777),
            .I(N__3770));
    InMux I__364 (
            .O(N__3774),
            .I(N__3767));
    InMux I__363 (
            .O(N__3773),
            .I(N__3764));
    LocalMux I__362 (
            .O(N__3770),
            .I(\U712_REG_SM.N_73 ));
    LocalMux I__361 (
            .O(N__3767),
            .I(\U712_REG_SM.N_73 ));
    LocalMux I__360 (
            .O(N__3764),
            .I(\U712_REG_SM.N_73 ));
    CascadeMux I__359 (
            .O(N__3757),
            .I(\U712_REG_SM.un1_STATE_COUNT_5_0_1_cascade_ ));
    InMux I__358 (
            .O(N__3754),
            .I(N__3750));
    InMux I__357 (
            .O(N__3753),
            .I(N__3747));
    LocalMux I__356 (
            .O(N__3750),
            .I(\U712_REG_SM.N_86 ));
    LocalMux I__355 (
            .O(N__3747),
            .I(\U712_REG_SM.N_86 ));
    CascadeMux I__354 (
            .O(N__3742),
            .I(\U712_REG_SM.N_68_cascade_ ));
    CascadeMux I__353 (
            .O(N__3739),
            .I(\U712_REG_SM.N_73_cascade_ ));
    IoInMux I__352 (
            .O(N__3736),
            .I(N__3733));
    LocalMux I__351 (
            .O(N__3733),
            .I(N__3730));
    IoSpan4Mux I__350 (
            .O(N__3730),
            .I(N__3727));
    Sp12to4 I__349 (
            .O(N__3727),
            .I(N__3724));
    Span12Mux_h I__348 (
            .O(N__3724),
            .I(N__3720));
    InMux I__347 (
            .O(N__3723),
            .I(N__3717));
    Odrv12 I__346 (
            .O(N__3720),
            .I(TACK_OUTn));
    LocalMux I__345 (
            .O(N__3717),
            .I(TACK_OUTn));
    IoInMux I__344 (
            .O(N__3712),
            .I(N__3708));
    InMux I__343 (
            .O(N__3711),
            .I(N__3705));
    LocalMux I__342 (
            .O(N__3708),
            .I(N__3702));
    LocalMux I__341 (
            .O(N__3705),
            .I(N__3699));
    Span4Mux_s3_h I__340 (
            .O(N__3702),
            .I(N__3696));
    Span12Mux_h I__339 (
            .O(N__3699),
            .I(N__3691));
    Sp12to4 I__338 (
            .O(N__3696),
            .I(N__3691));
    Span12Mux_v I__337 (
            .O(N__3691),
            .I(N__3688));
    Odrv12 I__336 (
            .O(N__3688),
            .I(C1_c));
    IoInMux I__335 (
            .O(N__3685),
            .I(N__3682));
    LocalMux I__334 (
            .O(N__3682),
            .I(N__3679));
    Span12Mux_s8_h I__333 (
            .O(N__3679),
            .I(N__3676));
    Odrv12 I__332 (
            .O(N__3676),
            .I(CLK40_OUT_i_i));
    InMux I__331 (
            .O(N__3673),
            .I(N__3670));
    LocalMux I__330 (
            .O(N__3670),
            .I(\U712_REG_SM.N_120 ));
    InMux I__329 (
            .O(N__3667),
            .I(N__3664));
    LocalMux I__328 (
            .O(N__3664),
            .I(N__3661));
    Span4Mux_v I__327 (
            .O(N__3661),
            .I(N__3658));
    Sp12to4 I__326 (
            .O(N__3658),
            .I(N__3655));
    Span12Mux_h I__325 (
            .O(N__3655),
            .I(N__3652));
    Odrv12 I__324 (
            .O(N__3652),
            .I(C3_c));
    IoInMux I__323 (
            .O(N__3649),
            .I(N__3646));
    LocalMux I__322 (
            .O(N__3646),
            .I(N__3643));
    Span4Mux_s2_h I__321 (
            .O(N__3643),
            .I(N__3640));
    Sp12to4 I__320 (
            .O(N__3640),
            .I(N__3637));
    Span12Mux_s11_v I__319 (
            .O(N__3637),
            .I(N__3634));
    Odrv12 I__318 (
            .O(N__3634),
            .I(N_677_i));
    InMux I__317 (
            .O(N__3631),
            .I(N__3628));
    LocalMux I__316 (
            .O(N__3628),
            .I(TACK_EN_i_ess));
    IoInMux I__315 (
            .O(N__3625),
            .I(N__3622));
    LocalMux I__314 (
            .O(N__3622),
            .I(N__3619));
    Span4Mux_s2_v I__313 (
            .O(N__3619),
            .I(N__3616));
    Span4Mux_v I__312 (
            .O(N__3616),
            .I(N__3613));
    Odrv4 I__311 (
            .O(N__3613),
            .I(CLK80_OUT_i_i));
    IoInMux I__310 (
            .O(N__3610),
            .I(N__3607));
    LocalMux I__309 (
            .O(N__3607),
            .I(N__3604));
    Span4Mux_s0_v I__308 (
            .O(N__3604),
            .I(N__3601));
    Span4Mux_v I__307 (
            .O(N__3601),
            .I(N__3598));
    Sp12to4 I__306 (
            .O(N__3598),
            .I(N__3595));
    Span12Mux_h I__305 (
            .O(N__3595),
            .I(N__3592));
    Span12Mux_v I__304 (
            .O(N__3592),
            .I(N__3589));
    Odrv12 I__303 (
            .O(N__3589),
            .I(CLK40_IN_c));
    defparam IN_MUX_bfv_14_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_4_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__4831),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__3712),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_2_1_7.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_2_1_7.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_2_1_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_2_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9577),
            .lcout(CLK80_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLK40C_obuf_RNO_LC_6_10_5.C_ON=1'b0;
    defparam CLK40C_obuf_RNO_LC_6_10_5.SEQ_MODE=4'b0000;
    defparam CLK40C_obuf_RNO_LC_6_10_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLK40C_obuf_RNO_LC_6_10_5 (
            .in0(N__3928),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_6_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_6_11_1 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_6_11_1  (
            .in0(N__4684),
            .in1(N__9158),
            .in2(N__4090),
            .in3(N__3673),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9569),
            .ce(),
            .sr(N__9366));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_11_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__4027),
            .in2(_gnd_net_),
            .in3(N__3753),
            .lcout(\U712_REG_SM.N_120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_0_LC_7_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_7_12_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_7_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3667),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9570),
            .ce(),
            .sr(N__9353));
    defparam TACKn_obuft_RNO_LC_7_15_4.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_7_15_4.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_7_15_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 TACKn_obuft_RNO_LC_7_15_4 (
            .in0(N__3631),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_677_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIVAPS2_3_LC_8_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIVAPS2_3_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIVAPS2_3_LC_8_12_5 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIVAPS2_3_LC_8_12_5  (
            .in0(N__3773),
            .in1(N__4929),
            .in2(N__4968),
            .in3(N__4676),
            .lcout(\U712_REG_SM.N_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_14_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_14_5 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_14_5 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_14_5  (
            .in0(N__3834),
            .in1(N__7816),
            .in2(_gnd_net_),
            .in3(N__3871),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9573),
            .ce(N__3805),
            .sr(N__9339));
    defparam \U712_REG_SM.C3_SYNC_2_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_2_LC_9_11_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_2_LC_9_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_2_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3957),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9555),
            .ce(),
            .sr(N__9349));
    defparam \U712_REG_SM.C1_SYNC_2_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_2_LC_9_11_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_2_LC_9_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_2_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4243),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9555),
            .ce(),
            .sr(N__9349));
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_11_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5044),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9555),
            .ce(),
            .sr(N__9349));
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_11_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_9_11_6  (
            .in0(N__4023),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9555),
            .ce(),
            .sr(N__9349));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_11_7 .LUT_INIT=16'b1011101110110000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_9_11_7  (
            .in0(N__4066),
            .in1(N__3754),
            .in2(N__3781),
            .in3(N__4022),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9555),
            .ce(),
            .sr(N__9349));
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_9_12_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__3976),
            .in2(_gnd_net_),
            .in3(N__3951),
            .lcout(\U712_REG_SM.N_68 ),
            .ltout(\U712_REG_SM.N_68_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI1FQR1_2_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI1FQR1_2_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI1FQR1_2_LC_9_12_2 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI1FQR1_2_LC_9_12_2  (
            .in0(N__5038),
            .in1(N__4213),
            .in2(N__3742),
            .in3(N__4239),
            .lcout(\U712_REG_SM.N_73 ),
            .ltout(\U712_REG_SM.N_73_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_12_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_12_3  (
            .in0(N__4969),
            .in1(N__4930),
            .in2(N__3739),
            .in3(N__4017),
            .lcout(\U712_REG_SM.N_117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_12_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_12_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_9_12_7  (
            .in0(N__4101),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4041),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_9_13_0  (
            .in0(N__4188),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9565),
            .ce(),
            .sr(N__9340));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_9_13_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_9_13_2 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_9_13_2 .LUT_INIT=16'b1111100011111100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_9_13_2  (
            .in0(N__3924),
            .in1(N__3723),
            .in2(N__4189),
            .in3(N__3885),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9565),
            .ce(),
            .sr(N__9340));
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_13_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3711),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9565),
            .ce(),
            .sr(N__9340));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_13_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_13_4 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_13_4 .LUT_INIT=16'b0011001000110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_9_13_4  (
            .in0(N__4159),
            .in1(N__3883),
            .in2(N__3853),
            .in3(N__3832),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9565),
            .ce(),
            .sr(N__9340));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_13_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4171),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9565),
            .ce(),
            .sr(N__9340));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_13_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_9_13_6  (
            .in0(N__3923),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3884),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9565),
            .ce(),
            .sr(N__9340));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_13_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_13_7 .LUT_INIT=16'b1010111110001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_9_13_7  (
            .in0(N__3886),
            .in1(N__3922),
            .in2(N__3835),
            .in3(N__3870),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9565),
            .ce(),
            .sr(N__9340));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_14_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_14_1 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_14_1  (
            .in0(N__7815),
            .in1(N__3869),
            .in2(N__3852),
            .in3(N__3833),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_45_0_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_14_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_14_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3808),
            .in3(N__9411),
            .lcout(\U712_CYCLE_TERM.N_45_0_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_LC_10_10_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_LC_10_10_2  (
            .in0(N__9173),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8116),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIFFKI2_4_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIFFKI2_4_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIFFKI2_4_LC_10_11_1 .LUT_INIT=16'b0011001100110001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIFFKI2_4_LC_10_11_1  (
            .in0(N__4065),
            .in1(N__4083),
            .in2(N__3780),
            .in3(N__4021),
            .lcout(\U712_REG_SM.un1_STATE_COUNT_5_0_1 ),
            .ltout(\U712_REG_SM.un1_STATE_COUNT_5_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_10_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_10_11_2 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_10_11_2  (
            .in0(N__3979),
            .in1(N__3956),
            .in2(N__3757),
            .in3(N__4455),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9550),
            .ce(),
            .sr(N__9344));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_10_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_10_11_4 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_10_11_4  (
            .in0(N__4111),
            .in1(N__8267),
            .in2(N__4105),
            .in3(N__4195),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9550),
            .ce(),
            .sr(N__9344));
    defparam \U712_REG_SM.STATE_COUNT_RNI1VLC2_5_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI1VLC2_5_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI1VLC2_5_LC_10_11_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI1VLC2_5_LC_10_11_5  (
            .in0(N__4454),
            .in1(N__3978),
            .in2(N__3958),
            .in3(N__4082),
            .lcout(\U712_REG_SM.N_173_0 ),
            .ltout(\U712_REG_SM.N_173_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_11_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(N__8189),
            .in2(N__4069),
            .in3(N__4064),
            .lcout(),
            .ltout(\U712_REG_SM.N_54_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_LC_10_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_10_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_10_11_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_10_11_7  (
            .in0(N__6415),
            .in1(N__4042),
            .in2(N__4051),
            .in3(N__4048),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9550),
            .ce(),
            .sr(N__9344));
    defparam \U712_REG_SM.C1_SYNC_RNIOEF21_2_LC_10_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIOEF21_2_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIOEF21_2_LC_10_12_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIOEF21_2_LC_10_12_0  (
            .in0(N__5036),
            .in1(N__4215),
            .in2(_gnd_net_),
            .in3(N__4240),
            .lcout(\U712_REG_SM.N_183_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_10_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_10_12_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(N__8179),
            .in2(_gnd_net_),
            .in3(N__4020),
            .lcout(\U712_REG_SM.RnW_m ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_12_2  (
            .in0(N__4018),
            .in1(N__4214),
            .in2(N__5043),
            .in3(N__4241),
            .lcout(\U712_REG_SM.N_162_0 ),
            .ltout(\U712_REG_SM.N_162_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_10_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_10_12_3 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__4440),
            .in2(N__4030),
            .in3(N__4470),
            .lcout(\U712_REG_SM.N_171_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIQU741_2_LC_10_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIQU741_2_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIQU741_2_LC_10_12_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIQU741_2_LC_10_12_4  (
            .in0(N__4019),
            .in1(N__3977),
            .in2(_gnd_net_),
            .in3(N__3952),
            .lcout(\U712_REG_SM.N_165_0 ),
            .ltout(\U712_REG_SM.N_165_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_10_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_10_12_5  (
            .in0(N__4242),
            .in1(N__5037),
            .in2(N__4219),
            .in3(N__4216),
            .lcout(\U712_REG_SM.N_167_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_12_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(N__8096),
            .in2(_gnd_net_),
            .in3(N__6981),
            .lcout(\U712_CHIP_RAM.CPU_TACK_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_13_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_13_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__4184),
            .in2(_gnd_net_),
            .in3(N__4170),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_7_1 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_7_1  (
            .in0(N__4117),
            .in1(N__8104),
            .in2(N__8702),
            .in3(N__6001),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_2 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_2  (
            .in0(N__8105),
            .in1(N__4153),
            .in2(N__4138),
            .in3(N__4135),
            .lcout(\U712_CHIP_RAM.N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_11_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_11_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5152),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9526),
            .ce(N__8953),
            .sr(N__9354));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_11_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_11_11_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__6387),
            .in2(_gnd_net_),
            .in3(N__6863),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_11_5 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_11_5  (
            .in0(N__6864),
            .in1(N__6982),
            .in2(N__7894),
            .in3(N__8349),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_11_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_11_11_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_11_11_6  (
            .in0(N__6411),
            .in1(N__6450),
            .in2(_gnd_net_),
            .in3(N__6426),
            .lcout(\U712_REG_SM.DS_EN_0_sqmuxa_1 ),
            .ltout(\U712_REG_SM.DS_EN_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_11_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_11_11_7 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_1_LC_11_11_7  (
            .in0(N__4733),
            .in1(N__4712),
            .in2(N__4477),
            .in3(N__4263),
            .lcout(\U712_REG_SM.un1_LDS_OUT_0_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_12_0 .LUT_INIT=16'b0000000011111011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_12_0  (
            .in0(N__4332),
            .in1(N__4343),
            .in2(N__4381),
            .in3(N__4441),
            .lcout(),
            .ltout(\U712_REG_SM.N_188_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_12_1 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_11_12_1  (
            .in0(N__4345),
            .in1(N__4474),
            .in2(N__4459),
            .in3(N__4456),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9551),
            .ce(),
            .sr(N__9329));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_11_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_11_12_3 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_11_12_3  (
            .in0(N__4734),
            .in1(N__4713),
            .in2(_gnd_net_),
            .in3(N__4264),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9551),
            .ce(),
            .sr(N__9329));
    defparam \U712_REG_SM.REGENn_1_LC_11_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_1_LC_11_12_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_1_LC_11_12_5 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_REG_SM.REGENn_1_LC_11_12_5  (
            .in0(N__4397),
            .in1(N__4353),
            .in2(_gnd_net_),
            .in3(N__4265),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9551),
            .ce(),
            .sr(N__9329));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_12_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_12_7 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_11_12_7  (
            .in0(N__4344),
            .in1(N__4377),
            .in2(N__4333),
            .in3(N__4354),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9551),
            .ce(),
            .sr(N__9329));
    defparam \U712_REG_SM.UDS_OUT_LC_11_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.UDS_OUT_LC_11_13_2 .LUT_INIT=16'b0111011111110000;
    LogicCell40 \U712_REG_SM.UDS_OUT_LC_11_13_2  (
            .in0(N__4654),
            .in1(N__4621),
            .in2(N__4869),
            .in3(N__4266),
            .lcout(\U712_REG_SM.UDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9556),
            .ce(),
            .sr(N__9322));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_13_3 .LUT_INIT=16'b0001000111110001;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_13_3  (
            .in0(N__4316),
            .in1(N__4294),
            .in2(N__5062),
            .in3(N__8075),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9556),
            .ce(),
            .sr(N__9322));
    defparam \U712_REG_SM.LDS_OUT_LC_11_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.LDS_OUT_LC_11_13_5 .LUT_INIT=16'b0111001011111010;
    LogicCell40 \U712_REG_SM.LDS_OUT_LC_11_13_5  (
            .in0(N__4267),
            .in1(N__4627),
            .in2(N__6288),
            .in3(N__4653),
            .lcout(\U712_REG_SM.LDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9556),
            .ce(),
            .sr(N__9322));
    defparam \U712_BYTE_ENABLE.LW_TRANS_LC_11_14_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LW_TRANS_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LW_TRANS_LC_11_14_1 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \U712_BYTE_ENABLE.LW_TRANS_LC_11_14_1  (
            .in0(N__4652),
            .in1(N__4902),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_BYTE_ENABLE.LW_TRANS_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDS_OUT_RNO_0_LC_11_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_RNO_0_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_RNO_0_LC_11_14_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_REG_SM.LDS_OUT_RNO_0_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__5475),
            .in2(_gnd_net_),
            .in3(N__8163),
            .lcout(\U712_REG_SM.LDS_OUT_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDS_OUT_RNO_0_LC_11_14_3 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_RNO_0_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDS_OUT_RNO_0_LC_11_14_3 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \U712_REG_SM.UDS_OUT_RNO_0_LC_11_14_3  (
            .in0(N__5476),
            .in1(_gnd_net_),
            .in2(N__8178),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.UDS_OUT_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_7_2 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_12_7_2  (
            .in0(N__5221),
            .in1(_gnd_net_),
            .in2(N__8821),
            .in3(N__8530),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9522),
            .ce(N__7395),
            .sr(N__9352));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_3 .LUT_INIT=16'b1010101010100011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_7_3  (
            .in0(N__4600),
            .in1(N__8691),
            .in2(N__8539),
            .in3(N__8812),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9522),
            .ce(N__7395),
            .sr(N__9352));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_7_7 .LUT_INIT=16'b1111110000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(N__8811),
            .in2(N__8540),
            .in3(N__4525),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9522),
            .ce(N__7395),
            .sr(N__9352));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_8_1 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_8_1  (
            .in0(N__8695),
            .in1(N__4744),
            .in2(N__8121),
            .in3(N__5113),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_2 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_2  (
            .in0(N__8092),
            .in1(N__4564),
            .in2(N__4543),
            .in3(N__4540),
            .lcout(\U712_CHIP_RAM.N_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_8_3 .LUT_INIT=16'b1101100001010101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_8_3  (
            .in0(N__5095),
            .in1(N__4519),
            .in2(N__4501),
            .in3(N__8090),
            .lcout(\U712_CHIP_RAM.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_6 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_6  (
            .in0(N__8089),
            .in1(N__6565),
            .in2(N__8699),
            .in3(N__5107),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_8_7 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_8_7  (
            .in0(N__4822),
            .in1(N__4807),
            .in2(N__4789),
            .in3(N__8091),
            .lcout(\U712_CHIP_RAM.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_12_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_12_9_4 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_12_9_4  (
            .in0(N__4750),
            .in1(N__8065),
            .in2(N__8703),
            .in3(N__5158),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_9_5 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_9_5  (
            .in0(N__8066),
            .in1(N__4786),
            .in2(N__4771),
            .in3(N__4768),
            .lcout(\U712_CHIP_RAM.N_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6549),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9530),
            .ce(N__8935),
            .sr(N__9338));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_10_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_10_4  (
            .in0(N__5184),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9530),
            .ce(N__8935),
            .sr(N__9338));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_12_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_12_11_2 .LUT_INIT=16'b0101011100000010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_12_11_2  (
            .in0(N__5617),
            .in1(N__6388),
            .in2(N__6873),
            .in3(N__8024),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9534),
            .ce(),
            .sr(N__9328));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_12_1 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_12_12_1  (
            .in0(N__4735),
            .in1(N__4717),
            .in2(N__4680),
            .in3(N__4696),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9544),
            .ce(),
            .sr(N__9321));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_12_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_12_12_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_12_12_3  (
            .in0(N__4917),
            .in1(N__4948),
            .in2(_gnd_net_),
            .in3(N__5055),
            .lcout(\U712_CHIP_RAM.un1_DBR_SYNC ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_LC_12_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_12_12_7 .LUT_INIT=16'b1010101011111100;
    LogicCell40 \U712_REG_SM.DS_EN_LC_12_12_7  (
            .in0(N__6305),
            .in1(N__5039),
            .in2(N__5002),
            .in3(N__4990),
            .lcout(\U712_REG_SM.DS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9544),
            .ce(),
            .sr(N__9321));
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_12_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_12_13_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_12_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DBR_SYNC_0_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4984),
            .lcout(U712_REG_SM_DBR_SYNC_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9549),
            .ce(),
            .sr(N__9320));
    defparam \U712_REG_SM.DBR_SYNC_1_LC_12_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_12_13_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_12_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_1_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4955),
            .lcout(U712_REG_SM_DBR_SYNC_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9549),
            .ce(),
            .sr(N__9320));
    defparam \U712_BYTE_ENABLE.LLBE_0_tz_LC_12_14_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_0_tz_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_0_tz_LC_12_14_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_0_tz_LC_12_14_6  (
            .in0(N__5477),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4906),
            .lcout(\U712_BYTE_ENABLE.LLBE_0_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_12_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_12_15_7 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_REG_SM.UDS_OUT_RNIUP9B_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__4870),
            .in2(_gnd_net_),
            .in3(N__6312),
            .lcout(U712_REG_SM_un1_UDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_2.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_2.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7780),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_13_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_13_4_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_13_4_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_13_4_1  (
            .in0(_gnd_net_),
            .in1(N__5643),
            .in2(_gnd_net_),
            .in3(N__5658),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_13_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_13_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_13_4_5 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_13_4_5  (
            .in0(N__5694),
            .in1(N__5709),
            .in2(N__5677),
            .in3(N__5724),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_7_1 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_7_1  (
            .in0(N__8680),
            .in1(N__5827),
            .in2(N__8122),
            .in3(N__5992),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_2  (
            .in0(N__8103),
            .in1(N__5263),
            .in2(N__5245),
            .in3(N__5242),
            .lcout(\U712_CHIP_RAM.N_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_7_7 .LUT_INIT=16'b1010100010101011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_13_7_7  (
            .in0(N__5215),
            .in1(N__8816),
            .in2(N__8541),
            .in3(N__8690),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9524),
            .ce(N__7394),
            .sr(N__9363));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_0  (
            .in0(N__5185),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9527),
            .ce(N__9064),
            .sr(N__9355));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5148),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9527),
            .ce(N__9064),
            .sr(N__9355));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5818),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9527),
            .ce(N__9064),
            .sr(N__9355));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_8_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_8_7  (
            .in0(N__5089),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9527),
            .ce(N__9064),
            .sr(N__9355));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_9_1 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_9_1  (
            .in0(N__8644),
            .in1(N__5794),
            .in2(N__8088),
            .in3(N__5101),
            .lcout(\U712_CHIP_RAM.CMA_5_3_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_13_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_13_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5088),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9531),
            .ce(N__8945),
            .sr(N__9350));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_10_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_13_10_3  (
            .in0(N__5374),
            .in1(N__8769),
            .in2(_gnd_net_),
            .in3(N__8511),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9538),
            .ce(N__7396),
            .sr(N__9345));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_10_5 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_10_5  (
            .in0(N__5347),
            .in1(N__6088),
            .in2(N__5329),
            .in3(N__8023),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_36_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_10_6 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__8768),
            .in2(N__5305),
            .in3(N__8510),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9538),
            .ce(N__7396),
            .sr(N__9345));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_13_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_13_11_0 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_13_11_0  (
            .in0(N__6069),
            .in1(N__5281),
            .in2(N__6055),
            .in3(N__7193),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9545),
            .ce(N__6123),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_13_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_13_11_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_13_11_1  (
            .in0(N__5404),
            .in1(N__7798),
            .in2(_gnd_net_),
            .in3(N__7236),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_13_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_13_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_13_11_2  (
            .in0(N__7014),
            .in1(N__7060),
            .in2(N__7089),
            .in3(N__7111),
            .lcout(\U712_CHIP_RAM.N_61 ),
            .ltout(\U712_CHIP_RAM.N_61_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_13_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_13_11_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5275),
            .in3(N__7855),
            .lcout(\U712_CHIP_RAM.N_65 ),
            .ltout(\U712_CHIP_RAM.N_65_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_13_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_13_11_4 .LUT_INIT=16'b0101010101011101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_13_11_4  (
            .in0(N__7799),
            .in1(N__5269),
            .in2(N__5272),
            .in3(N__7701),
            .lcout(\U712_CHIP_RAM.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_1_LC_13_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_1_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_1_LC_13_11_5 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_1_LC_13_11_5  (
            .in0(N__6847),
            .in1(_gnd_net_),
            .in2(N__6976),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_104_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI399Q7_LC_13_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI399Q7_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI399Q7_LC_13_11_6 .LUT_INIT=16'b0101000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI399Q7_LC_13_11_6  (
            .in0(N__7251),
            .in1(N__7192),
            .in2(N__6019),
            .in3(N__7702),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER16_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIEBLDE_LC_13_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIEBLDE_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIEBLDE_LC_13_11_7 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIEBLDE_LC_13_11_7  (
            .in0(N__5403),
            .in1(N__8218),
            .in2(N__5392),
            .in3(N__6081),
            .lcout(\U712_CHIP_RAM.N_158_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_13_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_13_12_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_13_12_0  (
            .in0(N__8350),
            .in1(N__7576),
            .in2(N__6874),
            .in3(N__8251),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_0_LC_13_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_0_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_0_LC_13_12_1 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_0_LC_13_12_1  (
            .in0(N__6504),
            .in1(_gnd_net_),
            .in2(N__5389),
            .in3(N__7197),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_13_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_13_12_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5386),
            .in3(N__9410),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI3EN62_0_LC_13_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI3EN62_0_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI3EN62_0_LC_13_12_3 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI3EN62_0_LC_13_12_3  (
            .in0(N__6380),
            .in1(N__7706),
            .in2(N__7630),
            .in3(N__6336),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_1_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_13_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_13_12_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_13_12_4  (
            .in0(N__6868),
            .in1(N__8250),
            .in2(N__6977),
            .in3(N__7853),
            .lcout(\U712_CHIP_RAM.N_67 ),
            .ltout(\U712_CHIP_RAM.N_67_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFQROA_LC_13_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFQROA_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFQROA_LC_13_12_5 .LUT_INIT=16'b0000010000110111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFQROA_LC_13_12_5  (
            .in0(N__7628),
            .in1(N__7707),
            .in2(N__5383),
            .in3(N__6103),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER18_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER18_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_13_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_13_12_6 .LUT_INIT=16'b0000001000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_13_12_6  (
            .in0(N__7198),
            .in1(N__6082),
            .in2(N__5380),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_m2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_13_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_13_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_13_12_7 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_13_12_7  (
            .in0(N__7808),
            .in1(_gnd_net_),
            .in2(N__5377),
            .in3(N__6053),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9552),
            .ce(N__6124),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_13_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_13_13_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_13_13_6 .LUT_INIT=16'b0010111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_13_13_6  (
            .in0(N__5768),
            .in1(N__5616),
            .in2(N__8968),
            .in3(N__5605),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9557),
            .ce(),
            .sr(N__9323));
    defparam \U712_BYTE_ENABLE.un2_CUMBEn_LC_13_14_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un2_CUMBEn_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un2_CUMBEn_LC_13_14_0 .LUT_INIT=16'b0001111100000000;
    LogicCell40 \U712_BYTE_ENABLE.un2_CUMBEn_LC_13_14_0  (
            .in0(N__5508),
            .in1(N__5566),
            .in2(N__5436),
            .in3(N__8119),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.un2_CUMBEnZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_LC_13_14_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_LC_13_14_1 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_LC_13_14_1  (
            .in0(N__9125),
            .in1(N__6744),
            .in2(N__5593),
            .in3(N__5771),
            .lcout(CUMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un2_CLLBEn_LC_13_14_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un2_CLLBEn_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un2_CLLBEn_LC_13_14_2 .LUT_INIT=16'b0010111100000000;
    LogicCell40 \U712_BYTE_ENABLE.un2_CLLBEn_LC_13_14_2  (
            .in0(N__5506),
            .in1(N__5565),
            .in2(N__5434),
            .in3(N__8117),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.un2_CLLBEnZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_LC_13_14_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_LC_13_14_3 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_LC_13_14_3  (
            .in0(N__9123),
            .in1(N__6743),
            .in2(N__5557),
            .in3(N__5769),
            .lcout(CLLBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un2_CLMBEn_LC_13_14_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un2_CLMBEn_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un2_CLMBEn_LC_13_14_4 .LUT_INIT=16'b0010111100000000;
    LogicCell40 \U712_BYTE_ENABLE.un2_CLMBEn_LC_13_14_4  (
            .in0(N__5507),
            .in1(N__5478),
            .in2(N__5435),
            .in3(N__8118),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.un2_CLMBEnZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_LC_13_14_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_LC_13_14_5 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_LC_13_14_5  (
            .in0(N__9124),
            .in1(N__6702),
            .in2(N__5533),
            .in3(N__5770),
            .lcout(CLMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un2_CUUBEn_LC_13_14_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un2_CUUBEn_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un2_CUUBEn_LC_13_14_6 .LUT_INIT=16'b0001111100000000;
    LogicCell40 \U712_BYTE_ENABLE.un2_CUUBEn_LC_13_14_6  (
            .in0(N__5509),
            .in1(N__5479),
            .in2(N__5437),
            .in3(N__8120),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.un2_CUUBEnZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_LC_13_14_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_LC_13_14_7 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_LC_13_14_7  (
            .in0(N__9126),
            .in1(N__6703),
            .in2(N__5407),
            .in3(N__5772),
            .lcout(CUUBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_14_4_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_14_4_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_14_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_14_4_0  (
            .in0(_gnd_net_),
            .in1(N__5725),
            .in2(_gnd_net_),
            .in3(N__5713),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_4_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__5626),
            .ce(),
            .sr(N__6010));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_14_4_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_14_4_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_14_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_14_4_1  (
            .in0(_gnd_net_),
            .in1(N__5710),
            .in2(_gnd_net_),
            .in3(N__5698),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__5626),
            .ce(),
            .sr(N__6010));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_14_4_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_14_4_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_14_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_14_4_2  (
            .in0(_gnd_net_),
            .in1(N__5695),
            .in2(_gnd_net_),
            .in3(N__5683),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__5626),
            .ce(),
            .sr(N__6010));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_14_4_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_14_4_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_14_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_14_4_3  (
            .in0(_gnd_net_),
            .in1(N__6241),
            .in2(_gnd_net_),
            .in3(N__5680),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__5626),
            .ce(),
            .sr(N__6010));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_14_4_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_14_4_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_14_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_14_4_4  (
            .in0(_gnd_net_),
            .in1(N__5676),
            .in2(_gnd_net_),
            .in3(N__5662),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__5626),
            .ce(),
            .sr(N__6010));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_14_4_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_14_4_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_14_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_14_4_5  (
            .in0(_gnd_net_),
            .in1(N__5659),
            .in2(_gnd_net_),
            .in3(N__5647),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__5626),
            .ce(),
            .sr(N__6010));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_14_4_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_14_4_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_14_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_14_4_6  (
            .in0(_gnd_net_),
            .in1(N__5644),
            .in2(_gnd_net_),
            .in3(N__5632),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__5626),
            .ce(),
            .sr(N__6010));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_14_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_14_4_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_14_4_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_14_4_7  (
            .in0(_gnd_net_),
            .in1(N__6228),
            .in2(_gnd_net_),
            .in3(N__5629),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5626),
            .ce(),
            .sr(N__6010));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_14_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_14_5_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_14_5_0  (
            .in0(N__8676),
            .in1(N__8515),
            .in2(N__8817),
            .in3(N__8879),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_7_1  (
            .in0(N__5860),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9528),
            .ce(N__9063),
            .sr(N__9367));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9007),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9528),
            .ce(N__9063),
            .sr(N__9367));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_2_LC_14_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_2_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_2_LC_14_8_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_2_LC_14_8_3  (
            .in0(N__8800),
            .in1(N__8663),
            .in2(_gnd_net_),
            .in3(N__8516),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(\U712_CHIP_RAM.CMA_5_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_8_4 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_14_8_4  (
            .in0(N__7264),
            .in1(N__5986),
            .in2(N__5965),
            .in3(N__8097),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9532),
            .ce(N__7392),
            .sr(N__9364));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_8_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_14_8_5  (
            .in0(N__8801),
            .in1(N__5941),
            .in2(_gnd_net_),
            .in3(N__8517),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9532),
            .ce(N__7392),
            .sr(N__9364));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_8_6 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_14_8_6  (
            .in0(N__8407),
            .in1(N__5911),
            .in2(N__5905),
            .in3(N__8098),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9532),
            .ce(N__7392),
            .sr(N__9364));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_14_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_14_9_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_14_9_1  (
            .in0(N__5856),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9539),
            .ce(N__8920),
            .sr(N__9356));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_14_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_14_9_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_14_9_7  (
            .in0(N__5814),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9539),
            .ce(N__8920),
            .sr(N__9356));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_14_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_14_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_14_10_1 .LUT_INIT=16'b1111110100110001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_14_10_1  (
            .in0(N__7795),
            .in1(N__6610),
            .in2(N__6054),
            .in3(N__8468),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9546),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_14_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_14_10_3 .LUT_INIT=16'b0001001000010011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_14_10_3  (
            .in0(N__8615),
            .in1(N__8866),
            .in2(N__8781),
            .in3(N__8467),
            .lcout(\U712_CHIP_RAM.un1_CMA31_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_10_6 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_10_6  (
            .in0(N__6517),
            .in1(N__8109),
            .in2(N__6097),
            .in3(N__8616),
            .lcout(\U712_CHIP_RAM.CMA_5_3_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_14_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_14_11_0 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_14_11_0  (
            .in0(N__6807),
            .in1(_gnd_net_),
            .in2(N__6975),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITC5T1_1_LC_14_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITC5T1_1_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITC5T1_1_LC_14_11_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITC5T1_1_LC_14_11_1  (
            .in0(N__6846),
            .in1(N__6954),
            .in2(_gnd_net_),
            .in3(N__8348),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_14_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_14_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_14_11_2 .LUT_INIT=16'b0000001101010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_14_11_2  (
            .in0(N__6025),
            .in1(N__6070),
            .in2(N__6058),
            .in3(N__6049),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9553),
            .ce(N__6601),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_14_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_14_11_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_14_11_3  (
            .in0(N__7753),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7235),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_1_LC_14_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_1_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_1_LC_14_11_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_1_LC_14_11_4  (
            .in0(N__6806),
            .in1(_gnd_net_),
            .in2(N__6974),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_2_1_LC_14_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_2_1_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_2_1_LC_14_11_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_2_1_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(N__6804),
            .in2(_gnd_net_),
            .in3(N__6947),
            .lcout(\U712_CHIP_RAM.N_124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_14_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_14_11_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_14_11_6  (
            .in0(N__6805),
            .in1(N__7754),
            .in2(_gnd_net_),
            .in3(N__8249),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_0 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIO007I_0_0_LC_14_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIO007I_0_0_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIO007I_0_0_LC_14_11_7 .LUT_INIT=16'b0000010100010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIO007I_0_0_LC_14_11_7  (
            .in0(N__6625),
            .in1(N__8323),
            .in2(N__6127),
            .in3(N__8299),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_14_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_14_12_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_14_12_0  (
            .in0(N__6990),
            .in1(N__7041),
            .in2(N__6862),
            .in3(N__7523),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_5 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI971H6_2_LC_14_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI971H6_2_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI971H6_2_LC_14_12_1 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI971H6_2_LC_14_12_1  (
            .in0(N__7042),
            .in1(N__7033),
            .in2(N__6106),
            .in3(N__6991),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2VVR2_LC_14_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2VVR2_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2VVR2_LC_14_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2VVR2_LC_14_12_2  (
            .in0(N__7796),
            .in1(N__8248),
            .in2(N__7708),
            .in3(N__7609),
            .lcout(\U712_CHIP_RAM.N_108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_14_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_14_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_14_12_3 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_14_12_3  (
            .in0(N__6586),
            .in1(N__9413),
            .in2(N__7026),
            .in3(N__7116),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9558),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_14_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_14_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_14_12_4 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_14_12_4  (
            .in0(N__6837),
            .in1(N__6973),
            .in2(_gnd_net_),
            .in3(N__6885),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9558),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_14_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_14_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_14_12_5 .LUT_INIT=16'b0001001000010010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_14_12_5  (
            .in0(N__6585),
            .in1(N__9412),
            .in2(N__7027),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9558),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_14_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_14_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_14_12_6 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_14_12_6  (
            .in0(N__9415),
            .in1(N__6487),
            .in2(N__7066),
            .in3(N__7088),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9558),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_14_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_14_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_14_12_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_14_12_7  (
            .in0(N__6486),
            .in1(N__9414),
            .in2(_gnd_net_),
            .in3(N__7065),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9558),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_14_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_14_13_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_14_13_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__6378),
            .in2(_gnd_net_),
            .in3(N__6861),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9561),
            .ce(N__6322),
            .sr(N__9330));
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_14_14_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_14_14_0 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_14_14_0  (
            .in0(N__9409),
            .in1(N__6651),
            .in2(_gnd_net_),
            .in3(N__6665),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_14_14_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_14_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_14_14_3 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_14_14_3  (
            .in0(N__6652),
            .in1(N__9122),
            .in2(N__6670),
            .in3(N__6377),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9566),
            .ce(),
            .sr(N__9324));
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_14_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_14_15_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_REG_SM.LDS_OUT_RNIL31J_LC_14_15_0  (
            .in0(N__6316),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6292),
            .lcout(U712_REG_SM_un1_LDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_15_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_15_4_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_15_4_7 .LUT_INIT=16'b1111010111111101;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_15_4_7  (
            .in0(N__6250),
            .in1(N__6240),
            .in2(N__6229),
            .in3(N__6214),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9523),
            .ce(),
            .sr(N__9376));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_5_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_15_5_7  (
            .in0(N__6139),
            .in1(N__8820),
            .in2(_gnd_net_),
            .in3(N__8534),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9525),
            .ce(N__7379),
            .sr(N__9374));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_6_2 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_6_2  (
            .in0(N__6184),
            .in1(N__6133),
            .in2(N__6163),
            .in3(N__8123),
            .lcout(\U712_CHIP_RAM.N_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_15_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_15_7_2 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_15_7_2  (
            .in0(N__6556),
            .in1(N__8099),
            .in2(N__8700),
            .in3(N__7303),
            .lcout(\U712_CHIP_RAM.CMA_5_3_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_15_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_15_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_15_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7330),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9540),
            .ce(N__8952),
            .sr(N__9368));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_15_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_15_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_15_8_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_15_8_4  (
            .in0(N__7297),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9540),
            .ce(N__8952),
            .sr(N__9368));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6550),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9547),
            .ce(N__9059),
            .sr(N__9365));
    defparam \U712_CHIP_RAM.DBDIR_LC_15_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_15_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_15_10_0 .LUT_INIT=16'b1111000001110100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_15_10_0  (
            .in0(N__7933),
            .in1(N__6511),
            .in2(N__7460),
            .in3(N__7219),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9554),
            .ce(),
            .sr(N__9357));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_15_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_15_10_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_15_10_4  (
            .in0(N__9417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6493),
            .lcout(\U712_CHIP_RAM.un1_CMA31_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_15_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_15_10_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_15_10_5  (
            .in0(N__7117),
            .in1(N__7025),
            .in2(_gnd_net_),
            .in3(N__6584),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_15_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_15_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_15_10_6 .LUT_INIT=16'b0011111100101010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_15_10_6  (
            .in0(N__6475),
            .in1(N__6460),
            .in2(N__6439),
            .in3(N__6404),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9554),
            .ce(),
            .sr(N__9357));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG7JB2_1_LC_15_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG7JB2_1_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG7JB2_1_LC_15_11_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIG7JB2_1_LC_15_11_0  (
            .in0(N__7839),
            .in1(N__7752),
            .in2(N__6853),
            .in3(N__6957),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI3EN62_LC_15_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI3EN62_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI3EN62_LC_15_11_1 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI3EN62_LC_15_11_1  (
            .in0(N__6379),
            .in1(N__7615),
            .in2(N__6343),
            .in3(N__7684),
            .lcout(\U712_CHIP_RAM.N_77 ),
            .ltout(\U712_CHIP_RAM.N_77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4B3NB_LC_15_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4B3NB_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4B3NB_LC_15_11_2 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4B3NB_LC_15_11_2  (
            .in0(N__6643),
            .in1(N__6637),
            .in2(N__6628),
            .in3(N__7483),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIO007I_0_LC_15_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIO007I_0_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIO007I_0_LC_15_11_3 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIO007I_0_LC_15_11_3  (
            .in0(N__6619),
            .in1(N__8322),
            .in2(N__6613),
            .in3(N__8298),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_15_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_15_11_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6604),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_15_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_15_11_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_15_11_5  (
            .in0(N__6833),
            .in1(N__7570),
            .in2(_gnd_net_),
            .in3(N__7522),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_15_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_15_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_15_11_6 .LUT_INIT=16'b0001001100010010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_15_11_6  (
            .in0(N__7217),
            .in1(N__6571),
            .in2(N__6854),
            .in3(N__7135),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9559),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_15_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_15_11_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_15_11_7  (
            .in0(N__6958),
            .in1(N__7840),
            .in2(N__7624),
            .in3(N__7683),
            .lcout(\U712_CHIP_RAM.N_121 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_15_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_15_12_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__8363),
            .in2(_gnd_net_),
            .in3(N__8376),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_2_LC_15_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_2_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_2_LC_15_12_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_2_LC_15_12_1  (
            .in0(N__6956),
            .in1(N__7882),
            .in2(N__7525),
            .in3(N__7682),
            .lcout(\U712_CHIP_RAM.N_122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJ42D8_0_LC_15_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJ42D8_0_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJ42D8_0_LC_15_12_2 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIJ42D8_0_LC_15_12_2  (
            .in0(N__6856),
            .in1(N__9416),
            .in2(N__8272),
            .in3(N__8281),
            .lcout(\U712_CHIP_RAM.N_80 ),
            .ltout(\U712_CHIP_RAM.N_80_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQU7BE_0_LC_15_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQU7BE_0_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQU7BE_0_LC_15_12_3 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQU7BE_0_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(N__7134),
            .in2(N__7123),
            .in3(N__7207),
            .lcout(\U712_CHIP_RAM.N_50 ),
            .ltout(\U712_CHIP_RAM.N_50_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_15_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_15_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_15_12_4 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_15_12_4  (
            .in0(N__6857),
            .in1(N__7521),
            .in2(N__7120),
            .in3(N__7575),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9562),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_15_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_15_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_15_12_5  (
            .in0(N__6955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7881),
            .lcout(\U712_CHIP_RAM.N_127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_15_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_15_12_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_15_12_6  (
            .in0(N__7112),
            .in1(N__7090),
            .in2(_gnd_net_),
            .in3(N__7061),
            .lcout(\U712_CHIP_RAM.N_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_15_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_15_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_15_12_7  (
            .in0(_gnd_net_),
            .in1(N__6855),
            .in2(_gnd_net_),
            .in3(N__7883),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER39_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_4_LC_15_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_4_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_4_LC_15_13_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_4_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__7015),
            .in2(_gnd_net_),
            .in3(N__6959),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER39_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_15_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_15_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_15_13_6 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_15_13_6  (
            .in0(N__6972),
            .in1(N__6886),
            .in2(N__6872),
            .in3(N__7887),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9567),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_15_14_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_15_14_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_15_14_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__6745),
            .in2(_gnd_net_),
            .in3(N__6696),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9571),
            .ce(),
            .sr(N__9331));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_15_14_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_15_14_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_15_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6669),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9571),
            .ce(),
            .sr(N__9331));
    defparam \U712_BUFFERS.DRDDIR_0_i_LC_15_15_3 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_0_i_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_0_i_LC_15_15_3 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \U712_BUFFERS.DRDDIR_0_i_LC_15_15_3  (
            .in0(N__9139),
            .in1(N__8200),
            .in2(N__7467),
            .in3(N__9180),
            .lcout(DRDDIR_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_16_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_16_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_16_5_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_16_5_3  (
            .in0(N__8819),
            .in1(N__8704),
            .in2(N__8886),
            .in3(N__8538),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9529),
            .ce(N__7393),
            .sr(N__9377));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7329),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9541),
            .ce(N__9058),
            .sr(N__9370));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_8_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_8_0  (
            .in0(N__7293),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9548),
            .ce(N__9045),
            .sr(N__9369));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_16_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_16_11_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_16_11_0  (
            .in0(N__7680),
            .in1(N__7255),
            .in2(N__7629),
            .in3(N__7240),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_16_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_16_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_16_11_1 .LUT_INIT=16'b0011111100110000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__7218),
            .in2(N__7162),
            .in3(N__8365),
            .lcout(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9563),
            .ce(),
            .sr(N__9358));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_16_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_16_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_16_11_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_16_11_3  (
            .in0(N__7159),
            .in1(N__9141),
            .in2(_gnd_net_),
            .in3(N__8127),
            .lcout(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9563),
            .ce(),
            .sr(N__9358));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_16_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_16_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_16_11_4 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_16_11_4  (
            .in0(N__7681),
            .in1(N__7147),
            .in2(_gnd_net_),
            .in3(N__8321),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9563),
            .ce(),
            .sr(N__9358));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI20AV_LC_16_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI20AV_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI20AV_LC_16_11_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI20AV_LC_16_11_5  (
            .in0(N__8377),
            .in1(N__8364),
            .in2(N__7524),
            .in3(N__7679),
            .lcout(\U712_CHIP_RAM.N_135 ),
            .ltout(\U712_CHIP_RAM.N_135_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMMGI5_LC_16_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMMGI5_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMMGI5_LC_16_11_6 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMMGI5_LC_16_11_6  (
            .in0(N__7571),
            .in1(N__8320),
            .in2(N__8302),
            .in3(N__8297),
            .lcout(\U712_CHIP_RAM.N_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_16_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_16_12_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_16_12_2  (
            .in0(N__7543),
            .in1(N__7611),
            .in2(N__7854),
            .in3(N__7678),
            .lcout(),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_16_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_16_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_16_12_3 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_16_12_3  (
            .in0(N__7900),
            .in1(N__8214),
            .in2(N__8275),
            .in3(N__8271),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9568),
            .ce(),
            .sr(N__9351));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_16_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_16_12_4 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_16_12_4  (
            .in0(N__8199),
            .in1(N__9140),
            .in2(N__8128),
            .in3(N__7929),
            .lcout(\U712_CHIP_RAM.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_16_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_16_12_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__7513),
            .in2(_gnd_net_),
            .in3(N__7880),
            .lcout(\U712_CHIP_RAM.N_63 ),
            .ltout(\U712_CHIP_RAM.N_63_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN14U1_LC_16_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN14U1_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN14U1_LC_16_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN14U1_LC_16_12_6  (
            .in0(N__7797),
            .in1(N__7677),
            .in2(N__7633),
            .in3(N__7610),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFMO84_3_LC_16_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFMO84_3_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFMO84_3_LC_16_12_7 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIFMO84_3_LC_16_12_7  (
            .in0(N__7569),
            .in1(N__7542),
            .in2(N__7528),
            .in3(N__7514),
            .lcout(\U712_CHIP_RAM.N_107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_DRDENn_LC_16_15_3 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_LC_16_15_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_LC_16_15_3  (
            .in0(N__9184),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9142),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_17_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_17_8_0 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_17_8_0  (
            .in0(N__9418),
            .in1(N__8548),
            .in2(_gnd_net_),
            .in3(N__9592),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_17_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_17_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_17_12_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_17_12_0  (
            .in0(N__9003),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9572),
            .ce(N__8934),
            .sr(N__9359));
    defparam \U712_CHIP_RAM.CRCSn_LC_18_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_18_4_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_18_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_18_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8887),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9533),
            .ce(),
            .sr(N__9380));
    defparam \U712_CHIP_RAM.RASn_LC_18_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_18_5_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_18_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_18_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8818),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9542),
            .ce(),
            .sr(N__9379));
    defparam \U712_CHIP_RAM.CASn_LC_18_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_18_5_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_18_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_18_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8701),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9542),
            .ce(),
            .sr(N__9379));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_18_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_18_8_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_18_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_18_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9591),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9560),
            .ce(),
            .sr(N__9375));
    defparam \U712_CHIP_RAM.WEn_LC_19_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_19_4_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_19_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_19_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8542),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9543),
            .ce(),
            .sr(N__9381));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_19_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_19_8_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_19_8_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_19_8_5  (
            .in0(_gnd_net_),
            .in1(N__8403),
            .in2(_gnd_net_),
            .in3(N__9601),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9564),
            .ce(),
            .sr(N__9378));
    defparam CONSTANT_ONE_LUT4_LC_20_4_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_20_4_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_20_4_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_20_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

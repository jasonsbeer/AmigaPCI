// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 8 2025 20:42:07

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    CMA,
    DRA,
    A,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    VBENn,
    CUMBEn,
    CLKRAM,
    C3,
    ASn,
    LDSn,
    CASUn,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40_OUT,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    DBRn,
    CLK40_IN,
    REGSPACEn,
    TSn,
    RASn,
    TACKn,
    C1);

    input [1:0] SIZ;
    output [10:0] CMA;
    input [9:0] DRA;
    input [20:0] A;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    input C3;
    output ASn;
    output LDSn;
    input CASUn;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40_OUT;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    input DBRn;
    input CLK40_IN;
    input REGSPACEn;
    input TSn;
    output RASn;
    output TACKn;
    input C1;

    wire N__10182;
    wire N__10181;
    wire N__10180;
    wire N__10173;
    wire N__10172;
    wire N__10171;
    wire N__10164;
    wire N__10163;
    wire N__10162;
    wire N__10155;
    wire N__10154;
    wire N__10153;
    wire N__10146;
    wire N__10145;
    wire N__10144;
    wire N__10137;
    wire N__10136;
    wire N__10135;
    wire N__10128;
    wire N__10127;
    wire N__10126;
    wire N__10119;
    wire N__10118;
    wire N__10117;
    wire N__10110;
    wire N__10109;
    wire N__10108;
    wire N__10101;
    wire N__10100;
    wire N__10099;
    wire N__10092;
    wire N__10091;
    wire N__10090;
    wire N__10083;
    wire N__10082;
    wire N__10081;
    wire N__10074;
    wire N__10073;
    wire N__10072;
    wire N__10065;
    wire N__10064;
    wire N__10063;
    wire N__10056;
    wire N__10055;
    wire N__10054;
    wire N__10047;
    wire N__10046;
    wire N__10045;
    wire N__10038;
    wire N__10037;
    wire N__10036;
    wire N__10029;
    wire N__10028;
    wire N__10027;
    wire N__10020;
    wire N__10019;
    wire N__10018;
    wire N__10011;
    wire N__10010;
    wire N__10009;
    wire N__10002;
    wire N__10001;
    wire N__10000;
    wire N__9993;
    wire N__9992;
    wire N__9991;
    wire N__9984;
    wire N__9983;
    wire N__9982;
    wire N__9975;
    wire N__9974;
    wire N__9973;
    wire N__9966;
    wire N__9965;
    wire N__9964;
    wire N__9957;
    wire N__9956;
    wire N__9955;
    wire N__9948;
    wire N__9947;
    wire N__9946;
    wire N__9939;
    wire N__9938;
    wire N__9937;
    wire N__9930;
    wire N__9929;
    wire N__9928;
    wire N__9921;
    wire N__9920;
    wire N__9919;
    wire N__9912;
    wire N__9911;
    wire N__9910;
    wire N__9903;
    wire N__9902;
    wire N__9901;
    wire N__9894;
    wire N__9893;
    wire N__9892;
    wire N__9885;
    wire N__9884;
    wire N__9883;
    wire N__9876;
    wire N__9875;
    wire N__9874;
    wire N__9867;
    wire N__9866;
    wire N__9865;
    wire N__9858;
    wire N__9857;
    wire N__9856;
    wire N__9849;
    wire N__9848;
    wire N__9847;
    wire N__9840;
    wire N__9839;
    wire N__9838;
    wire N__9831;
    wire N__9830;
    wire N__9829;
    wire N__9822;
    wire N__9821;
    wire N__9820;
    wire N__9813;
    wire N__9812;
    wire N__9811;
    wire N__9804;
    wire N__9803;
    wire N__9802;
    wire N__9795;
    wire N__9794;
    wire N__9793;
    wire N__9786;
    wire N__9785;
    wire N__9784;
    wire N__9777;
    wire N__9776;
    wire N__9775;
    wire N__9768;
    wire N__9767;
    wire N__9766;
    wire N__9759;
    wire N__9758;
    wire N__9757;
    wire N__9750;
    wire N__9749;
    wire N__9748;
    wire N__9741;
    wire N__9740;
    wire N__9739;
    wire N__9732;
    wire N__9731;
    wire N__9730;
    wire N__9723;
    wire N__9722;
    wire N__9721;
    wire N__9714;
    wire N__9713;
    wire N__9712;
    wire N__9705;
    wire N__9704;
    wire N__9703;
    wire N__9696;
    wire N__9695;
    wire N__9694;
    wire N__9687;
    wire N__9686;
    wire N__9685;
    wire N__9678;
    wire N__9677;
    wire N__9676;
    wire N__9669;
    wire N__9668;
    wire N__9667;
    wire N__9660;
    wire N__9659;
    wire N__9658;
    wire N__9651;
    wire N__9650;
    wire N__9649;
    wire N__9642;
    wire N__9641;
    wire N__9640;
    wire N__9633;
    wire N__9632;
    wire N__9631;
    wire N__9624;
    wire N__9623;
    wire N__9622;
    wire N__9615;
    wire N__9614;
    wire N__9613;
    wire N__9606;
    wire N__9605;
    wire N__9604;
    wire N__9597;
    wire N__9596;
    wire N__9595;
    wire N__9588;
    wire N__9587;
    wire N__9586;
    wire N__9579;
    wire N__9578;
    wire N__9577;
    wire N__9570;
    wire N__9569;
    wire N__9568;
    wire N__9561;
    wire N__9560;
    wire N__9559;
    wire N__9552;
    wire N__9551;
    wire N__9550;
    wire N__9543;
    wire N__9542;
    wire N__9541;
    wire N__9534;
    wire N__9533;
    wire N__9532;
    wire N__9525;
    wire N__9524;
    wire N__9523;
    wire N__9516;
    wire N__9515;
    wire N__9514;
    wire N__9507;
    wire N__9506;
    wire N__9505;
    wire N__9498;
    wire N__9497;
    wire N__9496;
    wire N__9489;
    wire N__9488;
    wire N__9487;
    wire N__9470;
    wire N__9469;
    wire N__9466;
    wire N__9463;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9427;
    wire N__9424;
    wire N__9421;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9391;
    wire N__9390;
    wire N__9389;
    wire N__9388;
    wire N__9387;
    wire N__9386;
    wire N__9385;
    wire N__9382;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9355;
    wire N__9354;
    wire N__9353;
    wire N__9352;
    wire N__9351;
    wire N__9348;
    wire N__9345;
    wire N__9342;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9294;
    wire N__9287;
    wire N__9286;
    wire N__9285;
    wire N__9284;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9274;
    wire N__9271;
    wire N__9268;
    wire N__9267;
    wire N__9266;
    wire N__9265;
    wire N__9264;
    wire N__9263;
    wire N__9262;
    wire N__9261;
    wire N__9260;
    wire N__9259;
    wire N__9258;
    wire N__9257;
    wire N__9256;
    wire N__9255;
    wire N__9254;
    wire N__9253;
    wire N__9250;
    wire N__9249;
    wire N__9248;
    wire N__9247;
    wire N__9246;
    wire N__9245;
    wire N__9244;
    wire N__9243;
    wire N__9240;
    wire N__9239;
    wire N__9238;
    wire N__9237;
    wire N__9236;
    wire N__9235;
    wire N__9234;
    wire N__9233;
    wire N__9232;
    wire N__9231;
    wire N__9230;
    wire N__9229;
    wire N__9228;
    wire N__9227;
    wire N__9224;
    wire N__9223;
    wire N__9222;
    wire N__9221;
    wire N__9218;
    wire N__9217;
    wire N__9216;
    wire N__9213;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8977;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8962;
    wire N__8959;
    wire N__8956;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8923;
    wire N__8922;
    wire N__8921;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8904;
    wire N__8899;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8875;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8836;
    wire N__8835;
    wire N__8834;
    wire N__8833;
    wire N__8832;
    wire N__8831;
    wire N__8830;
    wire N__8829;
    wire N__8828;
    wire N__8827;
    wire N__8826;
    wire N__8825;
    wire N__8824;
    wire N__8823;
    wire N__8822;
    wire N__8821;
    wire N__8820;
    wire N__8819;
    wire N__8818;
    wire N__8817;
    wire N__8816;
    wire N__8815;
    wire N__8814;
    wire N__8813;
    wire N__8810;
    wire N__8809;
    wire N__8808;
    wire N__8807;
    wire N__8806;
    wire N__8805;
    wire N__8804;
    wire N__8803;
    wire N__8802;
    wire N__8801;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8725;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8715;
    wire N__8712;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8704;
    wire N__8703;
    wire N__8700;
    wire N__8697;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8668;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8653;
    wire N__8650;
    wire N__8647;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8617;
    wire N__8614;
    wire N__8611;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8557;
    wire N__8554;
    wire N__8551;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8518;
    wire N__8517;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8503;
    wire N__8500;
    wire N__8497;
    wire N__8494;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8476;
    wire N__8475;
    wire N__8474;
    wire N__8473;
    wire N__8472;
    wire N__8471;
    wire N__8470;
    wire N__8467;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8443;
    wire N__8440;
    wire N__8439;
    wire N__8438;
    wire N__8437;
    wire N__8436;
    wire N__8435;
    wire N__8434;
    wire N__8433;
    wire N__8430;
    wire N__8429;
    wire N__8426;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8395;
    wire N__8394;
    wire N__8391;
    wire N__8388;
    wire N__8385;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8326;
    wire N__8325;
    wire N__8324;
    wire N__8319;
    wire N__8314;
    wire N__8313;
    wire N__8312;
    wire N__8309;
    wire N__8306;
    wire N__8301;
    wire N__8298;
    wire N__8295;
    wire N__8292;
    wire N__8289;
    wire N__8284;
    wire N__8279;
    wire N__8276;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8268;
    wire N__8265;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8237;
    wire N__8236;
    wire N__8231;
    wire N__8228;
    wire N__8227;
    wire N__8224;
    wire N__8221;
    wire N__8216;
    wire N__8213;
    wire N__8210;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8187;
    wire N__8182;
    wire N__8181;
    wire N__8178;
    wire N__8175;
    wire N__8172;
    wire N__8169;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8144;
    wire N__8141;
    wire N__8140;
    wire N__8137;
    wire N__8134;
    wire N__8133;
    wire N__8132;
    wire N__8131;
    wire N__8128;
    wire N__8127;
    wire N__8126;
    wire N__8123;
    wire N__8118;
    wire N__8115;
    wire N__8112;
    wire N__8107;
    wire N__8102;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8064;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8052;
    wire N__8051;
    wire N__8050;
    wire N__8047;
    wire N__8042;
    wire N__8037;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7966;
    wire N__7965;
    wire N__7960;
    wire N__7957;
    wire N__7956;
    wire N__7953;
    wire N__7948;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7921;
    wire N__7920;
    wire N__7919;
    wire N__7918;
    wire N__7915;
    wire N__7914;
    wire N__7913;
    wire N__7912;
    wire N__7911;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7903;
    wire N__7902;
    wire N__7899;
    wire N__7898;
    wire N__7897;
    wire N__7896;
    wire N__7891;
    wire N__7890;
    wire N__7889;
    wire N__7888;
    wire N__7887;
    wire N__7886;
    wire N__7885;
    wire N__7884;
    wire N__7881;
    wire N__7878;
    wire N__7875;
    wire N__7870;
    wire N__7865;
    wire N__7858;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7840;
    wire N__7837;
    wire N__7832;
    wire N__7825;
    wire N__7824;
    wire N__7819;
    wire N__7812;
    wire N__7811;
    wire N__7808;
    wire N__7801;
    wire N__7798;
    wire N__7795;
    wire N__7792;
    wire N__7789;
    wire N__7786;
    wire N__7783;
    wire N__7778;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7751;
    wire N__7748;
    wire N__7745;
    wire N__7742;
    wire N__7741;
    wire N__7738;
    wire N__7735;
    wire N__7730;
    wire N__7729;
    wire N__7726;
    wire N__7725;
    wire N__7722;
    wire N__7717;
    wire N__7714;
    wire N__7709;
    wire N__7708;
    wire N__7705;
    wire N__7702;
    wire N__7699;
    wire N__7696;
    wire N__7693;
    wire N__7690;
    wire N__7687;
    wire N__7684;
    wire N__7681;
    wire N__7678;
    wire N__7677;
    wire N__7672;
    wire N__7669;
    wire N__7664;
    wire N__7663;
    wire N__7662;
    wire N__7661;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7627;
    wire N__7624;
    wire N__7619;
    wire N__7616;
    wire N__7615;
    wire N__7612;
    wire N__7609;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7589;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7579;
    wire N__7578;
    wire N__7577;
    wire N__7568;
    wire N__7565;
    wire N__7564;
    wire N__7561;
    wire N__7560;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7548;
    wire N__7545;
    wire N__7538;
    wire N__7537;
    wire N__7536;
    wire N__7529;
    wire N__7526;
    wire N__7525;
    wire N__7524;
    wire N__7521;
    wire N__7514;
    wire N__7511;
    wire N__7510;
    wire N__7507;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7490;
    wire N__7489;
    wire N__7488;
    wire N__7485;
    wire N__7482;
    wire N__7479;
    wire N__7476;
    wire N__7473;
    wire N__7466;
    wire N__7465;
    wire N__7464;
    wire N__7461;
    wire N__7458;
    wire N__7455;
    wire N__7454;
    wire N__7453;
    wire N__7452;
    wire N__7451;
    wire N__7450;
    wire N__7449;
    wire N__7448;
    wire N__7447;
    wire N__7446;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7432;
    wire N__7431;
    wire N__7428;
    wire N__7425;
    wire N__7416;
    wire N__7413;
    wire N__7410;
    wire N__7407;
    wire N__7400;
    wire N__7397;
    wire N__7396;
    wire N__7395;
    wire N__7392;
    wire N__7391;
    wire N__7388;
    wire N__7387;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7374;
    wire N__7369;
    wire N__7368;
    wire N__7367;
    wire N__7366;
    wire N__7363;
    wire N__7360;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7342;
    wire N__7331;
    wire N__7324;
    wire N__7307;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7299;
    wire N__7298;
    wire N__7297;
    wire N__7296;
    wire N__7291;
    wire N__7286;
    wire N__7281;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7243;
    wire N__7240;
    wire N__7237;
    wire N__7234;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7220;
    wire N__7219;
    wire N__7218;
    wire N__7211;
    wire N__7208;
    wire N__7207;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7195;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7180;
    wire N__7175;
    wire N__7174;
    wire N__7173;
    wire N__7170;
    wire N__7167;
    wire N__7166;
    wire N__7163;
    wire N__7160;
    wire N__7155;
    wire N__7148;
    wire N__7147;
    wire N__7142;
    wire N__7141;
    wire N__7140;
    wire N__7139;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7124;
    wire N__7121;
    wire N__7112;
    wire N__7111;
    wire N__7110;
    wire N__7109;
    wire N__7108;
    wire N__7101;
    wire N__7096;
    wire N__7091;
    wire N__7090;
    wire N__7089;
    wire N__7088;
    wire N__7085;
    wire N__7078;
    wire N__7073;
    wire N__7072;
    wire N__7071;
    wire N__7070;
    wire N__7067;
    wire N__7064;
    wire N__7057;
    wire N__7052;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7042;
    wire N__7039;
    wire N__7034;
    wire N__7033;
    wire N__7032;
    wire N__7025;
    wire N__7022;
    wire N__7021;
    wire N__7018;
    wire N__7015;
    wire N__7012;
    wire N__7011;
    wire N__7010;
    wire N__7005;
    wire N__7000;
    wire N__6997;
    wire N__6992;
    wire N__6989;
    wire N__6988;
    wire N__6987;
    wire N__6980;
    wire N__6977;
    wire N__6974;
    wire N__6973;
    wire N__6970;
    wire N__6967;
    wire N__6962;
    wire N__6961;
    wire N__6958;
    wire N__6955;
    wire N__6950;
    wire N__6947;
    wire N__6944;
    wire N__6941;
    wire N__6938;
    wire N__6935;
    wire N__6932;
    wire N__6929;
    wire N__6926;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6911;
    wire N__6908;
    wire N__6905;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6883;
    wire N__6882;
    wire N__6881;
    wire N__6878;
    wire N__6877;
    wire N__6876;
    wire N__6873;
    wire N__6872;
    wire N__6871;
    wire N__6868;
    wire N__6863;
    wire N__6860;
    wire N__6859;
    wire N__6856;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6837;
    wire N__6834;
    wire N__6821;
    wire N__6818;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6800;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6787;
    wire N__6784;
    wire N__6781;
    wire N__6778;
    wire N__6775;
    wire N__6770;
    wire N__6767;
    wire N__6766;
    wire N__6765;
    wire N__6762;
    wire N__6759;
    wire N__6756;
    wire N__6753;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6727;
    wire N__6724;
    wire N__6721;
    wire N__6720;
    wire N__6719;
    wire N__6718;
    wire N__6715;
    wire N__6714;
    wire N__6711;
    wire N__6708;
    wire N__6707;
    wire N__6702;
    wire N__6701;
    wire N__6698;
    wire N__6697;
    wire N__6696;
    wire N__6695;
    wire N__6694;
    wire N__6693;
    wire N__6692;
    wire N__6691;
    wire N__6688;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6676;
    wire N__6673;
    wire N__6670;
    wire N__6667;
    wire N__6662;
    wire N__6657;
    wire N__6652;
    wire N__6629;
    wire N__6628;
    wire N__6627;
    wire N__6624;
    wire N__6623;
    wire N__6620;
    wire N__6617;
    wire N__6616;
    wire N__6615;
    wire N__6614;
    wire N__6613;
    wire N__6612;
    wire N__6611;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6599;
    wire N__6596;
    wire N__6593;
    wire N__6588;
    wire N__6585;
    wire N__6580;
    wire N__6563;
    wire N__6560;
    wire N__6557;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6542;
    wire N__6541;
    wire N__6540;
    wire N__6537;
    wire N__6534;
    wire N__6529;
    wire N__6528;
    wire N__6523;
    wire N__6520;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6500;
    wire N__6497;
    wire N__6494;
    wire N__6493;
    wire N__6490;
    wire N__6487;
    wire N__6482;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6452;
    wire N__6449;
    wire N__6446;
    wire N__6445;
    wire N__6444;
    wire N__6441;
    wire N__6438;
    wire N__6435;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6404;
    wire N__6403;
    wire N__6402;
    wire N__6401;
    wire N__6398;
    wire N__6397;
    wire N__6396;
    wire N__6391;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6381;
    wire N__6380;
    wire N__6377;
    wire N__6376;
    wire N__6375;
    wire N__6372;
    wire N__6369;
    wire N__6366;
    wire N__6363;
    wire N__6358;
    wire N__6353;
    wire N__6350;
    wire N__6347;
    wire N__6332;
    wire N__6329;
    wire N__6326;
    wire N__6323;
    wire N__6322;
    wire N__6321;
    wire N__6320;
    wire N__6317;
    wire N__6316;
    wire N__6313;
    wire N__6312;
    wire N__6309;
    wire N__6306;
    wire N__6305;
    wire N__6302;
    wire N__6299;
    wire N__6298;
    wire N__6297;
    wire N__6296;
    wire N__6295;
    wire N__6290;
    wire N__6285;
    wire N__6282;
    wire N__6277;
    wire N__6274;
    wire N__6273;
    wire N__6270;
    wire N__6269;
    wire N__6268;
    wire N__6267;
    wire N__6266;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6234;
    wire N__6227;
    wire N__6206;
    wire N__6203;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6191;
    wire N__6188;
    wire N__6187;
    wire N__6186;
    wire N__6185;
    wire N__6182;
    wire N__6181;
    wire N__6178;
    wire N__6177;
    wire N__6176;
    wire N__6175;
    wire N__6172;
    wire N__6171;
    wire N__6168;
    wire N__6165;
    wire N__6162;
    wire N__6161;
    wire N__6158;
    wire N__6157;
    wire N__6152;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6137;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6122;
    wire N__6119;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6088;
    wire N__6085;
    wire N__6084;
    wire N__6081;
    wire N__6080;
    wire N__6079;
    wire N__6078;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6065;
    wire N__6062;
    wire N__6061;
    wire N__6060;
    wire N__6057;
    wire N__6056;
    wire N__6055;
    wire N__6054;
    wire N__6053;
    wire N__6050;
    wire N__6045;
    wire N__6044;
    wire N__6043;
    wire N__6042;
    wire N__6041;
    wire N__6038;
    wire N__6033;
    wire N__6030;
    wire N__6027;
    wire N__6024;
    wire N__6021;
    wire N__6016;
    wire N__6013;
    wire N__6008;
    wire N__6003;
    wire N__5998;
    wire N__5993;
    wire N__5972;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5964;
    wire N__5963;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5932;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5915;
    wire N__5912;
    wire N__5911;
    wire N__5906;
    wire N__5903;
    wire N__5900;
    wire N__5897;
    wire N__5894;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5825;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5759;
    wire N__5756;
    wire N__5753;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5729;
    wire N__5726;
    wire N__5723;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5705;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5635;
    wire N__5634;
    wire N__5631;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5619;
    wire N__5616;
    wire N__5613;
    wire N__5610;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5526;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5512;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5489;
    wire N__5488;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5459;
    wire N__5458;
    wire N__5453;
    wire N__5452;
    wire N__5451;
    wire N__5448;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5434;
    wire N__5431;
    wire N__5428;
    wire N__5425;
    wire N__5420;
    wire N__5417;
    wire N__5416;
    wire N__5415;
    wire N__5414;
    wire N__5405;
    wire N__5402;
    wire N__5401;
    wire N__5396;
    wire N__5393;
    wire N__5390;
    wire N__5389;
    wire N__5388;
    wire N__5385;
    wire N__5380;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5336;
    wire N__5335;
    wire N__5334;
    wire N__5331;
    wire N__5326;
    wire N__5325;
    wire N__5320;
    wire N__5317;
    wire N__5316;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5304;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5242;
    wire N__5241;
    wire N__5240;
    wire N__5239;
    wire N__5236;
    wire N__5233;
    wire N__5230;
    wire N__5227;
    wire N__5224;
    wire N__5217;
    wire N__5214;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5192;
    wire N__5191;
    wire N__5188;
    wire N__5187;
    wire N__5184;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5156;
    wire N__5155;
    wire N__5154;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5143;
    wire N__5142;
    wire N__5141;
    wire N__5140;
    wire N__5139;
    wire N__5138;
    wire N__5137;
    wire N__5134;
    wire N__5133;
    wire N__5128;
    wire N__5123;
    wire N__5122;
    wire N__5119;
    wire N__5118;
    wire N__5117;
    wire N__5114;
    wire N__5113;
    wire N__5110;
    wire N__5105;
    wire N__5102;
    wire N__5097;
    wire N__5092;
    wire N__5089;
    wire N__5086;
    wire N__5081;
    wire N__5076;
    wire N__5057;
    wire N__5056;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5046;
    wire N__5045;
    wire N__5044;
    wire N__5043;
    wire N__5038;
    wire N__5031;
    wire N__5028;
    wire N__5021;
    wire N__5020;
    wire N__5017;
    wire N__5014;
    wire N__5011;
    wire N__5006;
    wire N__5005;
    wire N__5002;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4987;
    wire N__4982;
    wire N__4981;
    wire N__4980;
    wire N__4979;
    wire N__4976;
    wire N__4975;
    wire N__4972;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4960;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4948;
    wire N__4943;
    wire N__4936;
    wire N__4931;
    wire N__4930;
    wire N__4929;
    wire N__4926;
    wire N__4925;
    wire N__4924;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4902;
    wire N__4889;
    wire N__4888;
    wire N__4887;
    wire N__4886;
    wire N__4885;
    wire N__4884;
    wire N__4883;
    wire N__4882;
    wire N__4879;
    wire N__4872;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4799;
    wire N__4796;
    wire N__4795;
    wire N__4794;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4778;
    wire N__4775;
    wire N__4774;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4759;
    wire N__4758;
    wire N__4755;
    wire N__4750;
    wire N__4745;
    wire N__4744;
    wire N__4741;
    wire N__4738;
    wire N__4733;
    wire N__4732;
    wire N__4729;
    wire N__4726;
    wire N__4721;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4711;
    wire N__4706;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4694;
    wire N__4691;
    wire N__4690;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4673;
    wire N__4672;
    wire N__4669;
    wire N__4666;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4483;
    wire N__4482;
    wire N__4477;
    wire N__4474;
    wire N__4469;
    wire N__4466;
    wire N__4465;
    wire N__4464;
    wire N__4463;
    wire N__4458;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4445;
    wire N__4440;
    wire N__4433;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4397;
    wire N__4396;
    wire N__4395;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4363;
    wire N__4360;
    wire N__4357;
    wire N__4354;
    wire N__4351;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4309;
    wire N__4308;
    wire N__4305;
    wire N__4300;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4279;
    wire N__4276;
    wire N__4273;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4222;
    wire N__4219;
    wire N__4216;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4133;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4045;
    wire N__4042;
    wire N__4039;
    wire N__4038;
    wire N__4035;
    wire N__4032;
    wire N__4029;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3934;
    wire N__3929;
    wire N__3926;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3916;
    wire N__3913;
    wire N__3910;
    wire N__3905;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3887;
    wire N__3884;
    wire N__3881;
    wire N__3878;
    wire N__3875;
    wire N__3874;
    wire N__3873;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3859;
    wire N__3856;
    wire N__3853;
    wire N__3850;
    wire N__3847;
    wire N__3842;
    wire N__3839;
    wire N__3838;
    wire N__3835;
    wire N__3832;
    wire N__3827;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3815;
    wire N__3812;
    wire N__3811;
    wire N__3808;
    wire N__3805;
    wire N__3800;
    wire N__3797;
    wire N__3796;
    wire N__3793;
    wire N__3790;
    wire N__3785;
    wire N__3782;
    wire N__3779;
    wire N__3778;
    wire N__3775;
    wire N__3772;
    wire N__3769;
    wire N__3764;
    wire N__3761;
    wire N__3760;
    wire N__3757;
    wire N__3754;
    wire N__3749;
    wire N__3746;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3734;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3703;
    wire N__3702;
    wire N__3697;
    wire N__3694;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3680;
    wire N__3677;
    wire N__3674;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3662;
    wire N__3661;
    wire N__3660;
    wire N__3659;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3629;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3617;
    wire N__3614;
    wire N__3611;
    wire N__3608;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK40_PLL_i_i;
    wire N_981_i;
    wire CLK80_PLL_i_i;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire TACK_OUTn;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire CLK40_PLL_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_7_7_0_;
    wire \U712_CHIP_RAM.REFRESH5lto1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH5lto2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire DBDIR_c;
    wire TACK_EN_i_ess;
    wire VBENn_c;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1 ;
    wire \U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_2 ;
    wire RAMSPACEn_c;
    wire \U712_CHIP_RAM.un5_DMA_CYCLE_START_0 ;
    wire REG_CYCLEm;
    wire DRDENn_c;
    wire A_c_16;
    wire A_c_18;
    wire A_c_11;
    wire A_c_4;
    wire A_c_9;
    wire A_c_2;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_1_cascade_ ;
    wire A_c_12;
    wire A_c_5;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_1_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_i_i_a3_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_cascade_ ;
    wire \U712_CHIP_RAM.CLK_EN_e_1_cascade_ ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.N_176_cascade_ ;
    wire \U712_CHIP_RAM.N_166_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.N_313 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_9_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0_a3_0 ;
    wire \U712_CHIP_RAM.N_232_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0_a3_1 ;
    wire \U712_CHIP_RAM.N_232 ;
    wire \U712_CHIP_RAM.BANK0_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_167_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_9_0_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire SIZ_c_1;
    wire CONSTANT_ONE_NET;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire A_c_13;
    wire A_c_6;
    wire A_c_15;
    wire A_c_8;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNIIGLS1Z0Z_0 ;
    wire \U712_CHIP_RAM.N_176 ;
    wire \U712_CHIP_RAM.N_230_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_a3_1_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_285_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ;
    wire \U712_CHIP_RAM.N_314 ;
    wire bfn_10_9_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.N_167 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1 ;
    wire \U712_CHIP_RAM.N_53 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.N_196_cascade_ ;
    wire \U712_CHIP_RAM.N_315 ;
    wire \U712_CHIP_RAM.N_197_i_cascade_ ;
    wire \U712_CHIP_RAM.N_233 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8RZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.N_219_cascade_ ;
    wire \U712_CHIP_RAM.N_166 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_7_i_2_cascade_ ;
    wire \U712_CHIP_RAM.N_258 ;
    wire \U712_CHIP_RAM.N_49_cascade_ ;
    wire \U712_CHIP_RAM.N_206 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_1 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire DBENn_c;
    wire \U712_BYTE_ENABLE.N_268 ;
    wire N_185_i;
    wire \U712_BYTE_ENABLE.N_270_cascade_ ;
    wire N_186_i;
    wire \U712_BYTE_ENABLE.N_272 ;
    wire CASLn_c;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0 ;
    wire N_187_i;
    wire A_c_1;
    wire \U712_BYTE_ENABLE.N_265 ;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0 ;
    wire \U712_BYTE_ENABLE.N_266_cascade_ ;
    wire CASUn_c;
    wire N_184_i;
    wire DMA_CYCLEm;
    wire DRDDIR_i_m2;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_ ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire A_c_14;
    wire A_c_3;
    wire A_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire CMA_c_5;
    wire A_c_7;
    wire \U712_CHIP_RAM.N_324_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire RnW_c;
    wire AWEn_c;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.N_248 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2Z0Z_1 ;
    wire \U712_REG_SM.N_171_cascade_ ;
    wire \U712_REG_SM.DS_EN_0_sqmuxa_0_a2_0_a3_1_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_6 ;
    wire \U712_REG_SM.N_199_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.N_208_i_0_en_cascade_ ;
    wire \U712_CYCLE_TERM.N_208_i_0_en_0 ;
    wire \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a3_0_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_165 ;
    wire \U712_CHIP_RAM.N_249 ;
    wire CPU_TACKm;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_REG_SM.N_199 ;
    wire \U712_REG_SM.N_171 ;
    wire \U712_REG_SM.N_174_cascade_ ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_REG_SM.N_210 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_5 ;
    wire \U712_REG_SM.N_174 ;
    wire REG_TACK;
    wire DBR_SYNCZ0Z_0;
    wire CASn_c;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_ ;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire C3_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_2 ;
    wire C1_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_2 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire ASn_c;
    wire \U712_REG_SM.STATE_COUNT_RNITQLC2Z0Z_1 ;
    wire REGSPACEn_c;
    wire \U712_REG_SM.REG_CYCLE_GOZ0 ;
    wire TSn_c;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.DS_EN_0_sqmuxa ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_REG_SM.N_205 ;
    wire \U712_REG_SM.N_202 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire C1_c_g;
    wire RESETn_c;
    wire RESETn_c_i;
    wire N_118;
    wire A_c_0;
    wire SIZ_c_0;
    wire DS_ENm;
    wire N_113;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire WEn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire A_c_17;
    wire CPU_CYCLEm;
    wire CMA_c_8;
    wire CLK80_PLL;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire DBRn_c;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ;
    wire RAS0n_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire _gnd_net_;
    wire C3_c_g;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ;
    wire RESETn_c_i_g;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__3620),
            .RESETB(N__4373),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__10182),
            .DIN(N__10181),
            .DOUT(N__10180),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__10182),
            .PADOUT(N__10181),
            .PADIN(N__10180),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5645),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__10173),
            .DIN(N__10172),
            .DOUT(N__10171),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__10173),
            .PADOUT(N__10172),
            .PADIN(N__10171),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__10164),
            .DIN(N__10163),
            .DOUT(N__10162),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__10164),
            .PADOUT(N__10163),
            .PADIN(N__10162),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6950),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__10155),
            .DIN(N__10154),
            .DOUT(N__10153),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__10155),
            .PADOUT(N__10154),
            .PADIN(N__10153),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5297),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__10146),
            .DIN(N__10145),
            .DOUT(N__10144),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__10146),
            .PADOUT(N__10145),
            .PADIN(N__10144),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__10137),
            .DIN(N__10136),
            .DOUT(N__10135),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__10137),
            .PADOUT(N__10136),
            .PADIN(N__10135),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__10128),
            .DIN(N__10127),
            .DOUT(N__10126),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__10128),
            .PADOUT(N__10127),
            .PADIN(N__10126),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__10119),
            .DIN(N__10118),
            .DOUT(N__10117),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__10119),
            .PADOUT(N__10118),
            .PADIN(N__10117),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__10110),
            .DIN(N__10109),
            .DOUT(N__10108),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__10110),
            .PADOUT(N__10109),
            .PADIN(N__10108),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__10101),
            .DIN(N__10100),
            .DOUT(N__10099),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__10101),
            .PADOUT(N__10100),
            .PADIN(N__10099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5741),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__10092),
            .DIN(N__10091),
            .DOUT(N__10090),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__10092),
            .PADOUT(N__10091),
            .PADIN(N__10090),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__10083),
            .DIN(N__10082),
            .DOUT(N__10081),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__10083),
            .PADOUT(N__10082),
            .PADIN(N__10081),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__10074),
            .DIN(N__10073),
            .DOUT(N__10072),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__10074),
            .PADOUT(N__10073),
            .PADIN(N__10072),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__10065),
            .DIN(N__10064),
            .DOUT(N__10063),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__10065),
            .PADOUT(N__10064),
            .PADIN(N__10063),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3893),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__10056),
            .DIN(N__10055),
            .DOUT(N__10054),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__10056),
            .PADOUT(N__10055),
            .PADIN(N__10054),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__10047),
            .DIN(N__10046),
            .DOUT(N__10045),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__10047),
            .PADOUT(N__10046),
            .PADIN(N__10045),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__10038),
            .DIN(N__10037),
            .DOUT(N__10036),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__10038),
            .PADOUT(N__10037),
            .PADIN(N__10036),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5270),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__10029),
            .DIN(N__10028),
            .DOUT(N__10027),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__10029),
            .PADOUT(N__10028),
            .PADIN(N__10027),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__10020),
            .DIN(N__10019),
            .DOUT(N__10018),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__10020),
            .PADOUT(N__10019),
            .PADIN(N__10018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8162),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__10011),
            .DIN(N__10010),
            .DOUT(N__10009),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__10011),
            .PADOUT(N__10010),
            .PADIN(N__10009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__10002),
            .DIN(N__10001),
            .DOUT(N__10000),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__10002),
            .PADOUT(N__10001),
            .PADIN(N__10000),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__9993),
            .DIN(N__9992),
            .DOUT(N__9991),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__9993),
            .PADOUT(N__9992),
            .PADIN(N__9991),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__9984),
            .DIN(N__9983),
            .DOUT(N__9982),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__9984),
            .PADOUT(N__9983),
            .PADIN(N__9982),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__9975),
            .DIN(N__9974),
            .DOUT(N__9973),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__9975),
            .PADOUT(N__9974),
            .PADIN(N__9973),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__9966),
            .DIN(N__9965),
            .DOUT(N__9964),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__9966),
            .PADOUT(N__9965),
            .PADIN(N__9964),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4238),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__9957),
            .DIN(N__9956),
            .DOUT(N__9955),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__9957),
            .PADOUT(N__9956),
            .PADIN(N__9955),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__9948),
            .DIN(N__9947),
            .DOUT(N__9946),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__9948),
            .PADOUT(N__9947),
            .PADIN(N__9946),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__9939),
            .DIN(N__9938),
            .DOUT(N__9937),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__9939),
            .PADOUT(N__9938),
            .PADIN(N__9937),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__9930),
            .DIN(N__9929),
            .DOUT(N__9928),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__9930),
            .PADOUT(N__9929),
            .PADIN(N__9928),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__9921),
            .DIN(N__9920),
            .DOUT(N__9919),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__9921),
            .PADOUT(N__9920),
            .PADIN(N__9919),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__9912),
            .DIN(N__9911),
            .DOUT(N__9910),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__9912),
            .PADOUT(N__9911),
            .PADIN(N__9910),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5714),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__9903),
            .DIN(N__9902),
            .DOUT(N__9901),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__9903),
            .PADOUT(N__9902),
            .PADIN(N__9901),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__9894),
            .DIN(N__9893),
            .DOUT(N__9892),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__9894),
            .PADOUT(N__9893),
            .PADIN(N__9892),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__9885),
            .DIN(N__9884),
            .DOUT(N__9883),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__9885),
            .PADOUT(N__9884),
            .PADIN(N__9883),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__9876),
            .DIN(N__9875),
            .DOUT(N__9874),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__9876),
            .PADOUT(N__9875),
            .PADIN(N__9874),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__9867),
            .DIN(N__9866),
            .DOUT(N__9865),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__9867),
            .PADOUT(N__9866),
            .PADIN(N__9865),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8342),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__9858),
            .DIN(N__9857),
            .DOUT(N__9856),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__9858),
            .PADOUT(N__9857),
            .PADIN(N__9856),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__9849),
            .DIN(N__9848),
            .DOUT(N__9847),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__9849),
            .PADOUT(N__9848),
            .PADIN(N__9847),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8030),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__9840),
            .DIN(N__9839),
            .DOUT(N__9838),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__9840),
            .PADOUT(N__9839),
            .PADIN(N__9838),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__9831),
            .DIN(N__9830),
            .DOUT(N__9829),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__9831),
            .PADOUT(N__9830),
            .PADIN(N__9829),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__9822),
            .DIN(N__9821),
            .DOUT(N__9820),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__9822),
            .PADOUT(N__9821),
            .PADIN(N__9820),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3728),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__9813),
            .DIN(N__9812),
            .DOUT(N__9811),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__9813),
            .PADOUT(N__9812),
            .PADIN(N__9811),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7709),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__9804),
            .DIN(N__9803),
            .DOUT(N__9802),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__9804),
            .PADOUT(N__9803),
            .PADIN(N__9802),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6815),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__9795),
            .DIN(N__9794),
            .DOUT(N__9793),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__9795),
            .PADOUT(N__9794),
            .PADIN(N__9793),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__9786),
            .DIN(N__9785),
            .DOUT(N__9784),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__9786),
            .PADOUT(N__9785),
            .PADIN(N__9784),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_0_iopad (
            .OE(N__9777),
            .DIN(N__9776),
            .DOUT(N__9775),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__9777),
            .PADOUT(N__9776),
            .PADIN(N__9775),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__9768),
            .DIN(N__9767),
            .DOUT(N__9766),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__9768),
            .PADOUT(N__9767),
            .PADIN(N__9766),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6935),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__9759),
            .DIN(N__9758),
            .DOUT(N__9757),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__9759),
            .PADOUT(N__9758),
            .PADIN(N__9757),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__9750),
            .DIN(N__9749),
            .DOUT(N__9748),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__9750),
            .PADOUT(N__9749),
            .PADIN(N__9748),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5681),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__9741),
            .DIN(N__9740),
            .DOUT(N__9739),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__9741),
            .PADOUT(N__9740),
            .PADIN(N__9739),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4022),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__9732),
            .DIN(N__9731),
            .DOUT(N__9730),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__9732),
            .PADOUT(N__9731),
            .PADIN(N__9730),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5480),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__9723),
            .DIN(N__9722),
            .DOUT(N__9721),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__9723),
            .PADOUT(N__9722),
            .PADIN(N__9721),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7988),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__9714),
            .DIN(N__9713),
            .DOUT(N__9712),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__9714),
            .PADOUT(N__9713),
            .PADIN(N__9712),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7708),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__9705),
            .DIN(N__9704),
            .DOUT(N__9703),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__9705),
            .PADOUT(N__9704),
            .PADIN(N__9703),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__9696),
            .DIN(N__9695),
            .DOUT(N__9694),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__9696),
            .PADOUT(N__9695),
            .PADIN(N__9694),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__9687),
            .DIN(N__9686),
            .DOUT(N__9685),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__9687),
            .PADOUT(N__9686),
            .PADIN(N__9685),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5570),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__9678),
            .DIN(N__9677),
            .DOUT(N__9676),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__9678),
            .PADOUT(N__9677),
            .PADIN(N__9676),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8093),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__9669),
            .DIN(N__9668),
            .DOUT(N__9667),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__9669),
            .PADOUT(N__9668),
            .PADIN(N__9667),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3923),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_OUT_obuf_iopad (
            .OE(N__9660),
            .DIN(N__9659),
            .DOUT(N__9658),
            .PACKAGEPIN(CLK40_OUT));
    defparam CLK40_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40_OUT_obuf_preio (
            .PADOEN(N__9660),
            .PADOUT(N__9659),
            .PADIN(N__9658),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3647),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__9651),
            .DIN(N__9650),
            .DOUT(N__9649),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__9651),
            .PADOUT(N__9650),
            .PADIN(N__9649),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5597),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__9642),
            .DIN(N__9641),
            .DOUT(N__9640),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__9642),
            .PADOUT(N__9641),
            .PADIN(N__9640),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__9633),
            .DIN(N__9632),
            .DOUT(N__9631),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__9633),
            .PADOUT(N__9632),
            .PADIN(N__9631),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__9624),
            .DIN(N__9623),
            .DOUT(N__9622),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__9624),
            .PADOUT(N__9623),
            .PADIN(N__9622),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__9615),
            .DIN(N__9614),
            .DOUT(N__9613),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__9615),
            .PADOUT(N__9614),
            .PADIN(N__9613),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__9606),
            .DIN(N__9605),
            .DOUT(N__9604),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__9606),
            .PADOUT(N__9605),
            .PADIN(N__9604),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5831),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__9597),
            .DIN(N__9596),
            .DOUT(N__9595),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__9597),
            .PADOUT(N__9596),
            .PADIN(N__9595),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__9588),
            .DIN(N__9587),
            .DOUT(N__9586),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__9588),
            .PADOUT(N__9587),
            .PADIN(N__9586),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5366),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__9579),
            .DIN(N__9578),
            .DOUT(N__9577),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__9579),
            .PADOUT(N__9578),
            .PADIN(N__9577),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3638),
            .DIN0(),
            .DOUT0(N__3689),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__9570),
            .DIN(N__9569),
            .DOUT(N__9568),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__9570),
            .PADOUT(N__9569),
            .PADIN(N__9568),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6902),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__9561),
            .DIN(N__9560),
            .DOUT(N__9559),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__9561),
            .PADOUT(N__9560),
            .PADIN(N__9559),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__9552),
            .DIN(N__9551),
            .DOUT(N__9550),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__9552),
            .PADOUT(N__9551),
            .PADIN(N__9550),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__9543),
            .DIN(N__9542),
            .DOUT(N__9541),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__9543),
            .PADOUT(N__9542),
            .PADIN(N__9541),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7763),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__9534),
            .DIN(N__9533),
            .DOUT(N__9532),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__9534),
            .PADOUT(N__9533),
            .PADIN(N__9532),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__9525),
            .DIN(N__9524),
            .DOUT(N__9523),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__9525),
            .PADOUT(N__9524),
            .PADIN(N__9523),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__9516),
            .DIN(N__9515),
            .DOUT(N__9514),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__9516),
            .PADOUT(N__9515),
            .PADIN(N__9514),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__9507),
            .DIN(N__9506),
            .DOUT(N__9505),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__9507),
            .PADOUT(N__9506),
            .PADIN(N__9505),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__9498),
            .DIN(N__9497),
            .DOUT(N__9496),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__9498),
            .PADOUT(N__9497),
            .PADIN(N__9496),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5798),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__9489),
            .DIN(N__9488),
            .DOUT(N__9487),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__9489),
            .PADOUT(N__9488),
            .PADIN(N__9487),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8216),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2267 (
            .O(N__9470),
            .I(N__9466));
    InMux I__2266 (
            .O(N__9469),
            .I(N__9463));
    LocalMux I__2265 (
            .O(N__9466),
            .I(N__9458));
    LocalMux I__2264 (
            .O(N__9463),
            .I(N__9458));
    Span4Mux_v I__2263 (
            .O(N__9458),
            .I(N__9455));
    Span4Mux_v I__2262 (
            .O(N__9455),
            .I(N__9452));
    Sp12to4 I__2261 (
            .O(N__9452),
            .I(N__9449));
    Span12Mux_h I__2260 (
            .O(N__9449),
            .I(N__9446));
    Odrv12 I__2259 (
            .O(N__9446),
            .I(DRA_c_3));
    InMux I__2258 (
            .O(N__9443),
            .I(N__9440));
    LocalMux I__2257 (
            .O(N__9440),
            .I(N__9437));
    Span4Mux_h I__2256 (
            .O(N__9437),
            .I(N__9434));
    Odrv4 I__2255 (
            .O(N__9434),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__2254 (
            .O(N__9431),
            .I(N__9428));
    LocalMux I__2253 (
            .O(N__9428),
            .I(N__9424));
    InMux I__2252 (
            .O(N__9427),
            .I(N__9421));
    Span12Mux_v I__2251 (
            .O(N__9424),
            .I(N__9416));
    LocalMux I__2250 (
            .O(N__9421),
            .I(N__9416));
    Span12Mux_h I__2249 (
            .O(N__9416),
            .I(N__9413));
    Odrv12 I__2248 (
            .O(N__9413),
            .I(DRA_c_8));
    CascadeMux I__2247 (
            .O(N__9410),
            .I(N__9407));
    InMux I__2246 (
            .O(N__9407),
            .I(N__9404));
    LocalMux I__2245 (
            .O(N__9404),
            .I(N__9401));
    Span4Mux_h I__2244 (
            .O(N__9401),
            .I(N__9398));
    Odrv4 I__2243 (
            .O(N__9398),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2242 (
            .O(N__9395),
            .I(N__9392));
    LocalMux I__2241 (
            .O(N__9392),
            .I(N__9382));
    ClkMux I__2240 (
            .O(N__9391),
            .I(N__9365));
    ClkMux I__2239 (
            .O(N__9390),
            .I(N__9365));
    ClkMux I__2238 (
            .O(N__9389),
            .I(N__9365));
    ClkMux I__2237 (
            .O(N__9388),
            .I(N__9365));
    ClkMux I__2236 (
            .O(N__9387),
            .I(N__9365));
    ClkMux I__2235 (
            .O(N__9386),
            .I(N__9365));
    ClkMux I__2234 (
            .O(N__9385),
            .I(N__9365));
    Glb2LocalMux I__2233 (
            .O(N__9382),
            .I(N__9365));
    GlobalMux I__2232 (
            .O(N__9365),
            .I(N__9362));
    gio2CtrlBuf I__2231 (
            .O(N__9362),
            .I(C3_c_g));
    CEMux I__2230 (
            .O(N__9359),
            .I(N__9356));
    LocalMux I__2229 (
            .O(N__9356),
            .I(N__9348));
    CEMux I__2228 (
            .O(N__9355),
            .I(N__9345));
    CEMux I__2227 (
            .O(N__9354),
            .I(N__9342));
    CEMux I__2226 (
            .O(N__9353),
            .I(N__9338));
    CEMux I__2225 (
            .O(N__9352),
            .I(N__9335));
    CEMux I__2224 (
            .O(N__9351),
            .I(N__9332));
    Span4Mux_v I__2223 (
            .O(N__9348),
            .I(N__9329));
    LocalMux I__2222 (
            .O(N__9345),
            .I(N__9324));
    LocalMux I__2221 (
            .O(N__9342),
            .I(N__9324));
    CEMux I__2220 (
            .O(N__9341),
            .I(N__9321));
    LocalMux I__2219 (
            .O(N__9338),
            .I(N__9318));
    LocalMux I__2218 (
            .O(N__9335),
            .I(N__9315));
    LocalMux I__2217 (
            .O(N__9332),
            .I(N__9312));
    Span4Mux_h I__2216 (
            .O(N__9329),
            .I(N__9305));
    Span4Mux_v I__2215 (
            .O(N__9324),
            .I(N__9305));
    LocalMux I__2214 (
            .O(N__9321),
            .I(N__9305));
    Span4Mux_v I__2213 (
            .O(N__9318),
            .I(N__9302));
    Span4Mux_h I__2212 (
            .O(N__9315),
            .I(N__9299));
    Span4Mux_v I__2211 (
            .O(N__9312),
            .I(N__9294));
    Span4Mux_h I__2210 (
            .O(N__9305),
            .I(N__9294));
    Odrv4 I__2209 (
            .O(N__9302),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ));
    Odrv4 I__2208 (
            .O(N__9299),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ));
    Odrv4 I__2207 (
            .O(N__9294),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ));
    InMux I__2206 (
            .O(N__9287),
            .I(N__9280));
    InMux I__2205 (
            .O(N__9286),
            .I(N__9277));
    InMux I__2204 (
            .O(N__9285),
            .I(N__9274));
    InMux I__2203 (
            .O(N__9284),
            .I(N__9271));
    InMux I__2202 (
            .O(N__9283),
            .I(N__9268));
    LocalMux I__2201 (
            .O(N__9280),
            .I(N__9250));
    LocalMux I__2200 (
            .O(N__9277),
            .I(N__9240));
    LocalMux I__2199 (
            .O(N__9274),
            .I(N__9224));
    LocalMux I__2198 (
            .O(N__9271),
            .I(N__9218));
    LocalMux I__2197 (
            .O(N__9268),
            .I(N__9213));
    SRMux I__2196 (
            .O(N__9267),
            .I(N__9122));
    SRMux I__2195 (
            .O(N__9266),
            .I(N__9122));
    SRMux I__2194 (
            .O(N__9265),
            .I(N__9122));
    SRMux I__2193 (
            .O(N__9264),
            .I(N__9122));
    SRMux I__2192 (
            .O(N__9263),
            .I(N__9122));
    SRMux I__2191 (
            .O(N__9262),
            .I(N__9122));
    SRMux I__2190 (
            .O(N__9261),
            .I(N__9122));
    SRMux I__2189 (
            .O(N__9260),
            .I(N__9122));
    SRMux I__2188 (
            .O(N__9259),
            .I(N__9122));
    SRMux I__2187 (
            .O(N__9258),
            .I(N__9122));
    SRMux I__2186 (
            .O(N__9257),
            .I(N__9122));
    SRMux I__2185 (
            .O(N__9256),
            .I(N__9122));
    SRMux I__2184 (
            .O(N__9255),
            .I(N__9122));
    SRMux I__2183 (
            .O(N__9254),
            .I(N__9122));
    SRMux I__2182 (
            .O(N__9253),
            .I(N__9122));
    Glb2LocalMux I__2181 (
            .O(N__9250),
            .I(N__9122));
    SRMux I__2180 (
            .O(N__9249),
            .I(N__9122));
    SRMux I__2179 (
            .O(N__9248),
            .I(N__9122));
    SRMux I__2178 (
            .O(N__9247),
            .I(N__9122));
    SRMux I__2177 (
            .O(N__9246),
            .I(N__9122));
    SRMux I__2176 (
            .O(N__9245),
            .I(N__9122));
    SRMux I__2175 (
            .O(N__9244),
            .I(N__9122));
    SRMux I__2174 (
            .O(N__9243),
            .I(N__9122));
    Glb2LocalMux I__2173 (
            .O(N__9240),
            .I(N__9122));
    SRMux I__2172 (
            .O(N__9239),
            .I(N__9122));
    SRMux I__2171 (
            .O(N__9238),
            .I(N__9122));
    SRMux I__2170 (
            .O(N__9237),
            .I(N__9122));
    SRMux I__2169 (
            .O(N__9236),
            .I(N__9122));
    SRMux I__2168 (
            .O(N__9235),
            .I(N__9122));
    SRMux I__2167 (
            .O(N__9234),
            .I(N__9122));
    SRMux I__2166 (
            .O(N__9233),
            .I(N__9122));
    SRMux I__2165 (
            .O(N__9232),
            .I(N__9122));
    SRMux I__2164 (
            .O(N__9231),
            .I(N__9122));
    SRMux I__2163 (
            .O(N__9230),
            .I(N__9122));
    SRMux I__2162 (
            .O(N__9229),
            .I(N__9122));
    SRMux I__2161 (
            .O(N__9228),
            .I(N__9122));
    SRMux I__2160 (
            .O(N__9227),
            .I(N__9122));
    Glb2LocalMux I__2159 (
            .O(N__9224),
            .I(N__9122));
    SRMux I__2158 (
            .O(N__9223),
            .I(N__9122));
    SRMux I__2157 (
            .O(N__9222),
            .I(N__9122));
    SRMux I__2156 (
            .O(N__9221),
            .I(N__9122));
    Glb2LocalMux I__2155 (
            .O(N__9218),
            .I(N__9122));
    SRMux I__2154 (
            .O(N__9217),
            .I(N__9122));
    SRMux I__2153 (
            .O(N__9216),
            .I(N__9122));
    Glb2LocalMux I__2152 (
            .O(N__9213),
            .I(N__9122));
    GlobalMux I__2151 (
            .O(N__9122),
            .I(N__9119));
    gio2CtrlBuf I__2150 (
            .O(N__9119),
            .I(RESETn_c_i_g));
    InMux I__2149 (
            .O(N__9116),
            .I(N__9113));
    LocalMux I__2148 (
            .O(N__9113),
            .I(N__9109));
    InMux I__2147 (
            .O(N__9112),
            .I(N__9106));
    Sp12to4 I__2146 (
            .O(N__9109),
            .I(N__9101));
    LocalMux I__2145 (
            .O(N__9106),
            .I(N__9101));
    Span12Mux_v I__2144 (
            .O(N__9101),
            .I(N__9098));
    Span12Mux_h I__2143 (
            .O(N__9098),
            .I(N__9095));
    Odrv12 I__2142 (
            .O(N__9095),
            .I(DRA_c_6));
    InMux I__2141 (
            .O(N__9092),
            .I(N__9089));
    LocalMux I__2140 (
            .O(N__9089),
            .I(N__9086));
    Span4Mux_v I__2139 (
            .O(N__9086),
            .I(N__9083));
    Odrv4 I__2138 (
            .O(N__9083),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2137 (
            .O(N__9080),
            .I(N__9077));
    LocalMux I__2136 (
            .O(N__9077),
            .I(N__9073));
    InMux I__2135 (
            .O(N__9076),
            .I(N__9070));
    Span4Mux_h I__2134 (
            .O(N__9073),
            .I(N__9065));
    LocalMux I__2133 (
            .O(N__9070),
            .I(N__9065));
    Span4Mux_v I__2132 (
            .O(N__9065),
            .I(N__9062));
    Sp12to4 I__2131 (
            .O(N__9062),
            .I(N__9059));
    Span12Mux_h I__2130 (
            .O(N__9059),
            .I(N__9056));
    Span12Mux_v I__2129 (
            .O(N__9056),
            .I(N__9053));
    Odrv12 I__2128 (
            .O(N__9053),
            .I(DRA_c_4));
    InMux I__2127 (
            .O(N__9050),
            .I(N__9047));
    LocalMux I__2126 (
            .O(N__9047),
            .I(N__9044));
    Span4Mux_h I__2125 (
            .O(N__9044),
            .I(N__9041));
    Odrv4 I__2124 (
            .O(N__9041),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2123 (
            .O(N__9038),
            .I(N__9035));
    LocalMux I__2122 (
            .O(N__9035),
            .I(N__9032));
    Span4Mux_h I__2121 (
            .O(N__9032),
            .I(N__9029));
    Odrv4 I__2120 (
            .O(N__9029),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2119 (
            .O(N__9026),
            .I(N__9023));
    LocalMux I__2118 (
            .O(N__9023),
            .I(N__9020));
    Odrv4 I__2117 (
            .O(N__9020),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    CascadeMux I__2116 (
            .O(N__9017),
            .I(N__9014));
    InMux I__2115 (
            .O(N__9014),
            .I(N__9011));
    LocalMux I__2114 (
            .O(N__9011),
            .I(N__9008));
    Span4Mux_h I__2113 (
            .O(N__9008),
            .I(N__9005));
    Odrv4 I__2112 (
            .O(N__9005),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2111 (
            .O(N__9002),
            .I(N__8999));
    LocalMux I__2110 (
            .O(N__8999),
            .I(N__8995));
    InMux I__2109 (
            .O(N__8998),
            .I(N__8992));
    Sp12to4 I__2108 (
            .O(N__8995),
            .I(N__8987));
    LocalMux I__2107 (
            .O(N__8992),
            .I(N__8987));
    Span12Mux_v I__2106 (
            .O(N__8987),
            .I(N__8984));
    Span12Mux_h I__2105 (
            .O(N__8984),
            .I(N__8981));
    Odrv12 I__2104 (
            .O(N__8981),
            .I(DRA_c_2));
    InMux I__2103 (
            .O(N__8978),
            .I(N__8972));
    InMux I__2102 (
            .O(N__8977),
            .I(N__8972));
    LocalMux I__2101 (
            .O(N__8972),
            .I(N__8969));
    Span4Mux_h I__2100 (
            .O(N__8969),
            .I(N__8966));
    Odrv4 I__2099 (
            .O(N__8966),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__2098 (
            .O(N__8963),
            .I(N__8959));
    InMux I__2097 (
            .O(N__8962),
            .I(N__8956));
    LocalMux I__2096 (
            .O(N__8959),
            .I(N__8951));
    LocalMux I__2095 (
            .O(N__8956),
            .I(N__8951));
    Span12Mux_v I__2094 (
            .O(N__8951),
            .I(N__8948));
    Span12Mux_h I__2093 (
            .O(N__8948),
            .I(N__8945));
    Span12Mux_v I__2092 (
            .O(N__8945),
            .I(N__8942));
    Odrv12 I__2091 (
            .O(N__8942),
            .I(DRA_c_9));
    InMux I__2090 (
            .O(N__8939),
            .I(N__8936));
    LocalMux I__2089 (
            .O(N__8936),
            .I(N__8933));
    Span12Mux_v I__2088 (
            .O(N__8933),
            .I(N__8930));
    Odrv12 I__2087 (
            .O(N__8930),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    CEMux I__2086 (
            .O(N__8927),
            .I(N__8924));
    LocalMux I__2085 (
            .O(N__8924),
            .I(N__8917));
    CEMux I__2084 (
            .O(N__8923),
            .I(N__8914));
    CEMux I__2083 (
            .O(N__8922),
            .I(N__8911));
    CEMux I__2082 (
            .O(N__8921),
            .I(N__8908));
    CEMux I__2081 (
            .O(N__8920),
            .I(N__8905));
    Span4Mux_h I__2080 (
            .O(N__8917),
            .I(N__8899));
    LocalMux I__2079 (
            .O(N__8914),
            .I(N__8899));
    LocalMux I__2078 (
            .O(N__8911),
            .I(N__8896));
    LocalMux I__2077 (
            .O(N__8908),
            .I(N__8893));
    LocalMux I__2076 (
            .O(N__8905),
            .I(N__8890));
    CEMux I__2075 (
            .O(N__8904),
            .I(N__8887));
    Span4Mux_v I__2074 (
            .O(N__8899),
            .I(N__8884));
    Span4Mux_v I__2073 (
            .O(N__8896),
            .I(N__8875));
    Span4Mux_h I__2072 (
            .O(N__8893),
            .I(N__8875));
    Span4Mux_v I__2071 (
            .O(N__8890),
            .I(N__8875));
    LocalMux I__2070 (
            .O(N__8887),
            .I(N__8875));
    Odrv4 I__2069 (
            .O(N__8884),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ));
    Odrv4 I__2068 (
            .O(N__8875),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ));
    InMux I__2067 (
            .O(N__8870),
            .I(N__8867));
    LocalMux I__2066 (
            .O(N__8867),
            .I(N__8864));
    Span4Mux_v I__2065 (
            .O(N__8864),
            .I(N__8861));
    Sp12to4 I__2064 (
            .O(N__8861),
            .I(N__8858));
    Span12Mux_h I__2063 (
            .O(N__8858),
            .I(N__8855));
    Odrv12 I__2062 (
            .O(N__8855),
            .I(RAS0n_c));
    InMux I__2061 (
            .O(N__8852),
            .I(N__8849));
    LocalMux I__2060 (
            .O(N__8849),
            .I(N__8846));
    Span4Mux_v I__2059 (
            .O(N__8846),
            .I(N__8843));
    Odrv4 I__2058 (
            .O(N__8843),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    InMux I__2057 (
            .O(N__8840),
            .I(N__8837));
    LocalMux I__2056 (
            .O(N__8837),
            .I(N__8810));
    ClkMux I__2055 (
            .O(N__8836),
            .I(N__8732));
    ClkMux I__2054 (
            .O(N__8835),
            .I(N__8732));
    ClkMux I__2053 (
            .O(N__8834),
            .I(N__8732));
    ClkMux I__2052 (
            .O(N__8833),
            .I(N__8732));
    ClkMux I__2051 (
            .O(N__8832),
            .I(N__8732));
    ClkMux I__2050 (
            .O(N__8831),
            .I(N__8732));
    ClkMux I__2049 (
            .O(N__8830),
            .I(N__8732));
    ClkMux I__2048 (
            .O(N__8829),
            .I(N__8732));
    ClkMux I__2047 (
            .O(N__8828),
            .I(N__8732));
    ClkMux I__2046 (
            .O(N__8827),
            .I(N__8732));
    ClkMux I__2045 (
            .O(N__8826),
            .I(N__8732));
    ClkMux I__2044 (
            .O(N__8825),
            .I(N__8732));
    ClkMux I__2043 (
            .O(N__8824),
            .I(N__8732));
    ClkMux I__2042 (
            .O(N__8823),
            .I(N__8732));
    ClkMux I__2041 (
            .O(N__8822),
            .I(N__8732));
    ClkMux I__2040 (
            .O(N__8821),
            .I(N__8732));
    ClkMux I__2039 (
            .O(N__8820),
            .I(N__8732));
    ClkMux I__2038 (
            .O(N__8819),
            .I(N__8732));
    ClkMux I__2037 (
            .O(N__8818),
            .I(N__8732));
    ClkMux I__2036 (
            .O(N__8817),
            .I(N__8732));
    ClkMux I__2035 (
            .O(N__8816),
            .I(N__8732));
    ClkMux I__2034 (
            .O(N__8815),
            .I(N__8732));
    ClkMux I__2033 (
            .O(N__8814),
            .I(N__8732));
    ClkMux I__2032 (
            .O(N__8813),
            .I(N__8732));
    Glb2LocalMux I__2031 (
            .O(N__8810),
            .I(N__8732));
    ClkMux I__2030 (
            .O(N__8809),
            .I(N__8732));
    ClkMux I__2029 (
            .O(N__8808),
            .I(N__8732));
    ClkMux I__2028 (
            .O(N__8807),
            .I(N__8732));
    ClkMux I__2027 (
            .O(N__8806),
            .I(N__8732));
    ClkMux I__2026 (
            .O(N__8805),
            .I(N__8732));
    ClkMux I__2025 (
            .O(N__8804),
            .I(N__8732));
    ClkMux I__2024 (
            .O(N__8803),
            .I(N__8732));
    ClkMux I__2023 (
            .O(N__8802),
            .I(N__8732));
    ClkMux I__2022 (
            .O(N__8801),
            .I(N__8732));
    GlobalMux I__2021 (
            .O(N__8732),
            .I(CLK80_PLL));
    CEMux I__2020 (
            .O(N__8729),
            .I(N__8726));
    LocalMux I__2019 (
            .O(N__8726),
            .I(N__8721));
    CEMux I__2018 (
            .O(N__8725),
            .I(N__8718));
    CEMux I__2017 (
            .O(N__8724),
            .I(N__8715));
    Span4Mux_h I__2016 (
            .O(N__8721),
            .I(N__8712));
    LocalMux I__2015 (
            .O(N__8718),
            .I(N__8708));
    LocalMux I__2014 (
            .O(N__8715),
            .I(N__8705));
    Span4Mux_h I__2013 (
            .O(N__8712),
            .I(N__8700));
    CEMux I__2012 (
            .O(N__8711),
            .I(N__8697));
    Span12Mux_h I__2011 (
            .O(N__8708),
            .I(N__8692));
    Sp12to4 I__2010 (
            .O(N__8705),
            .I(N__8692));
    CEMux I__2009 (
            .O(N__8704),
            .I(N__8689));
    CEMux I__2008 (
            .O(N__8703),
            .I(N__8686));
    Odrv4 I__2007 (
            .O(N__8700),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__2006 (
            .O(N__8697),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv12 I__2005 (
            .O(N__8692),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__2004 (
            .O(N__8689),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__2003 (
            .O(N__8686),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    InMux I__2002 (
            .O(N__8675),
            .I(N__8672));
    LocalMux I__2001 (
            .O(N__8672),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2000 (
            .O(N__8669),
            .I(N__8663));
    InMux I__1999 (
            .O(N__8668),
            .I(N__8663));
    LocalMux I__1998 (
            .O(N__8663),
            .I(N__8660));
    Odrv4 I__1997 (
            .O(N__8660),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1996 (
            .O(N__8657),
            .I(N__8654));
    LocalMux I__1995 (
            .O(N__8654),
            .I(N__8650));
    InMux I__1994 (
            .O(N__8653),
            .I(N__8647));
    Span4Mux_h I__1993 (
            .O(N__8650),
            .I(N__8642));
    LocalMux I__1992 (
            .O(N__8647),
            .I(N__8642));
    Sp12to4 I__1991 (
            .O(N__8642),
            .I(N__8639));
    Span12Mux_v I__1990 (
            .O(N__8639),
            .I(N__8636));
    Span12Mux_h I__1989 (
            .O(N__8636),
            .I(N__8633));
    Odrv12 I__1988 (
            .O(N__8633),
            .I(DRA_c_5));
    InMux I__1987 (
            .O(N__8630),
            .I(N__8627));
    LocalMux I__1986 (
            .O(N__8627),
            .I(N__8624));
    Span4Mux_h I__1985 (
            .O(N__8624),
            .I(N__8621));
    Odrv4 I__1984 (
            .O(N__8621),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1983 (
            .O(N__8618),
            .I(N__8614));
    InMux I__1982 (
            .O(N__8617),
            .I(N__8611));
    LocalMux I__1981 (
            .O(N__8614),
            .I(N__8606));
    LocalMux I__1980 (
            .O(N__8611),
            .I(N__8606));
    Span4Mux_v I__1979 (
            .O(N__8606),
            .I(N__8603));
    Sp12to4 I__1978 (
            .O(N__8603),
            .I(N__8600));
    Span12Mux_h I__1977 (
            .O(N__8600),
            .I(N__8597));
    Odrv12 I__1976 (
            .O(N__8597),
            .I(DRA_c_7));
    InMux I__1975 (
            .O(N__8594),
            .I(N__8591));
    LocalMux I__1974 (
            .O(N__8591),
            .I(N__8588));
    Odrv4 I__1973 (
            .O(N__8588),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__1972 (
            .O(N__8585),
            .I(N__8582));
    LocalMux I__1971 (
            .O(N__8582),
            .I(N__8579));
    Span4Mux_h I__1970 (
            .O(N__8579),
            .I(N__8576));
    Odrv4 I__1969 (
            .O(N__8576),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1968 (
            .O(N__8573),
            .I(N__8570));
    LocalMux I__1967 (
            .O(N__8570),
            .I(N__8567));
    Span4Mux_h I__1966 (
            .O(N__8567),
            .I(N__8564));
    Span4Mux_v I__1965 (
            .O(N__8564),
            .I(N__8561));
    Odrv4 I__1964 (
            .O(N__8561),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__1963 (
            .O(N__8558),
            .I(N__8554));
    InMux I__1962 (
            .O(N__8557),
            .I(N__8551));
    LocalMux I__1961 (
            .O(N__8554),
            .I(N__8546));
    LocalMux I__1960 (
            .O(N__8551),
            .I(N__8546));
    Sp12to4 I__1959 (
            .O(N__8546),
            .I(N__8543));
    Span12Mux_v I__1958 (
            .O(N__8543),
            .I(N__8540));
    Span12Mux_h I__1957 (
            .O(N__8540),
            .I(N__8537));
    Odrv12 I__1956 (
            .O(N__8537),
            .I(DRA_c_1));
    InMux I__1955 (
            .O(N__8534),
            .I(N__8531));
    LocalMux I__1954 (
            .O(N__8531),
            .I(N__8528));
    Span4Mux_v I__1953 (
            .O(N__8528),
            .I(N__8525));
    Span4Mux_h I__1952 (
            .O(N__8525),
            .I(N__8522));
    Odrv4 I__1951 (
            .O(N__8522),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__1950 (
            .O(N__8519),
            .I(N__8514));
    InMux I__1949 (
            .O(N__8518),
            .I(N__8511));
    InMux I__1948 (
            .O(N__8517),
            .I(N__8508));
    LocalMux I__1947 (
            .O(N__8514),
            .I(N__8503));
    LocalMux I__1946 (
            .O(N__8511),
            .I(N__8503));
    LocalMux I__1945 (
            .O(N__8508),
            .I(N__8500));
    Span4Mux_v I__1944 (
            .O(N__8503),
            .I(N__8497));
    Span4Mux_v I__1943 (
            .O(N__8500),
            .I(N__8494));
    Sp12to4 I__1942 (
            .O(N__8497),
            .I(N__8489));
    Sp12to4 I__1941 (
            .O(N__8494),
            .I(N__8489));
    Span12Mux_h I__1940 (
            .O(N__8489),
            .I(N__8486));
    Span12Mux_v I__1939 (
            .O(N__8486),
            .I(N__8483));
    Odrv12 I__1938 (
            .O(N__8483),
            .I(DBRn_c));
    InMux I__1937 (
            .O(N__8480),
            .I(N__8477));
    LocalMux I__1936 (
            .O(N__8477),
            .I(N__8467));
    ClkMux I__1935 (
            .O(N__8476),
            .I(N__8450));
    ClkMux I__1934 (
            .O(N__8475),
            .I(N__8450));
    ClkMux I__1933 (
            .O(N__8474),
            .I(N__8450));
    ClkMux I__1932 (
            .O(N__8473),
            .I(N__8450));
    ClkMux I__1931 (
            .O(N__8472),
            .I(N__8450));
    ClkMux I__1930 (
            .O(N__8471),
            .I(N__8450));
    ClkMux I__1929 (
            .O(N__8470),
            .I(N__8450));
    Glb2LocalMux I__1928 (
            .O(N__8467),
            .I(N__8450));
    GlobalMux I__1927 (
            .O(N__8450),
            .I(N__8447));
    gio2CtrlBuf I__1926 (
            .O(N__8447),
            .I(C1_c_g));
    InMux I__1925 (
            .O(N__8444),
            .I(N__8440));
    InMux I__1924 (
            .O(N__8443),
            .I(N__8430));
    LocalMux I__1923 (
            .O(N__8440),
            .I(N__8426));
    InMux I__1922 (
            .O(N__8439),
            .I(N__8417));
    InMux I__1921 (
            .O(N__8438),
            .I(N__8417));
    InMux I__1920 (
            .O(N__8437),
            .I(N__8417));
    InMux I__1919 (
            .O(N__8436),
            .I(N__8417));
    InMux I__1918 (
            .O(N__8435),
            .I(N__8414));
    InMux I__1917 (
            .O(N__8434),
            .I(N__8411));
    InMux I__1916 (
            .O(N__8433),
            .I(N__8408));
    LocalMux I__1915 (
            .O(N__8430),
            .I(N__8405));
    InMux I__1914 (
            .O(N__8429),
            .I(N__8402));
    Span4Mux_v I__1913 (
            .O(N__8426),
            .I(N__8395));
    LocalMux I__1912 (
            .O(N__8417),
            .I(N__8395));
    LocalMux I__1911 (
            .O(N__8414),
            .I(N__8395));
    LocalMux I__1910 (
            .O(N__8411),
            .I(N__8391));
    LocalMux I__1909 (
            .O(N__8408),
            .I(N__8388));
    Span4Mux_v I__1908 (
            .O(N__8405),
            .I(N__8385));
    LocalMux I__1907 (
            .O(N__8402),
            .I(N__8380));
    Span4Mux_v I__1906 (
            .O(N__8395),
            .I(N__8380));
    InMux I__1905 (
            .O(N__8394),
            .I(N__8377));
    Span12Mux_v I__1904 (
            .O(N__8391),
            .I(N__8374));
    Span12Mux_v I__1903 (
            .O(N__8388),
            .I(N__8365));
    Sp12to4 I__1902 (
            .O(N__8385),
            .I(N__8365));
    Sp12to4 I__1901 (
            .O(N__8380),
            .I(N__8365));
    LocalMux I__1900 (
            .O(N__8377),
            .I(N__8365));
    Span12Mux_h I__1899 (
            .O(N__8374),
            .I(N__8362));
    Span12Mux_h I__1898 (
            .O(N__8365),
            .I(N__8359));
    Odrv12 I__1897 (
            .O(N__8362),
            .I(RESETn_c));
    Odrv12 I__1896 (
            .O(N__8359),
            .I(RESETn_c));
    IoInMux I__1895 (
            .O(N__8354),
            .I(N__8351));
    LocalMux I__1894 (
            .O(N__8351),
            .I(N__8348));
    Span12Mux_s4_v I__1893 (
            .O(N__8348),
            .I(N__8345));
    Odrv12 I__1892 (
            .O(N__8345),
            .I(RESETn_c_i));
    IoInMux I__1891 (
            .O(N__8342),
            .I(N__8339));
    LocalMux I__1890 (
            .O(N__8339),
            .I(N__8336));
    Span12Mux_s10_v I__1889 (
            .O(N__8336),
            .I(N__8333));
    Span12Mux_h I__1888 (
            .O(N__8333),
            .I(N__8330));
    Odrv12 I__1887 (
            .O(N__8330),
            .I(N_118));
    InMux I__1886 (
            .O(N__8327),
            .I(N__8319));
    InMux I__1885 (
            .O(N__8326),
            .I(N__8319));
    InMux I__1884 (
            .O(N__8325),
            .I(N__8314));
    InMux I__1883 (
            .O(N__8324),
            .I(N__8314));
    LocalMux I__1882 (
            .O(N__8319),
            .I(N__8309));
    LocalMux I__1881 (
            .O(N__8314),
            .I(N__8306));
    InMux I__1880 (
            .O(N__8313),
            .I(N__8301));
    InMux I__1879 (
            .O(N__8312),
            .I(N__8301));
    Span4Mux_v I__1878 (
            .O(N__8309),
            .I(N__8298));
    Span4Mux_v I__1877 (
            .O(N__8306),
            .I(N__8295));
    LocalMux I__1876 (
            .O(N__8301),
            .I(N__8292));
    Span4Mux_h I__1875 (
            .O(N__8298),
            .I(N__8289));
    Span4Mux_h I__1874 (
            .O(N__8295),
            .I(N__8284));
    Span4Mux_v I__1873 (
            .O(N__8292),
            .I(N__8284));
    Sp12to4 I__1872 (
            .O(N__8289),
            .I(N__8279));
    Sp12to4 I__1871 (
            .O(N__8284),
            .I(N__8279));
    Odrv12 I__1870 (
            .O(N__8279),
            .I(A_c_0));
    InMux I__1869 (
            .O(N__8276),
            .I(N__8272));
    CascadeMux I__1868 (
            .O(N__8275),
            .I(N__8269));
    LocalMux I__1867 (
            .O(N__8272),
            .I(N__8265));
    InMux I__1866 (
            .O(N__8269),
            .I(N__8260));
    InMux I__1865 (
            .O(N__8268),
            .I(N__8260));
    Span4Mux_h I__1864 (
            .O(N__8265),
            .I(N__8257));
    LocalMux I__1863 (
            .O(N__8260),
            .I(N__8254));
    Sp12to4 I__1862 (
            .O(N__8257),
            .I(N__8251));
    Span12Mux_v I__1861 (
            .O(N__8254),
            .I(N__8248));
    Span12Mux_v I__1860 (
            .O(N__8251),
            .I(N__8245));
    Span12Mux_h I__1859 (
            .O(N__8248),
            .I(N__8242));
    Odrv12 I__1858 (
            .O(N__8245),
            .I(SIZ_c_0));
    Odrv12 I__1857 (
            .O(N__8242),
            .I(SIZ_c_0));
    InMux I__1856 (
            .O(N__8237),
            .I(N__8231));
    InMux I__1855 (
            .O(N__8236),
            .I(N__8231));
    LocalMux I__1854 (
            .O(N__8231),
            .I(N__8228));
    Span12Mux_s9_v I__1853 (
            .O(N__8228),
            .I(N__8224));
    InMux I__1852 (
            .O(N__8227),
            .I(N__8221));
    Odrv12 I__1851 (
            .O(N__8224),
            .I(DS_ENm));
    LocalMux I__1850 (
            .O(N__8221),
            .I(DS_ENm));
    IoInMux I__1849 (
            .O(N__8216),
            .I(N__8213));
    LocalMux I__1848 (
            .O(N__8213),
            .I(N__8210));
    Span4Mux_s3_v I__1847 (
            .O(N__8210),
            .I(N__8207));
    Span4Mux_v I__1846 (
            .O(N__8207),
            .I(N__8204));
    Sp12to4 I__1845 (
            .O(N__8204),
            .I(N__8201));
    Odrv12 I__1844 (
            .O(N__8201),
            .I(N_113));
    InMux I__1843 (
            .O(N__8198),
            .I(N__8195));
    LocalMux I__1842 (
            .O(N__8195),
            .I(N__8191));
    InMux I__1841 (
            .O(N__8194),
            .I(N__8188));
    Span4Mux_v I__1840 (
            .O(N__8191),
            .I(N__8182));
    LocalMux I__1839 (
            .O(N__8188),
            .I(N__8182));
    CascadeMux I__1838 (
            .O(N__8187),
            .I(N__8178));
    Span4Mux_v I__1837 (
            .O(N__8182),
            .I(N__8175));
    InMux I__1836 (
            .O(N__8181),
            .I(N__8172));
    InMux I__1835 (
            .O(N__8178),
            .I(N__8169));
    Odrv4 I__1834 (
            .O(N__8175),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1833 (
            .O(N__8172),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1832 (
            .O(N__8169),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1831 (
            .O(N__8162),
            .I(N__8159));
    LocalMux I__1830 (
            .O(N__8159),
            .I(N__8156));
    Span4Mux_s2_v I__1829 (
            .O(N__8156),
            .I(N__8153));
    Span4Mux_v I__1828 (
            .O(N__8153),
            .I(N__8150));
    Span4Mux_h I__1827 (
            .O(N__8150),
            .I(N__8147));
    Odrv4 I__1826 (
            .O(N__8147),
            .I(CRCSn_c));
    CascadeMux I__1825 (
            .O(N__8144),
            .I(N__8141));
    InMux I__1824 (
            .O(N__8141),
            .I(N__8137));
    InMux I__1823 (
            .O(N__8140),
            .I(N__8134));
    LocalMux I__1822 (
            .O(N__8137),
            .I(N__8128));
    LocalMux I__1821 (
            .O(N__8134),
            .I(N__8123));
    InMux I__1820 (
            .O(N__8133),
            .I(N__8118));
    InMux I__1819 (
            .O(N__8132),
            .I(N__8118));
    InMux I__1818 (
            .O(N__8131),
            .I(N__8115));
    Span4Mux_v I__1817 (
            .O(N__8128),
            .I(N__8112));
    InMux I__1816 (
            .O(N__8127),
            .I(N__8107));
    InMux I__1815 (
            .O(N__8126),
            .I(N__8107));
    Span4Mux_h I__1814 (
            .O(N__8123),
            .I(N__8102));
    LocalMux I__1813 (
            .O(N__8118),
            .I(N__8102));
    LocalMux I__1812 (
            .O(N__8115),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1811 (
            .O(N__8112),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1810 (
            .O(N__8107),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1809 (
            .O(N__8102),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1808 (
            .O(N__8093),
            .I(N__8090));
    LocalMux I__1807 (
            .O(N__8090),
            .I(N__8087));
    IoSpan4Mux I__1806 (
            .O(N__8087),
            .I(N__8084));
    Span4Mux_s2_h I__1805 (
            .O(N__8084),
            .I(N__8081));
    Sp12to4 I__1804 (
            .O(N__8081),
            .I(N__8078));
    Span12Mux_h I__1803 (
            .O(N__8078),
            .I(N__8075));
    Odrv12 I__1802 (
            .O(N__8075),
            .I(WEn_c));
    InMux I__1801 (
            .O(N__8072),
            .I(N__8068));
    InMux I__1800 (
            .O(N__8071),
            .I(N__8065));
    LocalMux I__1799 (
            .O(N__8068),
            .I(N__8060));
    LocalMux I__1798 (
            .O(N__8065),
            .I(N__8057));
    InMux I__1797 (
            .O(N__8064),
            .I(N__8052));
    InMux I__1796 (
            .O(N__8063),
            .I(N__8052));
    Span4Mux_v I__1795 (
            .O(N__8060),
            .I(N__8047));
    Span4Mux_v I__1794 (
            .O(N__8057),
            .I(N__8042));
    LocalMux I__1793 (
            .O(N__8052),
            .I(N__8042));
    InMux I__1792 (
            .O(N__8051),
            .I(N__8037));
    InMux I__1791 (
            .O(N__8050),
            .I(N__8037));
    Odrv4 I__1790 (
            .O(N__8047),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1789 (
            .O(N__8042),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1788 (
            .O(N__8037),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__1787 (
            .O(N__8030),
            .I(N__8027));
    LocalMux I__1786 (
            .O(N__8027),
            .I(N__8024));
    Span4Mux_s2_v I__1785 (
            .O(N__8024),
            .I(N__8021));
    Span4Mux_v I__1784 (
            .O(N__8021),
            .I(N__8018));
    Span4Mux_v I__1783 (
            .O(N__8018),
            .I(N__8015));
    Span4Mux_h I__1782 (
            .O(N__8015),
            .I(N__8012));
    Odrv4 I__1781 (
            .O(N__8012),
            .I(RASn_c));
    InMux I__1780 (
            .O(N__8009),
            .I(N__8006));
    LocalMux I__1779 (
            .O(N__8006),
            .I(N__8003));
    Span4Mux_v I__1778 (
            .O(N__8003),
            .I(N__8000));
    Span4Mux_v I__1777 (
            .O(N__8000),
            .I(N__7997));
    Sp12to4 I__1776 (
            .O(N__7997),
            .I(N__7994));
    Span12Mux_h I__1775 (
            .O(N__7994),
            .I(N__7991));
    Odrv12 I__1774 (
            .O(N__7991),
            .I(A_c_19));
    IoInMux I__1773 (
            .O(N__7988),
            .I(N__7985));
    LocalMux I__1772 (
            .O(N__7985),
            .I(N__7982));
    IoSpan4Mux I__1771 (
            .O(N__7982),
            .I(N__7979));
    Span4Mux_s1_h I__1770 (
            .O(N__7979),
            .I(N__7976));
    Sp12to4 I__1769 (
            .O(N__7976),
            .I(N__7973));
    Span12Mux_h I__1768 (
            .O(N__7973),
            .I(N__7970));
    Odrv12 I__1767 (
            .O(N__7970),
            .I(CMA_c_9));
    InMux I__1766 (
            .O(N__7967),
            .I(N__7960));
    InMux I__1765 (
            .O(N__7966),
            .I(N__7960));
    CascadeMux I__1764 (
            .O(N__7965),
            .I(N__7957));
    LocalMux I__1763 (
            .O(N__7960),
            .I(N__7953));
    InMux I__1762 (
            .O(N__7957),
            .I(N__7948));
    InMux I__1761 (
            .O(N__7956),
            .I(N__7948));
    Odrv4 I__1760 (
            .O(N__7953),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1759 (
            .O(N__7948),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    InMux I__1758 (
            .O(N__7943),
            .I(N__7940));
    LocalMux I__1757 (
            .O(N__7940),
            .I(N__7937));
    Span4Mux_v I__1756 (
            .O(N__7937),
            .I(N__7934));
    Span4Mux_v I__1755 (
            .O(N__7934),
            .I(N__7931));
    Sp12to4 I__1754 (
            .O(N__7931),
            .I(N__7928));
    Span12Mux_h I__1753 (
            .O(N__7928),
            .I(N__7925));
    Odrv12 I__1752 (
            .O(N__7925),
            .I(A_c_17));
    CascadeMux I__1751 (
            .O(N__7922),
            .I(N__7915));
    InMux I__1750 (
            .O(N__7921),
            .I(N__7907));
    InMux I__1749 (
            .O(N__7920),
            .I(N__7904));
    CascadeMux I__1748 (
            .O(N__7919),
            .I(N__7899));
    InMux I__1747 (
            .O(N__7918),
            .I(N__7891));
    InMux I__1746 (
            .O(N__7915),
            .I(N__7891));
    CascadeMux I__1745 (
            .O(N__7914),
            .I(N__7881));
    CascadeMux I__1744 (
            .O(N__7913),
            .I(N__7878));
    InMux I__1743 (
            .O(N__7912),
            .I(N__7875));
    InMux I__1742 (
            .O(N__7911),
            .I(N__7870));
    InMux I__1741 (
            .O(N__7910),
            .I(N__7870));
    LocalMux I__1740 (
            .O(N__7907),
            .I(N__7865));
    LocalMux I__1739 (
            .O(N__7904),
            .I(N__7865));
    InMux I__1738 (
            .O(N__7903),
            .I(N__7858));
    InMux I__1737 (
            .O(N__7902),
            .I(N__7858));
    InMux I__1736 (
            .O(N__7899),
            .I(N__7858));
    InMux I__1735 (
            .O(N__7898),
            .I(N__7853));
    InMux I__1734 (
            .O(N__7897),
            .I(N__7853));
    InMux I__1733 (
            .O(N__7896),
            .I(N__7850));
    LocalMux I__1732 (
            .O(N__7891),
            .I(N__7847));
    InMux I__1731 (
            .O(N__7890),
            .I(N__7840));
    InMux I__1730 (
            .O(N__7889),
            .I(N__7840));
    InMux I__1729 (
            .O(N__7888),
            .I(N__7840));
    InMux I__1728 (
            .O(N__7887),
            .I(N__7837));
    InMux I__1727 (
            .O(N__7886),
            .I(N__7832));
    InMux I__1726 (
            .O(N__7885),
            .I(N__7832));
    InMux I__1725 (
            .O(N__7884),
            .I(N__7825));
    InMux I__1724 (
            .O(N__7881),
            .I(N__7825));
    InMux I__1723 (
            .O(N__7878),
            .I(N__7825));
    LocalMux I__1722 (
            .O(N__7875),
            .I(N__7819));
    LocalMux I__1721 (
            .O(N__7870),
            .I(N__7819));
    Span4Mux_v I__1720 (
            .O(N__7865),
            .I(N__7812));
    LocalMux I__1719 (
            .O(N__7858),
            .I(N__7812));
    LocalMux I__1718 (
            .O(N__7853),
            .I(N__7812));
    LocalMux I__1717 (
            .O(N__7850),
            .I(N__7808));
    Span4Mux_v I__1716 (
            .O(N__7847),
            .I(N__7801));
    LocalMux I__1715 (
            .O(N__7840),
            .I(N__7801));
    LocalMux I__1714 (
            .O(N__7837),
            .I(N__7801));
    LocalMux I__1713 (
            .O(N__7832),
            .I(N__7798));
    LocalMux I__1712 (
            .O(N__7825),
            .I(N__7795));
    InMux I__1711 (
            .O(N__7824),
            .I(N__7792));
    Span4Mux_v I__1710 (
            .O(N__7819),
            .I(N__7789));
    Span4Mux_v I__1709 (
            .O(N__7812),
            .I(N__7786));
    InMux I__1708 (
            .O(N__7811),
            .I(N__7783));
    Span4Mux_v I__1707 (
            .O(N__7808),
            .I(N__7778));
    Span4Mux_h I__1706 (
            .O(N__7801),
            .I(N__7778));
    Odrv4 I__1705 (
            .O(N__7798),
            .I(CPU_CYCLEm));
    Odrv4 I__1704 (
            .O(N__7795),
            .I(CPU_CYCLEm));
    LocalMux I__1703 (
            .O(N__7792),
            .I(CPU_CYCLEm));
    Odrv4 I__1702 (
            .O(N__7789),
            .I(CPU_CYCLEm));
    Odrv4 I__1701 (
            .O(N__7786),
            .I(CPU_CYCLEm));
    LocalMux I__1700 (
            .O(N__7783),
            .I(CPU_CYCLEm));
    Odrv4 I__1699 (
            .O(N__7778),
            .I(CPU_CYCLEm));
    IoInMux I__1698 (
            .O(N__7763),
            .I(N__7760));
    LocalMux I__1697 (
            .O(N__7760),
            .I(N__7757));
    IoSpan4Mux I__1696 (
            .O(N__7757),
            .I(N__7754));
    Span4Mux_s2_h I__1695 (
            .O(N__7754),
            .I(N__7751));
    Sp12to4 I__1694 (
            .O(N__7751),
            .I(N__7748));
    Span12Mux_h I__1693 (
            .O(N__7748),
            .I(N__7745));
    Odrv12 I__1692 (
            .O(N__7745),
            .I(CMA_c_8));
    InMux I__1691 (
            .O(N__7742),
            .I(N__7738));
    InMux I__1690 (
            .O(N__7741),
            .I(N__7735));
    LocalMux I__1689 (
            .O(N__7738),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1688 (
            .O(N__7735),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    CascadeMux I__1687 (
            .O(N__7730),
            .I(N__7726));
    CascadeMux I__1686 (
            .O(N__7729),
            .I(N__7722));
    InMux I__1685 (
            .O(N__7726),
            .I(N__7717));
    InMux I__1684 (
            .O(N__7725),
            .I(N__7717));
    InMux I__1683 (
            .O(N__7722),
            .I(N__7714));
    LocalMux I__1682 (
            .O(N__7717),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__1681 (
            .O(N__7714),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    IoInMux I__1680 (
            .O(N__7709),
            .I(N__7705));
    IoInMux I__1679 (
            .O(N__7708),
            .I(N__7702));
    LocalMux I__1678 (
            .O(N__7705),
            .I(N__7699));
    LocalMux I__1677 (
            .O(N__7702),
            .I(N__7696));
    Span4Mux_s3_v I__1676 (
            .O(N__7699),
            .I(N__7693));
    Span4Mux_s2_v I__1675 (
            .O(N__7696),
            .I(N__7690));
    Sp12to4 I__1674 (
            .O(N__7693),
            .I(N__7687));
    Span4Mux_h I__1673 (
            .O(N__7690),
            .I(N__7684));
    Span12Mux_s11_h I__1672 (
            .O(N__7687),
            .I(N__7681));
    Sp12to4 I__1671 (
            .O(N__7684),
            .I(N__7678));
    Span12Mux_v I__1670 (
            .O(N__7681),
            .I(N__7672));
    Span12Mux_v I__1669 (
            .O(N__7678),
            .I(N__7672));
    InMux I__1668 (
            .O(N__7677),
            .I(N__7669));
    Odrv12 I__1667 (
            .O(N__7672),
            .I(ASn_c));
    LocalMux I__1666 (
            .O(N__7669),
            .I(ASn_c));
    InMux I__1665 (
            .O(N__7664),
            .I(N__7652));
    InMux I__1664 (
            .O(N__7663),
            .I(N__7652));
    InMux I__1663 (
            .O(N__7662),
            .I(N__7652));
    InMux I__1662 (
            .O(N__7661),
            .I(N__7652));
    LocalMux I__1661 (
            .O(N__7652),
            .I(\U712_REG_SM.STATE_COUNT_RNITQLC2Z0Z_1 ));
    InMux I__1660 (
            .O(N__7649),
            .I(N__7646));
    LocalMux I__1659 (
            .O(N__7646),
            .I(N__7643));
    Span4Mux_v I__1658 (
            .O(N__7643),
            .I(N__7640));
    Sp12to4 I__1657 (
            .O(N__7640),
            .I(N__7637));
    Span12Mux_h I__1656 (
            .O(N__7637),
            .I(N__7634));
    Span12Mux_v I__1655 (
            .O(N__7634),
            .I(N__7631));
    Odrv12 I__1654 (
            .O(N__7631),
            .I(REGSPACEn_c));
    CascadeMux I__1653 (
            .O(N__7628),
            .I(N__7624));
    InMux I__1652 (
            .O(N__7627),
            .I(N__7619));
    InMux I__1651 (
            .O(N__7624),
            .I(N__7619));
    LocalMux I__1650 (
            .O(N__7619),
            .I(\U712_REG_SM.REG_CYCLE_GOZ0 ));
    CascadeMux I__1649 (
            .O(N__7616),
            .I(N__7612));
    InMux I__1648 (
            .O(N__7615),
            .I(N__7609));
    InMux I__1647 (
            .O(N__7612),
            .I(N__7606));
    LocalMux I__1646 (
            .O(N__7609),
            .I(N__7603));
    LocalMux I__1645 (
            .O(N__7606),
            .I(N__7600));
    Span4Mux_v I__1644 (
            .O(N__7603),
            .I(N__7597));
    Span4Mux_v I__1643 (
            .O(N__7600),
            .I(N__7594));
    Sp12to4 I__1642 (
            .O(N__7597),
            .I(N__7589));
    Sp12to4 I__1641 (
            .O(N__7594),
            .I(N__7589));
    Span12Mux_h I__1640 (
            .O(N__7589),
            .I(N__7586));
    Span12Mux_v I__1639 (
            .O(N__7586),
            .I(N__7583));
    Odrv12 I__1638 (
            .O(N__7583),
            .I(TSn_c));
    InMux I__1637 (
            .O(N__7580),
            .I(N__7568));
    InMux I__1636 (
            .O(N__7579),
            .I(N__7568));
    InMux I__1635 (
            .O(N__7578),
            .I(N__7568));
    InMux I__1634 (
            .O(N__7577),
            .I(N__7568));
    LocalMux I__1633 (
            .O(N__7568),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    CascadeMux I__1632 (
            .O(N__7565),
            .I(N__7561));
    InMux I__1631 (
            .O(N__7564),
            .I(N__7556));
    InMux I__1630 (
            .O(N__7561),
            .I(N__7553));
    InMux I__1629 (
            .O(N__7560),
            .I(N__7548));
    InMux I__1628 (
            .O(N__7559),
            .I(N__7548));
    LocalMux I__1627 (
            .O(N__7556),
            .I(N__7545));
    LocalMux I__1626 (
            .O(N__7553),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa ));
    LocalMux I__1625 (
            .O(N__7548),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa ));
    Odrv12 I__1624 (
            .O(N__7545),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa ));
    InMux I__1623 (
            .O(N__7538),
            .I(N__7529));
    InMux I__1622 (
            .O(N__7537),
            .I(N__7529));
    InMux I__1621 (
            .O(N__7536),
            .I(N__7529));
    LocalMux I__1620 (
            .O(N__7529),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    CascadeMux I__1619 (
            .O(N__7526),
            .I(N__7521));
    InMux I__1618 (
            .O(N__7525),
            .I(N__7514));
    InMux I__1617 (
            .O(N__7524),
            .I(N__7514));
    InMux I__1616 (
            .O(N__7521),
            .I(N__7514));
    LocalMux I__1615 (
            .O(N__7514),
            .I(\U712_REG_SM.N_205 ));
    InMux I__1614 (
            .O(N__7511),
            .I(N__7507));
    InMux I__1613 (
            .O(N__7510),
            .I(N__7503));
    LocalMux I__1612 (
            .O(N__7507),
            .I(N__7500));
    InMux I__1611 (
            .O(N__7506),
            .I(N__7497));
    LocalMux I__1610 (
            .O(N__7503),
            .I(\U712_REG_SM.N_202 ));
    Odrv4 I__1609 (
            .O(N__7500),
            .I(\U712_REG_SM.N_202 ));
    LocalMux I__1608 (
            .O(N__7497),
            .I(\U712_REG_SM.N_202 ));
    CascadeMux I__1607 (
            .O(N__7490),
            .I(N__7485));
    InMux I__1606 (
            .O(N__7489),
            .I(N__7482));
    InMux I__1605 (
            .O(N__7488),
            .I(N__7479));
    InMux I__1604 (
            .O(N__7485),
            .I(N__7476));
    LocalMux I__1603 (
            .O(N__7482),
            .I(N__7473));
    LocalMux I__1602 (
            .O(N__7479),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1601 (
            .O(N__7476),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv12 I__1600 (
            .O(N__7473),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    InMux I__1599 (
            .O(N__7466),
            .I(N__7461));
    CascadeMux I__1598 (
            .O(N__7465),
            .I(N__7458));
    CascadeMux I__1597 (
            .O(N__7464),
            .I(N__7455));
    LocalMux I__1596 (
            .O(N__7461),
            .I(N__7442));
    InMux I__1595 (
            .O(N__7458),
            .I(N__7439));
    InMux I__1594 (
            .O(N__7455),
            .I(N__7436));
    CascadeMux I__1593 (
            .O(N__7454),
            .I(N__7433));
    InMux I__1592 (
            .O(N__7453),
            .I(N__7428));
    InMux I__1591 (
            .O(N__7452),
            .I(N__7425));
    InMux I__1590 (
            .O(N__7451),
            .I(N__7416));
    InMux I__1589 (
            .O(N__7450),
            .I(N__7416));
    InMux I__1588 (
            .O(N__7449),
            .I(N__7416));
    InMux I__1587 (
            .O(N__7448),
            .I(N__7416));
    InMux I__1586 (
            .O(N__7447),
            .I(N__7413));
    CascadeMux I__1585 (
            .O(N__7446),
            .I(N__7410));
    CascadeMux I__1584 (
            .O(N__7445),
            .I(N__7407));
    Span4Mux_v I__1583 (
            .O(N__7442),
            .I(N__7400));
    LocalMux I__1582 (
            .O(N__7439),
            .I(N__7400));
    LocalMux I__1581 (
            .O(N__7436),
            .I(N__7400));
    InMux I__1580 (
            .O(N__7433),
            .I(N__7397));
    InMux I__1579 (
            .O(N__7432),
            .I(N__7392));
    CascadeMux I__1578 (
            .O(N__7431),
            .I(N__7388));
    LocalMux I__1577 (
            .O(N__7428),
            .I(N__7383));
    LocalMux I__1576 (
            .O(N__7425),
            .I(N__7380));
    LocalMux I__1575 (
            .O(N__7416),
            .I(N__7377));
    LocalMux I__1574 (
            .O(N__7413),
            .I(N__7374));
    InMux I__1573 (
            .O(N__7410),
            .I(N__7369));
    InMux I__1572 (
            .O(N__7407),
            .I(N__7369));
    Span4Mux_h I__1571 (
            .O(N__7400),
            .I(N__7363));
    LocalMux I__1570 (
            .O(N__7397),
            .I(N__7360));
    InMux I__1569 (
            .O(N__7396),
            .I(N__7355));
    InMux I__1568 (
            .O(N__7395),
            .I(N__7355));
    LocalMux I__1567 (
            .O(N__7392),
            .I(N__7352));
    InMux I__1566 (
            .O(N__7391),
            .I(N__7349));
    InMux I__1565 (
            .O(N__7388),
            .I(N__7342));
    InMux I__1564 (
            .O(N__7387),
            .I(N__7342));
    InMux I__1563 (
            .O(N__7386),
            .I(N__7342));
    Span4Mux_v I__1562 (
            .O(N__7383),
            .I(N__7331));
    Span4Mux_v I__1561 (
            .O(N__7380),
            .I(N__7331));
    Span4Mux_v I__1560 (
            .O(N__7377),
            .I(N__7331));
    Span4Mux_h I__1559 (
            .O(N__7374),
            .I(N__7331));
    LocalMux I__1558 (
            .O(N__7369),
            .I(N__7331));
    InMux I__1557 (
            .O(N__7368),
            .I(N__7324));
    InMux I__1556 (
            .O(N__7367),
            .I(N__7324));
    InMux I__1555 (
            .O(N__7366),
            .I(N__7324));
    Odrv4 I__1554 (
            .O(N__7363),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1553 (
            .O(N__7360),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1552 (
            .O(N__7355),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1551 (
            .O(N__7352),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1550 (
            .O(N__7349),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1549 (
            .O(N__7342),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1548 (
            .O(N__7331),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1547 (
            .O(N__7324),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    InMux I__1546 (
            .O(N__7307),
            .I(N__7303));
    InMux I__1545 (
            .O(N__7306),
            .I(N__7300));
    LocalMux I__1544 (
            .O(N__7303),
            .I(N__7291));
    LocalMux I__1543 (
            .O(N__7300),
            .I(N__7291));
    InMux I__1542 (
            .O(N__7299),
            .I(N__7286));
    InMux I__1541 (
            .O(N__7298),
            .I(N__7286));
    InMux I__1540 (
            .O(N__7297),
            .I(N__7281));
    InMux I__1539 (
            .O(N__7296),
            .I(N__7281));
    Odrv4 I__1538 (
            .O(N__7291),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1 ));
    LocalMux I__1537 (
            .O(N__7286),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1 ));
    LocalMux I__1536 (
            .O(N__7281),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1 ));
    InMux I__1535 (
            .O(N__7274),
            .I(N__7271));
    LocalMux I__1534 (
            .O(N__7271),
            .I(N__7268));
    Odrv4 I__1533 (
            .O(N__7268),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__1532 (
            .O(N__7265),
            .I(N__7262));
    LocalMux I__1531 (
            .O(N__7262),
            .I(N__7259));
    Span4Mux_h I__1530 (
            .O(N__7259),
            .I(N__7256));
    Odrv4 I__1529 (
            .O(N__7256),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    IoInMux I__1528 (
            .O(N__7253),
            .I(N__7249));
    InMux I__1527 (
            .O(N__7252),
            .I(N__7246));
    LocalMux I__1526 (
            .O(N__7249),
            .I(N__7243));
    LocalMux I__1525 (
            .O(N__7246),
            .I(N__7240));
    IoSpan4Mux I__1524 (
            .O(N__7243),
            .I(N__7237));
    Span12Mux_v I__1523 (
            .O(N__7240),
            .I(N__7234));
    IoSpan4Mux I__1522 (
            .O(N__7237),
            .I(N__7231));
    Span12Mux_h I__1521 (
            .O(N__7234),
            .I(N__7228));
    IoSpan4Mux I__1520 (
            .O(N__7231),
            .I(N__7225));
    Odrv12 I__1519 (
            .O(N__7228),
            .I(C3_c));
    Odrv4 I__1518 (
            .O(N__7225),
            .I(C3_c));
    InMux I__1517 (
            .O(N__7220),
            .I(N__7211));
    InMux I__1516 (
            .O(N__7219),
            .I(N__7211));
    InMux I__1515 (
            .O(N__7218),
            .I(N__7211));
    LocalMux I__1514 (
            .O(N__7211),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    IoInMux I__1513 (
            .O(N__7208),
            .I(N__7204));
    InMux I__1512 (
            .O(N__7207),
            .I(N__7201));
    LocalMux I__1511 (
            .O(N__7204),
            .I(N__7198));
    LocalMux I__1510 (
            .O(N__7201),
            .I(N__7195));
    Span4Mux_s3_h I__1509 (
            .O(N__7198),
            .I(N__7192));
    Span12Mux_v I__1508 (
            .O(N__7195),
            .I(N__7189));
    Sp12to4 I__1507 (
            .O(N__7192),
            .I(N__7186));
    Span12Mux_h I__1506 (
            .O(N__7189),
            .I(N__7183));
    Span12Mux_v I__1505 (
            .O(N__7186),
            .I(N__7180));
    Odrv12 I__1504 (
            .O(N__7183),
            .I(C1_c));
    Odrv12 I__1503 (
            .O(N__7180),
            .I(C1_c));
    CascadeMux I__1502 (
            .O(N__7175),
            .I(N__7170));
    CascadeMux I__1501 (
            .O(N__7174),
            .I(N__7167));
    InMux I__1500 (
            .O(N__7173),
            .I(N__7163));
    InMux I__1499 (
            .O(N__7170),
            .I(N__7160));
    InMux I__1498 (
            .O(N__7167),
            .I(N__7155));
    InMux I__1497 (
            .O(N__7166),
            .I(N__7155));
    LocalMux I__1496 (
            .O(N__7163),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__1495 (
            .O(N__7160),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__1494 (
            .O(N__7155),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__1493 (
            .O(N__7148),
            .I(N__7142));
    InMux I__1492 (
            .O(N__7147),
            .I(N__7142));
    LocalMux I__1491 (
            .O(N__7142),
            .I(N__7135));
    InMux I__1490 (
            .O(N__7141),
            .I(N__7132));
    InMux I__1489 (
            .O(N__7140),
            .I(N__7129));
    InMux I__1488 (
            .O(N__7139),
            .I(N__7124));
    InMux I__1487 (
            .O(N__7138),
            .I(N__7124));
    Sp12to4 I__1486 (
            .O(N__7135),
            .I(N__7121));
    LocalMux I__1485 (
            .O(N__7132),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1484 (
            .O(N__7129),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1483 (
            .O(N__7124),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv12 I__1482 (
            .O(N__7121),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__1481 (
            .O(N__7112),
            .I(N__7101));
    InMux I__1480 (
            .O(N__7111),
            .I(N__7101));
    InMux I__1479 (
            .O(N__7110),
            .I(N__7101));
    InMux I__1478 (
            .O(N__7109),
            .I(N__7096));
    InMux I__1477 (
            .O(N__7108),
            .I(N__7096));
    LocalMux I__1476 (
            .O(N__7101),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__1475 (
            .O(N__7096),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    InMux I__1474 (
            .O(N__7091),
            .I(N__7085));
    InMux I__1473 (
            .O(N__7090),
            .I(N__7078));
    InMux I__1472 (
            .O(N__7089),
            .I(N__7078));
    InMux I__1471 (
            .O(N__7088),
            .I(N__7078));
    LocalMux I__1470 (
            .O(N__7085),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__1469 (
            .O(N__7078),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    CascadeMux I__1468 (
            .O(N__7073),
            .I(N__7067));
    InMux I__1467 (
            .O(N__7072),
            .I(N__7064));
    InMux I__1466 (
            .O(N__7071),
            .I(N__7057));
    InMux I__1465 (
            .O(N__7070),
            .I(N__7057));
    InMux I__1464 (
            .O(N__7067),
            .I(N__7057));
    LocalMux I__1463 (
            .O(N__7064),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1462 (
            .O(N__7057),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    InMux I__1461 (
            .O(N__7052),
            .I(N__7048));
    InMux I__1460 (
            .O(N__7051),
            .I(N__7045));
    LocalMux I__1459 (
            .O(N__7048),
            .I(N__7042));
    LocalMux I__1458 (
            .O(N__7045),
            .I(N__7039));
    Odrv4 I__1457 (
            .O(N__7042),
            .I(\U712_REG_SM.N_210 ));
    Odrv4 I__1456 (
            .O(N__7039),
            .I(\U712_REG_SM.N_210 ));
    InMux I__1455 (
            .O(N__7034),
            .I(N__7025));
    InMux I__1454 (
            .O(N__7033),
            .I(N__7025));
    InMux I__1453 (
            .O(N__7032),
            .I(N__7025));
    LocalMux I__1452 (
            .O(N__7025),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    CascadeMux I__1451 (
            .O(N__7022),
            .I(N__7018));
    InMux I__1450 (
            .O(N__7021),
            .I(N__7015));
    InMux I__1449 (
            .O(N__7018),
            .I(N__7012));
    LocalMux I__1448 (
            .O(N__7015),
            .I(N__7005));
    LocalMux I__1447 (
            .O(N__7012),
            .I(N__7005));
    InMux I__1446 (
            .O(N__7011),
            .I(N__7000));
    InMux I__1445 (
            .O(N__7010),
            .I(N__7000));
    Span4Mux_v I__1444 (
            .O(N__7005),
            .I(N__6997));
    LocalMux I__1443 (
            .O(N__7000),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    Odrv4 I__1442 (
            .O(N__6997),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    CascadeMux I__1441 (
            .O(N__6992),
            .I(N__6989));
    InMux I__1440 (
            .O(N__6989),
            .I(N__6980));
    InMux I__1439 (
            .O(N__6988),
            .I(N__6980));
    InMux I__1438 (
            .O(N__6987),
            .I(N__6980));
    LocalMux I__1437 (
            .O(N__6980),
            .I(\U712_REG_SM.N_174 ));
    CascadeMux I__1436 (
            .O(N__6977),
            .I(N__6974));
    InMux I__1435 (
            .O(N__6974),
            .I(N__6970));
    InMux I__1434 (
            .O(N__6973),
            .I(N__6967));
    LocalMux I__1433 (
            .O(N__6970),
            .I(REG_TACK));
    LocalMux I__1432 (
            .O(N__6967),
            .I(REG_TACK));
    InMux I__1431 (
            .O(N__6962),
            .I(N__6958));
    InMux I__1430 (
            .O(N__6961),
            .I(N__6955));
    LocalMux I__1429 (
            .O(N__6958),
            .I(DBR_SYNCZ0Z_0));
    LocalMux I__1428 (
            .O(N__6955),
            .I(DBR_SYNCZ0Z_0));
    IoInMux I__1427 (
            .O(N__6950),
            .I(N__6947));
    LocalMux I__1426 (
            .O(N__6947),
            .I(N__6944));
    Span12Mux_s1_v I__1425 (
            .O(N__6944),
            .I(N__6941));
    Span12Mux_h I__1424 (
            .O(N__6941),
            .I(N__6938));
    Odrv12 I__1423 (
            .O(N__6938),
            .I(CASn_c));
    IoInMux I__1422 (
            .O(N__6935),
            .I(N__6932));
    LocalMux I__1421 (
            .O(N__6932),
            .I(N__6929));
    Span4Mux_s3_v I__1420 (
            .O(N__6929),
            .I(N__6926));
    Span4Mux_v I__1419 (
            .O(N__6926),
            .I(N__6923));
    Span4Mux_h I__1418 (
            .O(N__6923),
            .I(N__6920));
    Span4Mux_h I__1417 (
            .O(N__6920),
            .I(N__6917));
    Odrv4 I__1416 (
            .O(N__6917),
            .I(CMA_c_10));
    InMux I__1415 (
            .O(N__6914),
            .I(N__6911));
    LocalMux I__1414 (
            .O(N__6911),
            .I(N__6908));
    Odrv12 I__1413 (
            .O(N__6908),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    CascadeMux I__1412 (
            .O(N__6905),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_ ));
    IoInMux I__1411 (
            .O(N__6902),
            .I(N__6899));
    LocalMux I__1410 (
            .O(N__6899),
            .I(N__6896));
    IoSpan4Mux I__1409 (
            .O(N__6896),
            .I(N__6893));
    Span4Mux_s3_v I__1408 (
            .O(N__6893),
            .I(N__6890));
    Span4Mux_v I__1407 (
            .O(N__6890),
            .I(N__6887));
    Odrv4 I__1406 (
            .O(N__6887),
            .I(CMA_c_2));
    CascadeMux I__1405 (
            .O(N__6884),
            .I(N__6878));
    CascadeMux I__1404 (
            .O(N__6883),
            .I(N__6873));
    CascadeMux I__1403 (
            .O(N__6882),
            .I(N__6868));
    InMux I__1402 (
            .O(N__6881),
            .I(N__6863));
    InMux I__1401 (
            .O(N__6878),
            .I(N__6863));
    CascadeMux I__1400 (
            .O(N__6877),
            .I(N__6860));
    InMux I__1399 (
            .O(N__6876),
            .I(N__6856));
    InMux I__1398 (
            .O(N__6873),
            .I(N__6851));
    InMux I__1397 (
            .O(N__6872),
            .I(N__6851));
    InMux I__1396 (
            .O(N__6871),
            .I(N__6848));
    InMux I__1395 (
            .O(N__6868),
            .I(N__6845));
    LocalMux I__1394 (
            .O(N__6863),
            .I(N__6842));
    InMux I__1393 (
            .O(N__6860),
            .I(N__6837));
    InMux I__1392 (
            .O(N__6859),
            .I(N__6837));
    LocalMux I__1391 (
            .O(N__6856),
            .I(N__6834));
    LocalMux I__1390 (
            .O(N__6851),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1389 (
            .O(N__6848),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1388 (
            .O(N__6845),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__1387 (
            .O(N__6842),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1386 (
            .O(N__6837),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__1385 (
            .O(N__6834),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    InMux I__1384 (
            .O(N__6821),
            .I(N__6818));
    LocalMux I__1383 (
            .O(N__6818),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__1382 (
            .O(N__6815),
            .I(N__6812));
    LocalMux I__1381 (
            .O(N__6812),
            .I(N__6809));
    IoSpan4Mux I__1380 (
            .O(N__6809),
            .I(N__6806));
    IoSpan4Mux I__1379 (
            .O(N__6806),
            .I(N__6803));
    Span4Mux_s2_h I__1378 (
            .O(N__6803),
            .I(N__6800));
    Sp12to4 I__1377 (
            .O(N__6800),
            .I(N__6797));
    Span12Mux_h I__1376 (
            .O(N__6797),
            .I(N__6794));
    Odrv12 I__1375 (
            .O(N__6794),
            .I(CMA_c_3));
    CascadeMux I__1374 (
            .O(N__6791),
            .I(\U712_REG_SM.N_199_cascade_ ));
    CascadeMux I__1373 (
            .O(N__6788),
            .I(N__6784));
    InMux I__1372 (
            .O(N__6787),
            .I(N__6781));
    InMux I__1371 (
            .O(N__6784),
            .I(N__6778));
    LocalMux I__1370 (
            .O(N__6781),
            .I(N__6775));
    LocalMux I__1369 (
            .O(N__6778),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    Odrv12 I__1368 (
            .O(N__6775),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__1367 (
            .O(N__6770),
            .I(N__6767));
    InMux I__1366 (
            .O(N__6767),
            .I(N__6762));
    InMux I__1365 (
            .O(N__6766),
            .I(N__6759));
    InMux I__1364 (
            .O(N__6765),
            .I(N__6756));
    LocalMux I__1363 (
            .O(N__6762),
            .I(N__6753));
    LocalMux I__1362 (
            .O(N__6759),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__1361 (
            .O(N__6756),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    Odrv12 I__1360 (
            .O(N__6753),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__1359 (
            .O(N__6746),
            .I(\U712_CYCLE_TERM.N_208_i_0_en_cascade_ ));
    CEMux I__1358 (
            .O(N__6743),
            .I(N__6740));
    LocalMux I__1357 (
            .O(N__6740),
            .I(N__6737));
    Odrv12 I__1356 (
            .O(N__6737),
            .I(\U712_CYCLE_TERM.N_208_i_0_en_0 ));
    InMux I__1355 (
            .O(N__6734),
            .I(N__6731));
    LocalMux I__1354 (
            .O(N__6731),
            .I(\U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a3_0_2 ));
    CascadeMux I__1353 (
            .O(N__6728),
            .I(N__6724));
    InMux I__1352 (
            .O(N__6727),
            .I(N__6721));
    InMux I__1351 (
            .O(N__6724),
            .I(N__6715));
    LocalMux I__1350 (
            .O(N__6721),
            .I(N__6711));
    InMux I__1349 (
            .O(N__6720),
            .I(N__6708));
    InMux I__1348 (
            .O(N__6719),
            .I(N__6702));
    InMux I__1347 (
            .O(N__6718),
            .I(N__6702));
    LocalMux I__1346 (
            .O(N__6715),
            .I(N__6698));
    InMux I__1345 (
            .O(N__6714),
            .I(N__6688));
    Span4Mux_v I__1344 (
            .O(N__6711),
            .I(N__6685));
    LocalMux I__1343 (
            .O(N__6708),
            .I(N__6682));
    InMux I__1342 (
            .O(N__6707),
            .I(N__6679));
    LocalMux I__1341 (
            .O(N__6702),
            .I(N__6676));
    InMux I__1340 (
            .O(N__6701),
            .I(N__6673));
    Span4Mux_v I__1339 (
            .O(N__6698),
            .I(N__6670));
    InMux I__1338 (
            .O(N__6697),
            .I(N__6667));
    InMux I__1337 (
            .O(N__6696),
            .I(N__6662));
    InMux I__1336 (
            .O(N__6695),
            .I(N__6662));
    InMux I__1335 (
            .O(N__6694),
            .I(N__6657));
    InMux I__1334 (
            .O(N__6693),
            .I(N__6657));
    InMux I__1333 (
            .O(N__6692),
            .I(N__6652));
    InMux I__1332 (
            .O(N__6691),
            .I(N__6652));
    LocalMux I__1331 (
            .O(N__6688),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1330 (
            .O(N__6685),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1329 (
            .O(N__6682),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1328 (
            .O(N__6679),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1327 (
            .O(N__6676),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1326 (
            .O(N__6673),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1325 (
            .O(N__6670),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1324 (
            .O(N__6667),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1323 (
            .O(N__6662),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1322 (
            .O(N__6657),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1321 (
            .O(N__6652),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1320 (
            .O(N__6629),
            .I(N__6624));
    CascadeMux I__1319 (
            .O(N__6628),
            .I(N__6620));
    CascadeMux I__1318 (
            .O(N__6627),
            .I(N__6617));
    LocalMux I__1317 (
            .O(N__6624),
            .I(N__6607));
    InMux I__1316 (
            .O(N__6623),
            .I(N__6604));
    InMux I__1315 (
            .O(N__6620),
            .I(N__6599));
    InMux I__1314 (
            .O(N__6617),
            .I(N__6599));
    InMux I__1313 (
            .O(N__6616),
            .I(N__6596));
    InMux I__1312 (
            .O(N__6615),
            .I(N__6593));
    InMux I__1311 (
            .O(N__6614),
            .I(N__6588));
    InMux I__1310 (
            .O(N__6613),
            .I(N__6588));
    InMux I__1309 (
            .O(N__6612),
            .I(N__6585));
    InMux I__1308 (
            .O(N__6611),
            .I(N__6580));
    InMux I__1307 (
            .O(N__6610),
            .I(N__6580));
    Odrv4 I__1306 (
            .O(N__6607),
            .I(\U712_CHIP_RAM.N_165 ));
    LocalMux I__1305 (
            .O(N__6604),
            .I(\U712_CHIP_RAM.N_165 ));
    LocalMux I__1304 (
            .O(N__6599),
            .I(\U712_CHIP_RAM.N_165 ));
    LocalMux I__1303 (
            .O(N__6596),
            .I(\U712_CHIP_RAM.N_165 ));
    LocalMux I__1302 (
            .O(N__6593),
            .I(\U712_CHIP_RAM.N_165 ));
    LocalMux I__1301 (
            .O(N__6588),
            .I(\U712_CHIP_RAM.N_165 ));
    LocalMux I__1300 (
            .O(N__6585),
            .I(\U712_CHIP_RAM.N_165 ));
    LocalMux I__1299 (
            .O(N__6580),
            .I(\U712_CHIP_RAM.N_165 ));
    InMux I__1298 (
            .O(N__6563),
            .I(N__6560));
    LocalMux I__1297 (
            .O(N__6560),
            .I(\U712_CHIP_RAM.N_249 ));
    InMux I__1296 (
            .O(N__6557),
            .I(N__6553));
    InMux I__1295 (
            .O(N__6556),
            .I(N__6550));
    LocalMux I__1294 (
            .O(N__6553),
            .I(N__6547));
    LocalMux I__1293 (
            .O(N__6550),
            .I(CPU_TACKm));
    Odrv4 I__1292 (
            .O(N__6547),
            .I(CPU_TACKm));
    CascadeMux I__1291 (
            .O(N__6542),
            .I(N__6537));
    InMux I__1290 (
            .O(N__6541),
            .I(N__6534));
    InMux I__1289 (
            .O(N__6540),
            .I(N__6529));
    InMux I__1288 (
            .O(N__6537),
            .I(N__6529));
    LocalMux I__1287 (
            .O(N__6534),
            .I(N__6523));
    LocalMux I__1286 (
            .O(N__6529),
            .I(N__6523));
    InMux I__1285 (
            .O(N__6528),
            .I(N__6520));
    Odrv12 I__1284 (
            .O(N__6523),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__1283 (
            .O(N__6520),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CascadeMux I__1282 (
            .O(N__6515),
            .I(N__6512));
    InMux I__1281 (
            .O(N__6512),
            .I(N__6509));
    LocalMux I__1280 (
            .O(N__6509),
            .I(N__6506));
    Odrv4 I__1279 (
            .O(N__6506),
            .I(\U712_REG_SM.N_199 ));
    InMux I__1278 (
            .O(N__6503),
            .I(N__6500));
    LocalMux I__1277 (
            .O(N__6500),
            .I(\U712_REG_SM.N_171 ));
    CascadeMux I__1276 (
            .O(N__6497),
            .I(\U712_REG_SM.N_174_cascade_ ));
    InMux I__1275 (
            .O(N__6494),
            .I(N__6490));
    InMux I__1274 (
            .O(N__6493),
            .I(N__6487));
    LocalMux I__1273 (
            .O(N__6490),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1272 (
            .O(N__6487),
            .I(DBR_SYNCZ0Z_1));
    InMux I__1271 (
            .O(N__6482),
            .I(N__6478));
    InMux I__1270 (
            .O(N__6481),
            .I(N__6475));
    LocalMux I__1269 (
            .O(N__6478),
            .I(N__6472));
    LocalMux I__1268 (
            .O(N__6475),
            .I(N__6469));
    Sp12to4 I__1267 (
            .O(N__6472),
            .I(N__6466));
    Span4Mux_v I__1266 (
            .O(N__6469),
            .I(N__6463));
    Span12Mux_h I__1265 (
            .O(N__6466),
            .I(N__6460));
    Sp12to4 I__1264 (
            .O(N__6463),
            .I(N__6457));
    Span12Mux_v I__1263 (
            .O(N__6460),
            .I(N__6452));
    Span12Mux_h I__1262 (
            .O(N__6457),
            .I(N__6452));
    Odrv12 I__1261 (
            .O(N__6452),
            .I(RnW_c));
    InMux I__1260 (
            .O(N__6449),
            .I(N__6446));
    LocalMux I__1259 (
            .O(N__6446),
            .I(N__6441));
    InMux I__1258 (
            .O(N__6445),
            .I(N__6438));
    InMux I__1257 (
            .O(N__6444),
            .I(N__6435));
    Span4Mux_h I__1256 (
            .O(N__6441),
            .I(N__6430));
    LocalMux I__1255 (
            .O(N__6438),
            .I(N__6430));
    LocalMux I__1254 (
            .O(N__6435),
            .I(N__6427));
    Span4Mux_h I__1253 (
            .O(N__6430),
            .I(N__6424));
    Span4Mux_v I__1252 (
            .O(N__6427),
            .I(N__6421));
    Sp12to4 I__1251 (
            .O(N__6424),
            .I(N__6418));
    IoSpan4Mux I__1250 (
            .O(N__6421),
            .I(N__6415));
    Span12Mux_v I__1249 (
            .O(N__6418),
            .I(N__6412));
    IoSpan4Mux I__1248 (
            .O(N__6415),
            .I(N__6409));
    Odrv12 I__1247 (
            .O(N__6412),
            .I(AWEn_c));
    Odrv4 I__1246 (
            .O(N__6409),
            .I(AWEn_c));
    InMux I__1245 (
            .O(N__6404),
            .I(N__6398));
    InMux I__1244 (
            .O(N__6403),
            .I(N__6391));
    InMux I__1243 (
            .O(N__6402),
            .I(N__6391));
    InMux I__1242 (
            .O(N__6401),
            .I(N__6388));
    LocalMux I__1241 (
            .O(N__6398),
            .I(N__6385));
    InMux I__1240 (
            .O(N__6397),
            .I(N__6382));
    CascadeMux I__1239 (
            .O(N__6396),
            .I(N__6377));
    LocalMux I__1238 (
            .O(N__6391),
            .I(N__6372));
    LocalMux I__1237 (
            .O(N__6388),
            .I(N__6369));
    Span4Mux_h I__1236 (
            .O(N__6385),
            .I(N__6366));
    LocalMux I__1235 (
            .O(N__6382),
            .I(N__6363));
    InMux I__1234 (
            .O(N__6381),
            .I(N__6358));
    InMux I__1233 (
            .O(N__6380),
            .I(N__6358));
    InMux I__1232 (
            .O(N__6377),
            .I(N__6353));
    InMux I__1231 (
            .O(N__6376),
            .I(N__6353));
    InMux I__1230 (
            .O(N__6375),
            .I(N__6350));
    Span4Mux_h I__1229 (
            .O(N__6372),
            .I(N__6347));
    Odrv4 I__1228 (
            .O(N__6369),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1227 (
            .O(N__6366),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1226 (
            .O(N__6363),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1225 (
            .O(N__6358),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1224 (
            .O(N__6353),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1223 (
            .O(N__6350),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1222 (
            .O(N__6347),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1221 (
            .O(N__6332),
            .I(N__6329));
    LocalMux I__1220 (
            .O(N__6329),
            .I(N__6326));
    Odrv4 I__1219 (
            .O(N__6326),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_RNOZ0Z_0 ));
    CascadeMux I__1218 (
            .O(N__6323),
            .I(N__6317));
    CascadeMux I__1217 (
            .O(N__6322),
            .I(N__6313));
    InMux I__1216 (
            .O(N__6321),
            .I(N__6309));
    InMux I__1215 (
            .O(N__6320),
            .I(N__6306));
    InMux I__1214 (
            .O(N__6317),
            .I(N__6302));
    InMux I__1213 (
            .O(N__6316),
            .I(N__6299));
    InMux I__1212 (
            .O(N__6313),
            .I(N__6290));
    InMux I__1211 (
            .O(N__6312),
            .I(N__6290));
    LocalMux I__1210 (
            .O(N__6309),
            .I(N__6285));
    LocalMux I__1209 (
            .O(N__6306),
            .I(N__6285));
    InMux I__1208 (
            .O(N__6305),
            .I(N__6282));
    LocalMux I__1207 (
            .O(N__6302),
            .I(N__6277));
    LocalMux I__1206 (
            .O(N__6299),
            .I(N__6277));
    CascadeMux I__1205 (
            .O(N__6298),
            .I(N__6274));
    CascadeMux I__1204 (
            .O(N__6297),
            .I(N__6270));
    InMux I__1203 (
            .O(N__6296),
            .I(N__6262));
    InMux I__1202 (
            .O(N__6295),
            .I(N__6259));
    LocalMux I__1201 (
            .O(N__6290),
            .I(N__6256));
    Span4Mux_h I__1200 (
            .O(N__6285),
            .I(N__6251));
    LocalMux I__1199 (
            .O(N__6282),
            .I(N__6251));
    Span4Mux_v I__1198 (
            .O(N__6277),
            .I(N__6248));
    InMux I__1197 (
            .O(N__6274),
            .I(N__6245));
    InMux I__1196 (
            .O(N__6273),
            .I(N__6242));
    InMux I__1195 (
            .O(N__6270),
            .I(N__6239));
    InMux I__1194 (
            .O(N__6269),
            .I(N__6234));
    InMux I__1193 (
            .O(N__6268),
            .I(N__6234));
    InMux I__1192 (
            .O(N__6267),
            .I(N__6227));
    InMux I__1191 (
            .O(N__6266),
            .I(N__6227));
    InMux I__1190 (
            .O(N__6265),
            .I(N__6227));
    LocalMux I__1189 (
            .O(N__6262),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1188 (
            .O(N__6259),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1187 (
            .O(N__6256),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1186 (
            .O(N__6251),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1185 (
            .O(N__6248),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1184 (
            .O(N__6245),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1183 (
            .O(N__6242),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1182 (
            .O(N__6239),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1181 (
            .O(N__6234),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1180 (
            .O(N__6227),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1179 (
            .O(N__6206),
            .I(N__6203));
    LocalMux I__1178 (
            .O(N__6203),
            .I(N__6199));
    InMux I__1177 (
            .O(N__6202),
            .I(N__6196));
    Odrv4 I__1176 (
            .O(N__6199),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1 ));
    LocalMux I__1175 (
            .O(N__6196),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1 ));
    CascadeMux I__1174 (
            .O(N__6191),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1_cascade_ ));
    InMux I__1173 (
            .O(N__6188),
            .I(N__6182));
    CascadeMux I__1172 (
            .O(N__6187),
            .I(N__6178));
    InMux I__1171 (
            .O(N__6186),
            .I(N__6172));
    InMux I__1170 (
            .O(N__6185),
            .I(N__6168));
    LocalMux I__1169 (
            .O(N__6182),
            .I(N__6165));
    InMux I__1168 (
            .O(N__6181),
            .I(N__6162));
    InMux I__1167 (
            .O(N__6178),
            .I(N__6158));
    InMux I__1166 (
            .O(N__6177),
            .I(N__6152));
    InMux I__1165 (
            .O(N__6176),
            .I(N__6152));
    InMux I__1164 (
            .O(N__6175),
            .I(N__6148));
    LocalMux I__1163 (
            .O(N__6172),
            .I(N__6145));
    InMux I__1162 (
            .O(N__6171),
            .I(N__6142));
    LocalMux I__1161 (
            .O(N__6168),
            .I(N__6137));
    Span4Mux_v I__1160 (
            .O(N__6165),
            .I(N__6137));
    LocalMux I__1159 (
            .O(N__6162),
            .I(N__6134));
    InMux I__1158 (
            .O(N__6161),
            .I(N__6131));
    LocalMux I__1157 (
            .O(N__6158),
            .I(N__6128));
    InMux I__1156 (
            .O(N__6157),
            .I(N__6125));
    LocalMux I__1155 (
            .O(N__6152),
            .I(N__6122));
    InMux I__1154 (
            .O(N__6151),
            .I(N__6119));
    LocalMux I__1153 (
            .O(N__6148),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1152 (
            .O(N__6145),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1151 (
            .O(N__6142),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1150 (
            .O(N__6137),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1149 (
            .O(N__6134),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1148 (
            .O(N__6131),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv12 I__1147 (
            .O(N__6128),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1146 (
            .O(N__6125),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1145 (
            .O(N__6122),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1144 (
            .O(N__6119),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__1143 (
            .O(N__6098),
            .I(N__6095));
    LocalMux I__1142 (
            .O(N__6095),
            .I(N__6092));
    Odrv4 I__1141 (
            .O(N__6092),
            .I(\U712_CHIP_RAM.N_248 ));
    CascadeMux I__1140 (
            .O(N__6089),
            .I(N__6085));
    CascadeMux I__1139 (
            .O(N__6088),
            .I(N__6081));
    InMux I__1138 (
            .O(N__6085),
            .I(N__6074));
    InMux I__1137 (
            .O(N__6084),
            .I(N__6071));
    InMux I__1136 (
            .O(N__6081),
            .I(N__6068));
    InMux I__1135 (
            .O(N__6080),
            .I(N__6065));
    InMux I__1134 (
            .O(N__6079),
            .I(N__6062));
    InMux I__1133 (
            .O(N__6078),
            .I(N__6057));
    InMux I__1132 (
            .O(N__6077),
            .I(N__6050));
    LocalMux I__1131 (
            .O(N__6074),
            .I(N__6045));
    LocalMux I__1130 (
            .O(N__6071),
            .I(N__6045));
    LocalMux I__1129 (
            .O(N__6068),
            .I(N__6038));
    LocalMux I__1128 (
            .O(N__6065),
            .I(N__6033));
    LocalMux I__1127 (
            .O(N__6062),
            .I(N__6033));
    InMux I__1126 (
            .O(N__6061),
            .I(N__6030));
    InMux I__1125 (
            .O(N__6060),
            .I(N__6027));
    LocalMux I__1124 (
            .O(N__6057),
            .I(N__6024));
    InMux I__1123 (
            .O(N__6056),
            .I(N__6021));
    InMux I__1122 (
            .O(N__6055),
            .I(N__6016));
    InMux I__1121 (
            .O(N__6054),
            .I(N__6016));
    InMux I__1120 (
            .O(N__6053),
            .I(N__6013));
    LocalMux I__1119 (
            .O(N__6050),
            .I(N__6008));
    Span4Mux_v I__1118 (
            .O(N__6045),
            .I(N__6008));
    InMux I__1117 (
            .O(N__6044),
            .I(N__6003));
    InMux I__1116 (
            .O(N__6043),
            .I(N__6003));
    InMux I__1115 (
            .O(N__6042),
            .I(N__5998));
    InMux I__1114 (
            .O(N__6041),
            .I(N__5998));
    Span4Mux_v I__1113 (
            .O(N__6038),
            .I(N__5993));
    Span4Mux_v I__1112 (
            .O(N__6033),
            .I(N__5993));
    LocalMux I__1111 (
            .O(N__6030),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1110 (
            .O(N__6027),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1109 (
            .O(N__6024),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1108 (
            .O(N__6021),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1107 (
            .O(N__6016),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1106 (
            .O(N__6013),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1105 (
            .O(N__6008),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1104 (
            .O(N__6003),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1103 (
            .O(N__5998),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1102 (
            .O(N__5993),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1101 (
            .O(N__5972),
            .I(N__5968));
    InMux I__1100 (
            .O(N__5971),
            .I(N__5965));
    LocalMux I__1099 (
            .O(N__5968),
            .I(N__5958));
    LocalMux I__1098 (
            .O(N__5965),
            .I(N__5958));
    InMux I__1097 (
            .O(N__5964),
            .I(N__5955));
    InMux I__1096 (
            .O(N__5963),
            .I(N__5952));
    Span4Mux_h I__1095 (
            .O(N__5958),
            .I(N__5949));
    LocalMux I__1094 (
            .O(N__5955),
            .I(N__5946));
    LocalMux I__1093 (
            .O(N__5952),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2Z0Z_1 ));
    Odrv4 I__1092 (
            .O(N__5949),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2Z0Z_1 ));
    Odrv4 I__1091 (
            .O(N__5946),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2Z0Z_1 ));
    CascadeMux I__1090 (
            .O(N__5939),
            .I(\U712_REG_SM.N_171_cascade_ ));
    CascadeMux I__1089 (
            .O(N__5936),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa_0_a2_0_a3_1_cascade_ ));
    CascadeMux I__1088 (
            .O(N__5933),
            .I(N__5929));
    InMux I__1087 (
            .O(N__5932),
            .I(N__5926));
    InMux I__1086 (
            .O(N__5929),
            .I(N__5923));
    LocalMux I__1085 (
            .O(N__5926),
            .I(N__5920));
    LocalMux I__1084 (
            .O(N__5923),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    Odrv4 I__1083 (
            .O(N__5920),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    CascadeMux I__1082 (
            .O(N__5915),
            .I(N__5912));
    InMux I__1081 (
            .O(N__5912),
            .I(N__5906));
    InMux I__1080 (
            .O(N__5911),
            .I(N__5906));
    LocalMux I__1079 (
            .O(N__5906),
            .I(N__5903));
    Span4Mux_v I__1078 (
            .O(N__5903),
            .I(N__5900));
    Span4Mux_v I__1077 (
            .O(N__5900),
            .I(N__5897));
    Sp12to4 I__1076 (
            .O(N__5897),
            .I(N__5894));
    Span12Mux_h I__1075 (
            .O(N__5894),
            .I(N__5891));
    Odrv12 I__1074 (
            .O(N__5891),
            .I(A_c_14));
    InMux I__1073 (
            .O(N__5888),
            .I(N__5885));
    LocalMux I__1072 (
            .O(N__5885),
            .I(N__5882));
    Span4Mux_v I__1071 (
            .O(N__5882),
            .I(N__5879));
    Sp12to4 I__1070 (
            .O(N__5879),
            .I(N__5876));
    Span12Mux_h I__1069 (
            .O(N__5876),
            .I(N__5873));
    Span12Mux_v I__1068 (
            .O(N__5873),
            .I(N__5870));
    Odrv12 I__1067 (
            .O(N__5870),
            .I(A_c_3));
    InMux I__1066 (
            .O(N__5867),
            .I(N__5864));
    LocalMux I__1065 (
            .O(N__5864),
            .I(N__5861));
    Span4Mux_v I__1064 (
            .O(N__5861),
            .I(N__5858));
    Sp12to4 I__1063 (
            .O(N__5858),
            .I(N__5855));
    Span12Mux_h I__1062 (
            .O(N__5855),
            .I(N__5852));
    Odrv12 I__1061 (
            .O(N__5852),
            .I(A_c_10));
    CascadeMux I__1060 (
            .O(N__5849),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ));
    InMux I__1059 (
            .O(N__5846),
            .I(N__5843));
    LocalMux I__1058 (
            .O(N__5843),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    CascadeMux I__1057 (
            .O(N__5840),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ));
    InMux I__1056 (
            .O(N__5837),
            .I(N__5834));
    LocalMux I__1055 (
            .O(N__5834),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    IoInMux I__1054 (
            .O(N__5831),
            .I(N__5828));
    LocalMux I__1053 (
            .O(N__5828),
            .I(N__5825));
    Span4Mux_s3_v I__1052 (
            .O(N__5825),
            .I(N__5822));
    Span4Mux_v I__1051 (
            .O(N__5822),
            .I(N__5819));
    Span4Mux_v I__1050 (
            .O(N__5819),
            .I(N__5816));
    Odrv4 I__1049 (
            .O(N__5816),
            .I(CMA_c_1));
    InMux I__1048 (
            .O(N__5813),
            .I(N__5810));
    LocalMux I__1047 (
            .O(N__5810),
            .I(N__5807));
    Odrv4 I__1046 (
            .O(N__5807),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__1045 (
            .O(N__5804),
            .I(N__5801));
    LocalMux I__1044 (
            .O(N__5801),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    IoInMux I__1043 (
            .O(N__5798),
            .I(N__5795));
    LocalMux I__1042 (
            .O(N__5795),
            .I(N__5792));
    Span4Mux_s1_h I__1041 (
            .O(N__5792),
            .I(N__5789));
    Span4Mux_h I__1040 (
            .O(N__5789),
            .I(N__5786));
    Sp12to4 I__1039 (
            .O(N__5786),
            .I(N__5783));
    Span12Mux_s8_v I__1038 (
            .O(N__5783),
            .I(N__5780));
    Span12Mux_h I__1037 (
            .O(N__5780),
            .I(N__5777));
    Odrv12 I__1036 (
            .O(N__5777),
            .I(CMA_c_5));
    InMux I__1035 (
            .O(N__5774),
            .I(N__5771));
    LocalMux I__1034 (
            .O(N__5771),
            .I(N__5768));
    Span4Mux_v I__1033 (
            .O(N__5768),
            .I(N__5765));
    Span4Mux_h I__1032 (
            .O(N__5765),
            .I(N__5762));
    Sp12to4 I__1031 (
            .O(N__5762),
            .I(N__5759));
    Odrv12 I__1030 (
            .O(N__5759),
            .I(A_c_7));
    CascadeMux I__1029 (
            .O(N__5756),
            .I(\U712_CHIP_RAM.N_324_cascade_ ));
    InMux I__1028 (
            .O(N__5753),
            .I(N__5750));
    LocalMux I__1027 (
            .O(N__5750),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    InMux I__1026 (
            .O(N__5747),
            .I(N__5744));
    LocalMux I__1025 (
            .O(N__5744),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__1024 (
            .O(N__5741),
            .I(N__5738));
    LocalMux I__1023 (
            .O(N__5738),
            .I(N__5735));
    IoSpan4Mux I__1022 (
            .O(N__5735),
            .I(N__5732));
    Span4Mux_s3_h I__1021 (
            .O(N__5732),
            .I(N__5729));
    Sp12to4 I__1020 (
            .O(N__5729),
            .I(N__5726));
    Span12Mux_h I__1019 (
            .O(N__5726),
            .I(N__5723));
    Odrv12 I__1018 (
            .O(N__5723),
            .I(CMA_c_7));
    InMux I__1017 (
            .O(N__5720),
            .I(N__5717));
    LocalMux I__1016 (
            .O(N__5717),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__1015 (
            .O(N__5714),
            .I(N__5711));
    LocalMux I__1014 (
            .O(N__5711),
            .I(N__5708));
    Span4Mux_s2_h I__1013 (
            .O(N__5708),
            .I(N__5705));
    Span4Mux_v I__1012 (
            .O(N__5705),
            .I(N__5702));
    Span4Mux_v I__1011 (
            .O(N__5702),
            .I(N__5699));
    Sp12to4 I__1010 (
            .O(N__5699),
            .I(N__5696));
    Span12Mux_s9_h I__1009 (
            .O(N__5696),
            .I(N__5693));
    Odrv12 I__1008 (
            .O(N__5693),
            .I(CMA_c_6));
    InMux I__1007 (
            .O(N__5690),
            .I(N__5687));
    LocalMux I__1006 (
            .O(N__5687),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    CascadeMux I__1005 (
            .O(N__5684),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_ ));
    IoInMux I__1004 (
            .O(N__5681),
            .I(N__5678));
    LocalMux I__1003 (
            .O(N__5678),
            .I(N__5675));
    IoSpan4Mux I__1002 (
            .O(N__5675),
            .I(N__5672));
    Span4Mux_s1_h I__1001 (
            .O(N__5672),
            .I(N__5669));
    Sp12to4 I__1000 (
            .O(N__5669),
            .I(N__5666));
    Span12Mux_s11_v I__999 (
            .O(N__5666),
            .I(N__5663));
    Span12Mux_h I__998 (
            .O(N__5663),
            .I(N__5660));
    Odrv12 I__997 (
            .O(N__5660),
            .I(CMA_c_4));
    CascadeMux I__996 (
            .O(N__5657),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ));
    InMux I__995 (
            .O(N__5654),
            .I(N__5651));
    LocalMux I__994 (
            .O(N__5651),
            .I(N__5648));
    Odrv4 I__993 (
            .O(N__5648),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    IoInMux I__992 (
            .O(N__5645),
            .I(N__5642));
    LocalMux I__991 (
            .O(N__5642),
            .I(N__5639));
    IoSpan4Mux I__990 (
            .O(N__5639),
            .I(N__5636));
    Span4Mux_s2_v I__989 (
            .O(N__5636),
            .I(N__5631));
    InMux I__988 (
            .O(N__5635),
            .I(N__5626));
    InMux I__987 (
            .O(N__5634),
            .I(N__5626));
    Sp12to4 I__986 (
            .O(N__5631),
            .I(N__5623));
    LocalMux I__985 (
            .O(N__5626),
            .I(N__5620));
    Span12Mux_v I__984 (
            .O(N__5623),
            .I(N__5616));
    Span4Mux_v I__983 (
            .O(N__5620),
            .I(N__5613));
    InMux I__982 (
            .O(N__5619),
            .I(N__5610));
    Odrv12 I__981 (
            .O(N__5616),
            .I(DBENn_c));
    Odrv4 I__980 (
            .O(N__5613),
            .I(DBENn_c));
    LocalMux I__979 (
            .O(N__5610),
            .I(DBENn_c));
    InMux I__978 (
            .O(N__5603),
            .I(N__5600));
    LocalMux I__977 (
            .O(N__5600),
            .I(\U712_BYTE_ENABLE.N_268 ));
    IoInMux I__976 (
            .O(N__5597),
            .I(N__5594));
    LocalMux I__975 (
            .O(N__5594),
            .I(N__5591));
    IoSpan4Mux I__974 (
            .O(N__5591),
            .I(N__5588));
    IoSpan4Mux I__973 (
            .O(N__5588),
            .I(N__5585));
    Sp12to4 I__972 (
            .O(N__5585),
            .I(N__5582));
    Span12Mux_s7_v I__971 (
            .O(N__5582),
            .I(N__5579));
    Span12Mux_h I__970 (
            .O(N__5579),
            .I(N__5576));
    Odrv12 I__969 (
            .O(N__5576),
            .I(N_185_i));
    CascadeMux I__968 (
            .O(N__5573),
            .I(\U712_BYTE_ENABLE.N_270_cascade_ ));
    IoInMux I__967 (
            .O(N__5570),
            .I(N__5567));
    LocalMux I__966 (
            .O(N__5567),
            .I(N__5564));
    IoSpan4Mux I__965 (
            .O(N__5564),
            .I(N__5561));
    Sp12to4 I__964 (
            .O(N__5561),
            .I(N__5558));
    Span12Mux_s7_v I__963 (
            .O(N__5558),
            .I(N__5555));
    Span12Mux_h I__962 (
            .O(N__5555),
            .I(N__5552));
    Span12Mux_v I__961 (
            .O(N__5552),
            .I(N__5549));
    Odrv12 I__960 (
            .O(N__5549),
            .I(N_186_i));
    InMux I__959 (
            .O(N__5546),
            .I(N__5543));
    LocalMux I__958 (
            .O(N__5543),
            .I(\U712_BYTE_ENABLE.N_272 ));
    CascadeMux I__957 (
            .O(N__5540),
            .I(N__5536));
    CascadeMux I__956 (
            .O(N__5539),
            .I(N__5533));
    InMux I__955 (
            .O(N__5536),
            .I(N__5530));
    InMux I__954 (
            .O(N__5533),
            .I(N__5527));
    LocalMux I__953 (
            .O(N__5530),
            .I(N__5523));
    LocalMux I__952 (
            .O(N__5527),
            .I(N__5520));
    InMux I__951 (
            .O(N__5526),
            .I(N__5517));
    Span4Mux_v I__950 (
            .O(N__5523),
            .I(N__5512));
    Span4Mux_v I__949 (
            .O(N__5520),
            .I(N__5512));
    LocalMux I__948 (
            .O(N__5517),
            .I(N__5509));
    Sp12to4 I__947 (
            .O(N__5512),
            .I(N__5506));
    Span12Mux_h I__946 (
            .O(N__5509),
            .I(N__5503));
    Span12Mux_h I__945 (
            .O(N__5506),
            .I(N__5500));
    Span12Mux_v I__944 (
            .O(N__5503),
            .I(N__5497));
    Span12Mux_v I__943 (
            .O(N__5500),
            .I(N__5494));
    Odrv12 I__942 (
            .O(N__5497),
            .I(CASLn_c));
    Odrv12 I__941 (
            .O(N__5494),
            .I(CASLn_c));
    InMux I__940 (
            .O(N__5489),
            .I(N__5483));
    InMux I__939 (
            .O(N__5488),
            .I(N__5483));
    LocalMux I__938 (
            .O(N__5483),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0 ));
    IoInMux I__937 (
            .O(N__5480),
            .I(N__5477));
    LocalMux I__936 (
            .O(N__5477),
            .I(N__5474));
    IoSpan4Mux I__935 (
            .O(N__5474),
            .I(N__5471));
    Sp12to4 I__934 (
            .O(N__5471),
            .I(N__5468));
    Span12Mux_s7_v I__933 (
            .O(N__5468),
            .I(N__5465));
    Span12Mux_v I__932 (
            .O(N__5465),
            .I(N__5462));
    Odrv12 I__931 (
            .O(N__5462),
            .I(N_187_i));
    InMux I__930 (
            .O(N__5459),
            .I(N__5453));
    InMux I__929 (
            .O(N__5458),
            .I(N__5453));
    LocalMux I__928 (
            .O(N__5453),
            .I(N__5448));
    InMux I__927 (
            .O(N__5452),
            .I(N__5443));
    InMux I__926 (
            .O(N__5451),
            .I(N__5443));
    Span4Mux_v I__925 (
            .O(N__5448),
            .I(N__5440));
    LocalMux I__924 (
            .O(N__5443),
            .I(N__5437));
    Span4Mux_v I__923 (
            .O(N__5440),
            .I(N__5434));
    Span4Mux_v I__922 (
            .O(N__5437),
            .I(N__5431));
    Span4Mux_h I__921 (
            .O(N__5434),
            .I(N__5428));
    Span4Mux_v I__920 (
            .O(N__5431),
            .I(N__5425));
    Sp12to4 I__919 (
            .O(N__5428),
            .I(N__5420));
    Sp12to4 I__918 (
            .O(N__5425),
            .I(N__5420));
    Odrv12 I__917 (
            .O(N__5420),
            .I(A_c_1));
    InMux I__916 (
            .O(N__5417),
            .I(N__5405));
    InMux I__915 (
            .O(N__5416),
            .I(N__5405));
    InMux I__914 (
            .O(N__5415),
            .I(N__5405));
    InMux I__913 (
            .O(N__5414),
            .I(N__5405));
    LocalMux I__912 (
            .O(N__5405),
            .I(\U712_BYTE_ENABLE.N_265 ));
    InMux I__911 (
            .O(N__5402),
            .I(N__5396));
    InMux I__910 (
            .O(N__5401),
            .I(N__5396));
    LocalMux I__909 (
            .O(N__5396),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0 ));
    CascadeMux I__908 (
            .O(N__5393),
            .I(\U712_BYTE_ENABLE.N_266_cascade_ ));
    InMux I__907 (
            .O(N__5390),
            .I(N__5385));
    InMux I__906 (
            .O(N__5389),
            .I(N__5380));
    InMux I__905 (
            .O(N__5388),
            .I(N__5380));
    LocalMux I__904 (
            .O(N__5385),
            .I(N__5375));
    LocalMux I__903 (
            .O(N__5380),
            .I(N__5375));
    Span12Mux_v I__902 (
            .O(N__5375),
            .I(N__5372));
    Span12Mux_h I__901 (
            .O(N__5372),
            .I(N__5369));
    Odrv12 I__900 (
            .O(N__5369),
            .I(CASUn_c));
    IoInMux I__899 (
            .O(N__5366),
            .I(N__5363));
    LocalMux I__898 (
            .O(N__5363),
            .I(N__5360));
    Span4Mux_s2_h I__897 (
            .O(N__5360),
            .I(N__5357));
    Span4Mux_h I__896 (
            .O(N__5357),
            .I(N__5354));
    Sp12to4 I__895 (
            .O(N__5354),
            .I(N__5351));
    Span12Mux_v I__894 (
            .O(N__5351),
            .I(N__5348));
    Span12Mux_h I__893 (
            .O(N__5348),
            .I(N__5345));
    Odrv12 I__892 (
            .O(N__5345),
            .I(N_184_i));
    InMux I__891 (
            .O(N__5342),
            .I(N__5339));
    LocalMux I__890 (
            .O(N__5339),
            .I(N__5336));
    Span4Mux_v I__889 (
            .O(N__5336),
            .I(N__5331));
    InMux I__888 (
            .O(N__5335),
            .I(N__5326));
    InMux I__887 (
            .O(N__5334),
            .I(N__5326));
    Span4Mux_v I__886 (
            .O(N__5331),
            .I(N__5320));
    LocalMux I__885 (
            .O(N__5326),
            .I(N__5320));
    InMux I__884 (
            .O(N__5325),
            .I(N__5317));
    Span4Mux_v I__883 (
            .O(N__5320),
            .I(N__5312));
    LocalMux I__882 (
            .O(N__5317),
            .I(N__5309));
    InMux I__881 (
            .O(N__5316),
            .I(N__5304));
    InMux I__880 (
            .O(N__5315),
            .I(N__5304));
    Odrv4 I__879 (
            .O(N__5312),
            .I(DMA_CYCLEm));
    Odrv12 I__878 (
            .O(N__5309),
            .I(DMA_CYCLEm));
    LocalMux I__877 (
            .O(N__5304),
            .I(DMA_CYCLEm));
    IoInMux I__876 (
            .O(N__5297),
            .I(N__5294));
    LocalMux I__875 (
            .O(N__5294),
            .I(N__5291));
    Span4Mux_s1_h I__874 (
            .O(N__5291),
            .I(N__5288));
    Sp12to4 I__873 (
            .O(N__5288),
            .I(N__5285));
    Span12Mux_s6_v I__872 (
            .O(N__5285),
            .I(N__5282));
    Span12Mux_h I__871 (
            .O(N__5282),
            .I(N__5279));
    Odrv12 I__870 (
            .O(N__5279),
            .I(DRDDIR_i_m2));
    InMux I__869 (
            .O(N__5276),
            .I(N__5273));
    LocalMux I__868 (
            .O(N__5273),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__867 (
            .O(N__5270),
            .I(N__5267));
    LocalMux I__866 (
            .O(N__5267),
            .I(N__5264));
    Span4Mux_s2_v I__865 (
            .O(N__5264),
            .I(N__5261));
    Span4Mux_v I__864 (
            .O(N__5261),
            .I(N__5258));
    Span4Mux_v I__863 (
            .O(N__5258),
            .I(N__5255));
    Span4Mux_h I__862 (
            .O(N__5255),
            .I(N__5252));
    Odrv4 I__861 (
            .O(N__5252),
            .I(CMA_c_0));
    CascadeMux I__860 (
            .O(N__5249),
            .I(\U712_CHIP_RAM.N_219_cascade_ ));
    InMux I__859 (
            .O(N__5246),
            .I(N__5243));
    LocalMux I__858 (
            .O(N__5243),
            .I(N__5236));
    InMux I__857 (
            .O(N__5242),
            .I(N__5233));
    InMux I__856 (
            .O(N__5241),
            .I(N__5230));
    InMux I__855 (
            .O(N__5240),
            .I(N__5227));
    InMux I__854 (
            .O(N__5239),
            .I(N__5224));
    Span4Mux_v I__853 (
            .O(N__5236),
            .I(N__5217));
    LocalMux I__852 (
            .O(N__5233),
            .I(N__5217));
    LocalMux I__851 (
            .O(N__5230),
            .I(N__5217));
    LocalMux I__850 (
            .O(N__5227),
            .I(N__5214));
    LocalMux I__849 (
            .O(N__5224),
            .I(\U712_CHIP_RAM.N_166 ));
    Odrv4 I__848 (
            .O(N__5217),
            .I(\U712_CHIP_RAM.N_166 ));
    Odrv4 I__847 (
            .O(N__5214),
            .I(\U712_CHIP_RAM.N_166 ));
    CascadeMux I__846 (
            .O(N__5207),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_7_i_2_cascade_ ));
    InMux I__845 (
            .O(N__5204),
            .I(N__5201));
    LocalMux I__844 (
            .O(N__5201),
            .I(N__5198));
    Odrv12 I__843 (
            .O(N__5198),
            .I(\U712_CHIP_RAM.N_258 ));
    CascadeMux I__842 (
            .O(N__5195),
            .I(\U712_CHIP_RAM.N_49_cascade_ ));
    InMux I__841 (
            .O(N__5192),
            .I(N__5188));
    CascadeMux I__840 (
            .O(N__5191),
            .I(N__5184));
    LocalMux I__839 (
            .O(N__5188),
            .I(N__5181));
    InMux I__838 (
            .O(N__5187),
            .I(N__5178));
    InMux I__837 (
            .O(N__5184),
            .I(N__5175));
    Span4Mux_v I__836 (
            .O(N__5181),
            .I(N__5172));
    LocalMux I__835 (
            .O(N__5178),
            .I(\U712_CHIP_RAM.N_206 ));
    LocalMux I__834 (
            .O(N__5175),
            .I(\U712_CHIP_RAM.N_206 ));
    Odrv4 I__833 (
            .O(N__5172),
            .I(\U712_CHIP_RAM.N_206 ));
    CascadeMux I__832 (
            .O(N__5165),
            .I(N__5162));
    InMux I__831 (
            .O(N__5162),
            .I(N__5159));
    LocalMux I__830 (
            .O(N__5159),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_1 ));
    InMux I__829 (
            .O(N__5156),
            .I(N__5150));
    InMux I__828 (
            .O(N__5155),
            .I(N__5147));
    CascadeMux I__827 (
            .O(N__5154),
            .I(N__5144));
    CascadeMux I__826 (
            .O(N__5153),
            .I(N__5134));
    LocalMux I__825 (
            .O(N__5150),
            .I(N__5128));
    LocalMux I__824 (
            .O(N__5147),
            .I(N__5128));
    InMux I__823 (
            .O(N__5144),
            .I(N__5123));
    InMux I__822 (
            .O(N__5143),
            .I(N__5123));
    InMux I__821 (
            .O(N__5142),
            .I(N__5119));
    CascadeMux I__820 (
            .O(N__5141),
            .I(N__5114));
    InMux I__819 (
            .O(N__5140),
            .I(N__5110));
    InMux I__818 (
            .O(N__5139),
            .I(N__5105));
    InMux I__817 (
            .O(N__5138),
            .I(N__5105));
    InMux I__816 (
            .O(N__5137),
            .I(N__5102));
    InMux I__815 (
            .O(N__5134),
            .I(N__5097));
    InMux I__814 (
            .O(N__5133),
            .I(N__5097));
    Span4Mux_h I__813 (
            .O(N__5128),
            .I(N__5092));
    LocalMux I__812 (
            .O(N__5123),
            .I(N__5092));
    InMux I__811 (
            .O(N__5122),
            .I(N__5089));
    LocalMux I__810 (
            .O(N__5119),
            .I(N__5086));
    InMux I__809 (
            .O(N__5118),
            .I(N__5081));
    InMux I__808 (
            .O(N__5117),
            .I(N__5081));
    InMux I__807 (
            .O(N__5114),
            .I(N__5076));
    InMux I__806 (
            .O(N__5113),
            .I(N__5076));
    LocalMux I__805 (
            .O(N__5110),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__804 (
            .O(N__5105),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__803 (
            .O(N__5102),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__802 (
            .O(N__5097),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__801 (
            .O(N__5092),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__800 (
            .O(N__5089),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__799 (
            .O(N__5086),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__798 (
            .O(N__5081),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__797 (
            .O(N__5076),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__796 (
            .O(N__5057),
            .I(N__5053));
    InMux I__795 (
            .O(N__5056),
            .I(N__5050));
    LocalMux I__794 (
            .O(N__5053),
            .I(N__5047));
    LocalMux I__793 (
            .O(N__5050),
            .I(N__5038));
    Span4Mux_h I__792 (
            .O(N__5047),
            .I(N__5038));
    InMux I__791 (
            .O(N__5046),
            .I(N__5031));
    InMux I__790 (
            .O(N__5045),
            .I(N__5031));
    InMux I__789 (
            .O(N__5044),
            .I(N__5031));
    InMux I__788 (
            .O(N__5043),
            .I(N__5028));
    Odrv4 I__787 (
            .O(N__5038),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__786 (
            .O(N__5031),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__785 (
            .O(N__5028),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    InMux I__784 (
            .O(N__5021),
            .I(N__5017));
    InMux I__783 (
            .O(N__5020),
            .I(N__5014));
    LocalMux I__782 (
            .O(N__5017),
            .I(N__5011));
    LocalMux I__781 (
            .O(N__5014),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    Odrv4 I__780 (
            .O(N__5011),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__779 (
            .O(N__5006),
            .I(N__5002));
    InMux I__778 (
            .O(N__5005),
            .I(N__4998));
    LocalMux I__777 (
            .O(N__5002),
            .I(N__4995));
    InMux I__776 (
            .O(N__5001),
            .I(N__4992));
    LocalMux I__775 (
            .O(N__4998),
            .I(N__4987));
    Span4Mux_h I__774 (
            .O(N__4995),
            .I(N__4987));
    LocalMux I__773 (
            .O(N__4992),
            .I(\U712_CHIP_RAM.N_167 ));
    Odrv4 I__772 (
            .O(N__4987),
            .I(\U712_CHIP_RAM.N_167 ));
    CascadeMux I__771 (
            .O(N__4982),
            .I(N__4976));
    InMux I__770 (
            .O(N__4981),
            .I(N__4972));
    InMux I__769 (
            .O(N__4980),
            .I(N__4967));
    InMux I__768 (
            .O(N__4979),
            .I(N__4967));
    InMux I__767 (
            .O(N__4976),
            .I(N__4964));
    InMux I__766 (
            .O(N__4975),
            .I(N__4961));
    LocalMux I__765 (
            .O(N__4972),
            .I(N__4956));
    LocalMux I__764 (
            .O(N__4967),
            .I(N__4953));
    LocalMux I__763 (
            .O(N__4964),
            .I(N__4948));
    LocalMux I__762 (
            .O(N__4961),
            .I(N__4948));
    InMux I__761 (
            .O(N__4960),
            .I(N__4943));
    InMux I__760 (
            .O(N__4959),
            .I(N__4943));
    Span4Mux_v I__759 (
            .O(N__4956),
            .I(N__4936));
    Span4Mux_h I__758 (
            .O(N__4953),
            .I(N__4936));
    Span4Mux_v I__757 (
            .O(N__4948),
            .I(N__4936));
    LocalMux I__756 (
            .O(N__4943),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__755 (
            .O(N__4936),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__754 (
            .O(N__4931),
            .I(N__4926));
    InMux I__753 (
            .O(N__4930),
            .I(N__4920));
    InMux I__752 (
            .O(N__4929),
            .I(N__4917));
    LocalMux I__751 (
            .O(N__4926),
            .I(N__4914));
    InMux I__750 (
            .O(N__4925),
            .I(N__4911));
    InMux I__749 (
            .O(N__4924),
            .I(N__4908));
    InMux I__748 (
            .O(N__4923),
            .I(N__4905));
    LocalMux I__747 (
            .O(N__4920),
            .I(N__4902));
    LocalMux I__746 (
            .O(N__4917),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1 ));
    Odrv4 I__745 (
            .O(N__4914),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1 ));
    LocalMux I__744 (
            .O(N__4911),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1 ));
    LocalMux I__743 (
            .O(N__4908),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1 ));
    LocalMux I__742 (
            .O(N__4905),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1 ));
    Odrv4 I__741 (
            .O(N__4902),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1 ));
    InMux I__740 (
            .O(N__4889),
            .I(N__4879));
    InMux I__739 (
            .O(N__4888),
            .I(N__4872));
    InMux I__738 (
            .O(N__4887),
            .I(N__4872));
    InMux I__737 (
            .O(N__4886),
            .I(N__4872));
    InMux I__736 (
            .O(N__4885),
            .I(N__4865));
    InMux I__735 (
            .O(N__4884),
            .I(N__4865));
    InMux I__734 (
            .O(N__4883),
            .I(N__4865));
    InMux I__733 (
            .O(N__4882),
            .I(N__4862));
    LocalMux I__732 (
            .O(N__4879),
            .I(N__4859));
    LocalMux I__731 (
            .O(N__4872),
            .I(\U712_CHIP_RAM.N_53 ));
    LocalMux I__730 (
            .O(N__4865),
            .I(\U712_CHIP_RAM.N_53 ));
    LocalMux I__729 (
            .O(N__4862),
            .I(\U712_CHIP_RAM.N_53 ));
    Odrv4 I__728 (
            .O(N__4859),
            .I(\U712_CHIP_RAM.N_53 ));
    InMux I__727 (
            .O(N__4850),
            .I(N__4847));
    LocalMux I__726 (
            .O(N__4847),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    CascadeMux I__725 (
            .O(N__4844),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_1_cascade_ ));
    CEMux I__724 (
            .O(N__4841),
            .I(N__4837));
    CEMux I__723 (
            .O(N__4840),
            .I(N__4834));
    LocalMux I__722 (
            .O(N__4837),
            .I(N__4830));
    LocalMux I__721 (
            .O(N__4834),
            .I(N__4827));
    CEMux I__720 (
            .O(N__4833),
            .I(N__4824));
    Span4Mux_h I__719 (
            .O(N__4830),
            .I(N__4821));
    Span4Mux_h I__718 (
            .O(N__4827),
            .I(N__4818));
    LocalMux I__717 (
            .O(N__4824),
            .I(N__4815));
    Span4Mux_h I__716 (
            .O(N__4821),
            .I(N__4812));
    Span4Mux_h I__715 (
            .O(N__4818),
            .I(N__4809));
    Span4Mux_v I__714 (
            .O(N__4815),
            .I(N__4806));
    Odrv4 I__713 (
            .O(N__4812),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv4 I__712 (
            .O(N__4809),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv4 I__711 (
            .O(N__4806),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    CascadeMux I__710 (
            .O(N__4799),
            .I(\U712_CHIP_RAM.N_196_cascade_ ));
    InMux I__709 (
            .O(N__4796),
            .I(N__4789));
    InMux I__708 (
            .O(N__4795),
            .I(N__4789));
    InMux I__707 (
            .O(N__4794),
            .I(N__4786));
    LocalMux I__706 (
            .O(N__4789),
            .I(N__4783));
    LocalMux I__705 (
            .O(N__4786),
            .I(\U712_CHIP_RAM.N_315 ));
    Odrv4 I__704 (
            .O(N__4783),
            .I(\U712_CHIP_RAM.N_315 ));
    CascadeMux I__703 (
            .O(N__4778),
            .I(\U712_CHIP_RAM.N_197_i_cascade_ ));
    InMux I__702 (
            .O(N__4775),
            .I(N__4769));
    InMux I__701 (
            .O(N__4774),
            .I(N__4769));
    LocalMux I__700 (
            .O(N__4769),
            .I(N__4766));
    Odrv4 I__699 (
            .O(N__4766),
            .I(\U712_CHIP_RAM.N_233 ));
    InMux I__698 (
            .O(N__4763),
            .I(N__4760));
    LocalMux I__697 (
            .O(N__4760),
            .I(N__4755));
    InMux I__696 (
            .O(N__4759),
            .I(N__4750));
    InMux I__695 (
            .O(N__4758),
            .I(N__4750));
    Odrv4 I__694 (
            .O(N__4755),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8RZ0 ));
    LocalMux I__693 (
            .O(N__4750),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8RZ0 ));
    InMux I__692 (
            .O(N__4745),
            .I(N__4741));
    InMux I__691 (
            .O(N__4744),
            .I(N__4738));
    LocalMux I__690 (
            .O(N__4741),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__689 (
            .O(N__4738),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__688 (
            .O(N__4733),
            .I(N__4729));
    InMux I__687 (
            .O(N__4732),
            .I(N__4726));
    LocalMux I__686 (
            .O(N__4729),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__685 (
            .O(N__4726),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__684 (
            .O(N__4721),
            .I(N__4717));
    InMux I__683 (
            .O(N__4720),
            .I(N__4714));
    InMux I__682 (
            .O(N__4717),
            .I(N__4711));
    LocalMux I__681 (
            .O(N__4714),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__680 (
            .O(N__4711),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__679 (
            .O(N__4706),
            .I(N__4702));
    InMux I__678 (
            .O(N__4705),
            .I(N__4699));
    LocalMux I__677 (
            .O(N__4702),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__676 (
            .O(N__4699),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__675 (
            .O(N__4694),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1_cascade_ ));
    CEMux I__674 (
            .O(N__4691),
            .I(N__4687));
    CEMux I__673 (
            .O(N__4690),
            .I(N__4684));
    LocalMux I__672 (
            .O(N__4687),
            .I(N__4681));
    LocalMux I__671 (
            .O(N__4684),
            .I(N__4678));
    Odrv4 I__670 (
            .O(N__4681),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ));
    Odrv4 I__669 (
            .O(N__4678),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ));
    InMux I__668 (
            .O(N__4673),
            .I(N__4669));
    InMux I__667 (
            .O(N__4672),
            .I(N__4666));
    LocalMux I__666 (
            .O(N__4669),
            .I(N__4662));
    LocalMux I__665 (
            .O(N__4666),
            .I(N__4659));
    InMux I__664 (
            .O(N__4665),
            .I(N__4656));
    Odrv4 I__663 (
            .O(N__4662),
            .I(\U712_CHIP_RAM.N_314 ));
    Odrv4 I__662 (
            .O(N__4659),
            .I(\U712_CHIP_RAM.N_314 ));
    LocalMux I__661 (
            .O(N__4656),
            .I(\U712_CHIP_RAM.N_314 ));
    InMux I__660 (
            .O(N__4649),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__659 (
            .O(N__4646),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__658 (
            .O(N__4643),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__657 (
            .O(N__4640),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__656 (
            .O(N__4637),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__655 (
            .O(N__4634),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__654 (
            .O(N__4631),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    CascadeMux I__653 (
            .O(N__4628),
            .I(\U712_CHIP_RAM.N_230_cascade_ ));
    CascadeMux I__652 (
            .O(N__4625),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_0_cascade_ ));
    InMux I__651 (
            .O(N__4622),
            .I(N__4619));
    LocalMux I__650 (
            .O(N__4619),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_1 ));
    InMux I__649 (
            .O(N__4616),
            .I(N__4613));
    LocalMux I__648 (
            .O(N__4613),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_1 ));
    InMux I__647 (
            .O(N__4610),
            .I(N__4607));
    LocalMux I__646 (
            .O(N__4607),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_a3_1_1 ));
    CascadeMux I__645 (
            .O(N__4604),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_cascade_ ));
    InMux I__644 (
            .O(N__4601),
            .I(N__4598));
    LocalMux I__643 (
            .O(N__4598),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ));
    CascadeMux I__642 (
            .O(N__4595),
            .I(\U712_CHIP_RAM.N_285_cascade_ ));
    CascadeMux I__641 (
            .O(N__4592),
            .I(N__4589));
    InMux I__640 (
            .O(N__4589),
            .I(N__4586));
    LocalMux I__639 (
            .O(N__4586),
            .I(N__4583));
    Odrv4 I__638 (
            .O(N__4583),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_1 ));
    CascadeMux I__637 (
            .O(N__4580),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_1_cascade_ ));
    CascadeMux I__636 (
            .O(N__4577),
            .I(N__4574));
    InMux I__635 (
            .O(N__4574),
            .I(N__4571));
    LocalMux I__634 (
            .O(N__4571),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1 ));
    SRMux I__633 (
            .O(N__4568),
            .I(N__4565));
    LocalMux I__632 (
            .O(N__4565),
            .I(N__4562));
    Span4Mux_h I__631 (
            .O(N__4562),
            .I(N__4559));
    Odrv4 I__630 (
            .O(N__4559),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__629 (
            .O(N__4556),
            .I(N__4553));
    LocalMux I__628 (
            .O(N__4553),
            .I(N__4550));
    Span4Mux_v I__627 (
            .O(N__4550),
            .I(N__4547));
    Span4Mux_h I__626 (
            .O(N__4547),
            .I(N__4544));
    Sp12to4 I__625 (
            .O(N__4544),
            .I(N__4541));
    Odrv12 I__624 (
            .O(N__4541),
            .I(A_c_13));
    CascadeMux I__623 (
            .O(N__4538),
            .I(N__4535));
    InMux I__622 (
            .O(N__4535),
            .I(N__4532));
    LocalMux I__621 (
            .O(N__4532),
            .I(N__4529));
    Span12Mux_v I__620 (
            .O(N__4529),
            .I(N__4526));
    Span12Mux_h I__619 (
            .O(N__4526),
            .I(N__4523));
    Odrv12 I__618 (
            .O(N__4523),
            .I(A_c_6));
    InMux I__617 (
            .O(N__4520),
            .I(N__4517));
    LocalMux I__616 (
            .O(N__4517),
            .I(N__4514));
    Span4Mux_h I__615 (
            .O(N__4514),
            .I(N__4511));
    Sp12to4 I__614 (
            .O(N__4511),
            .I(N__4508));
    Span12Mux_v I__613 (
            .O(N__4508),
            .I(N__4505));
    Odrv12 I__612 (
            .O(N__4505),
            .I(A_c_15));
    InMux I__611 (
            .O(N__4502),
            .I(N__4499));
    LocalMux I__610 (
            .O(N__4499),
            .I(N__4496));
    Span12Mux_v I__609 (
            .O(N__4496),
            .I(N__4493));
    Span12Mux_h I__608 (
            .O(N__4493),
            .I(N__4490));
    Odrv12 I__607 (
            .O(N__4490),
            .I(A_c_8));
    CascadeMux I__606 (
            .O(N__4487),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ));
    InMux I__605 (
            .O(N__4484),
            .I(N__4477));
    InMux I__604 (
            .O(N__4483),
            .I(N__4477));
    InMux I__603 (
            .O(N__4482),
            .I(N__4474));
    LocalMux I__602 (
            .O(N__4477),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIIGLS1Z0Z_0 ));
    LocalMux I__601 (
            .O(N__4474),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIIGLS1Z0Z_0 ));
    CascadeMux I__600 (
            .O(N__4469),
            .I(N__4466));
    InMux I__599 (
            .O(N__4466),
            .I(N__4458));
    InMux I__598 (
            .O(N__4465),
            .I(N__4458));
    InMux I__597 (
            .O(N__4464),
            .I(N__4454));
    InMux I__596 (
            .O(N__4463),
            .I(N__4451));
    LocalMux I__595 (
            .O(N__4458),
            .I(N__4448));
    InMux I__594 (
            .O(N__4457),
            .I(N__4445));
    LocalMux I__593 (
            .O(N__4454),
            .I(N__4440));
    LocalMux I__592 (
            .O(N__4451),
            .I(N__4440));
    Odrv4 I__591 (
            .O(N__4448),
            .I(\U712_CHIP_RAM.N_176 ));
    LocalMux I__590 (
            .O(N__4445),
            .I(\U712_CHIP_RAM.N_176 ));
    Odrv4 I__589 (
            .O(N__4440),
            .I(\U712_CHIP_RAM.N_176 ));
    InMux I__588 (
            .O(N__4433),
            .I(N__4429));
    InMux I__587 (
            .O(N__4432),
            .I(N__4426));
    LocalMux I__586 (
            .O(N__4429),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__585 (
            .O(N__4426),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__584 (
            .O(N__4421),
            .I(\U712_CHIP_RAM.N_167_cascade_ ));
    CEMux I__583 (
            .O(N__4418),
            .I(N__4415));
    LocalMux I__582 (
            .O(N__4415),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_9_0_0 ));
    InMux I__581 (
            .O(N__4412),
            .I(N__4409));
    LocalMux I__580 (
            .O(N__4409),
            .I(N__4405));
    InMux I__579 (
            .O(N__4408),
            .I(N__4402));
    Odrv4 I__578 (
            .O(N__4405),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__577 (
            .O(N__4402),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__576 (
            .O(N__4397),
            .I(N__4388));
    InMux I__575 (
            .O(N__4396),
            .I(N__4388));
    InMux I__574 (
            .O(N__4395),
            .I(N__4388));
    LocalMux I__573 (
            .O(N__4388),
            .I(N__4385));
    Sp12to4 I__572 (
            .O(N__4385),
            .I(N__4382));
    Span12Mux_v I__571 (
            .O(N__4382),
            .I(N__4379));
    Span12Mux_h I__570 (
            .O(N__4379),
            .I(N__4376));
    Odrv12 I__569 (
            .O(N__4376),
            .I(SIZ_c_1));
    IoInMux I__568 (
            .O(N__4373),
            .I(N__4370));
    LocalMux I__567 (
            .O(N__4370),
            .I(N__4367));
    Span4Mux_s0_v I__566 (
            .O(N__4367),
            .I(N__4364));
    Sp12to4 I__565 (
            .O(N__4364),
            .I(N__4360));
    InMux I__564 (
            .O(N__4363),
            .I(N__4357));
    Span12Mux_h I__563 (
            .O(N__4360),
            .I(N__4354));
    LocalMux I__562 (
            .O(N__4357),
            .I(N__4351));
    Odrv12 I__561 (
            .O(N__4354),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__560 (
            .O(N__4351),
            .I(CONSTANT_ONE_NET));
    InMux I__559 (
            .O(N__4346),
            .I(N__4343));
    LocalMux I__558 (
            .O(N__4343),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__557 (
            .O(N__4340),
            .I(N__4337));
    LocalMux I__556 (
            .O(N__4337),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    CascadeMux I__555 (
            .O(N__4334),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1_cascade_ ));
    InMux I__554 (
            .O(N__4331),
            .I(N__4327));
    InMux I__553 (
            .O(N__4330),
            .I(N__4324));
    LocalMux I__552 (
            .O(N__4327),
            .I(\U712_CHIP_RAM.N_313 ));
    LocalMux I__551 (
            .O(N__4324),
            .I(\U712_CHIP_RAM.N_313 ));
    InMux I__550 (
            .O(N__4319),
            .I(N__4316));
    LocalMux I__549 (
            .O(N__4316),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ));
    CascadeMux I__548 (
            .O(N__4313),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_9_0_cascade_ ));
    InMux I__547 (
            .O(N__4310),
            .I(N__4305));
    InMux I__546 (
            .O(N__4309),
            .I(N__4300));
    InMux I__545 (
            .O(N__4308),
            .I(N__4300));
    LocalMux I__544 (
            .O(N__4305),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0_a3_0 ));
    LocalMux I__543 (
            .O(N__4300),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0_a3_0 ));
    CascadeMux I__542 (
            .O(N__4295),
            .I(\U712_CHIP_RAM.N_232_cascade_ ));
    InMux I__541 (
            .O(N__4292),
            .I(N__4289));
    LocalMux I__540 (
            .O(N__4289),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0_a3_1 ));
    InMux I__539 (
            .O(N__4286),
            .I(N__4283));
    LocalMux I__538 (
            .O(N__4283),
            .I(\U712_CHIP_RAM.N_232 ));
    InMux I__537 (
            .O(N__4280),
            .I(N__4276));
    InMux I__536 (
            .O(N__4279),
            .I(N__4273));
    LocalMux I__535 (
            .O(N__4276),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    LocalMux I__534 (
            .O(N__4273),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    InMux I__533 (
            .O(N__4268),
            .I(N__4265));
    LocalMux I__532 (
            .O(N__4265),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0 ));
    InMux I__531 (
            .O(N__4262),
            .I(N__4259));
    LocalMux I__530 (
            .O(N__4259),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_i_i_a3_0 ));
    CascadeMux I__529 (
            .O(N__4256),
            .I(N__4253));
    InMux I__528 (
            .O(N__4253),
            .I(N__4250));
    LocalMux I__527 (
            .O(N__4250),
            .I(N__4247));
    Odrv4 I__526 (
            .O(N__4247),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    CascadeMux I__525 (
            .O(N__4244),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_cascade_ ));
    CascadeMux I__524 (
            .O(N__4241),
            .I(\U712_CHIP_RAM.CLK_EN_e_1_cascade_ ));
    IoInMux I__523 (
            .O(N__4238),
            .I(N__4235));
    LocalMux I__522 (
            .O(N__4235),
            .I(N__4232));
    IoSpan4Mux I__521 (
            .O(N__4232),
            .I(N__4229));
    Sp12to4 I__520 (
            .O(N__4229),
            .I(N__4226));
    Span12Mux_s7_h I__519 (
            .O(N__4226),
            .I(N__4223));
    Span12Mux_h I__518 (
            .O(N__4223),
            .I(N__4219));
    InMux I__517 (
            .O(N__4222),
            .I(N__4216));
    Odrv12 I__516 (
            .O(N__4219),
            .I(CLK_EN_c));
    LocalMux I__515 (
            .O(N__4216),
            .I(CLK_EN_c));
    CascadeMux I__514 (
            .O(N__4211),
            .I(\U712_CHIP_RAM.N_176_cascade_ ));
    CascadeMux I__513 (
            .O(N__4208),
            .I(\U712_CHIP_RAM.N_166_cascade_ ));
    InMux I__512 (
            .O(N__4205),
            .I(N__4202));
    LocalMux I__511 (
            .O(N__4202),
            .I(N__4199));
    Span12Mux_h I__510 (
            .O(N__4199),
            .I(N__4196));
    Odrv12 I__509 (
            .O(N__4196),
            .I(A_c_11));
    InMux I__508 (
            .O(N__4193),
            .I(N__4190));
    LocalMux I__507 (
            .O(N__4190),
            .I(N__4187));
    Span4Mux_h I__506 (
            .O(N__4187),
            .I(N__4184));
    Sp12to4 I__505 (
            .O(N__4184),
            .I(N__4181));
    Span12Mux_v I__504 (
            .O(N__4181),
            .I(N__4178));
    Odrv12 I__503 (
            .O(N__4178),
            .I(A_c_4));
    InMux I__502 (
            .O(N__4175),
            .I(N__4172));
    LocalMux I__501 (
            .O(N__4172),
            .I(N__4169));
    Span4Mux_h I__500 (
            .O(N__4169),
            .I(N__4166));
    Span4Mux_v I__499 (
            .O(N__4166),
            .I(N__4163));
    Sp12to4 I__498 (
            .O(N__4163),
            .I(N__4160));
    Odrv12 I__497 (
            .O(N__4160),
            .I(A_c_9));
    InMux I__496 (
            .O(N__4157),
            .I(N__4154));
    LocalMux I__495 (
            .O(N__4154),
            .I(N__4151));
    Span4Mux_v I__494 (
            .O(N__4151),
            .I(N__4148));
    Sp12to4 I__493 (
            .O(N__4148),
            .I(N__4145));
    Span12Mux_h I__492 (
            .O(N__4145),
            .I(N__4142));
    Span12Mux_v I__491 (
            .O(N__4142),
            .I(N__4139));
    Odrv12 I__490 (
            .O(N__4139),
            .I(A_c_2));
    CascadeMux I__489 (
            .O(N__4136),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_1_cascade_ ));
    InMux I__488 (
            .O(N__4133),
            .I(N__4130));
    LocalMux I__487 (
            .O(N__4130),
            .I(N__4127));
    Span4Mux_v I__486 (
            .O(N__4127),
            .I(N__4124));
    Span4Mux_h I__485 (
            .O(N__4124),
            .I(N__4121));
    Sp12to4 I__484 (
            .O(N__4121),
            .I(N__4118));
    Odrv12 I__483 (
            .O(N__4118),
            .I(A_c_12));
    InMux I__482 (
            .O(N__4115),
            .I(N__4112));
    LocalMux I__481 (
            .O(N__4112),
            .I(N__4109));
    Span4Mux_v I__480 (
            .O(N__4109),
            .I(N__4106));
    Span4Mux_v I__479 (
            .O(N__4106),
            .I(N__4103));
    Sp12to4 I__478 (
            .O(N__4103),
            .I(N__4100));
    Odrv12 I__477 (
            .O(N__4100),
            .I(A_c_5));
    CascadeMux I__476 (
            .O(N__4097),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2_cascade_ ));
    InMux I__475 (
            .O(N__4094),
            .I(N__4091));
    LocalMux I__474 (
            .O(N__4091),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_0 ));
    InMux I__473 (
            .O(N__4088),
            .I(N__4085));
    LocalMux I__472 (
            .O(N__4085),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_1_0 ));
    CascadeMux I__471 (
            .O(N__4082),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_ ));
    InMux I__470 (
            .O(N__4079),
            .I(N__4076));
    LocalMux I__469 (
            .O(N__4076),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_2 ));
    InMux I__468 (
            .O(N__4073),
            .I(N__4070));
    LocalMux I__467 (
            .O(N__4070),
            .I(N__4067));
    Span4Mux_h I__466 (
            .O(N__4067),
            .I(N__4064));
    Sp12to4 I__465 (
            .O(N__4064),
            .I(N__4061));
    Span12Mux_v I__464 (
            .O(N__4061),
            .I(N__4058));
    Odrv12 I__463 (
            .O(N__4058),
            .I(RAMSPACEn_c));
    InMux I__462 (
            .O(N__4055),
            .I(N__4052));
    LocalMux I__461 (
            .O(N__4052),
            .I(N__4049));
    Odrv4 I__460 (
            .O(N__4049),
            .I(\U712_CHIP_RAM.un5_DMA_CYCLE_START_0 ));
    InMux I__459 (
            .O(N__4046),
            .I(N__4042));
    InMux I__458 (
            .O(N__4045),
            .I(N__4039));
    LocalMux I__457 (
            .O(N__4042),
            .I(N__4035));
    LocalMux I__456 (
            .O(N__4039),
            .I(N__4032));
    InMux I__455 (
            .O(N__4038),
            .I(N__4029));
    Odrv12 I__454 (
            .O(N__4035),
            .I(REG_CYCLEm));
    Odrv4 I__453 (
            .O(N__4032),
            .I(REG_CYCLEm));
    LocalMux I__452 (
            .O(N__4029),
            .I(REG_CYCLEm));
    IoInMux I__451 (
            .O(N__4022),
            .I(N__4019));
    LocalMux I__450 (
            .O(N__4019),
            .I(N__4016));
    Span4Mux_s0_v I__449 (
            .O(N__4016),
            .I(N__4013));
    Sp12to4 I__448 (
            .O(N__4013),
            .I(N__4010));
    Span12Mux_s9_h I__447 (
            .O(N__4010),
            .I(N__4007));
    Span12Mux_v I__446 (
            .O(N__4007),
            .I(N__4004));
    Odrv12 I__445 (
            .O(N__4004),
            .I(DRDENn_c));
    InMux I__444 (
            .O(N__4001),
            .I(N__3998));
    LocalMux I__443 (
            .O(N__3998),
            .I(N__3995));
    Span4Mux_h I__442 (
            .O(N__3995),
            .I(N__3992));
    Sp12to4 I__441 (
            .O(N__3992),
            .I(N__3989));
    Span12Mux_v I__440 (
            .O(N__3989),
            .I(N__3986));
    Odrv12 I__439 (
            .O(N__3986),
            .I(A_c_16));
    InMux I__438 (
            .O(N__3983),
            .I(N__3980));
    LocalMux I__437 (
            .O(N__3980),
            .I(N__3977));
    Span4Mux_v I__436 (
            .O(N__3977),
            .I(N__3974));
    Span4Mux_v I__435 (
            .O(N__3974),
            .I(N__3971));
    Sp12to4 I__434 (
            .O(N__3971),
            .I(N__3968));
    Span12Mux_h I__433 (
            .O(N__3968),
            .I(N__3965));
    Odrv12 I__432 (
            .O(N__3965),
            .I(A_c_18));
    InMux I__431 (
            .O(N__3962),
            .I(N__3958));
    InMux I__430 (
            .O(N__3961),
            .I(N__3955));
    LocalMux I__429 (
            .O(N__3958),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__428 (
            .O(N__3955),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__427 (
            .O(N__3950),
            .I(N__3947));
    LocalMux I__426 (
            .O(N__3947),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ));
    CascadeMux I__425 (
            .O(N__3944),
            .I(N__3940));
    InMux I__424 (
            .O(N__3943),
            .I(N__3937));
    InMux I__423 (
            .O(N__3940),
            .I(N__3934));
    LocalMux I__422 (
            .O(N__3937),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__421 (
            .O(N__3934),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__420 (
            .O(N__3929),
            .I(N__3926));
    LocalMux I__419 (
            .O(N__3926),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    IoInMux I__418 (
            .O(N__3923),
            .I(N__3920));
    LocalMux I__417 (
            .O(N__3920),
            .I(N__3917));
    Span12Mux_s4_v I__416 (
            .O(N__3917),
            .I(N__3913));
    InMux I__415 (
            .O(N__3916),
            .I(N__3910));
    Odrv12 I__414 (
            .O(N__3913),
            .I(DBDIR_c));
    LocalMux I__413 (
            .O(N__3910),
            .I(DBDIR_c));
    InMux I__412 (
            .O(N__3905),
            .I(N__3902));
    LocalMux I__411 (
            .O(N__3902),
            .I(N__3899));
    Span4Mux_v I__410 (
            .O(N__3899),
            .I(N__3896));
    Odrv4 I__409 (
            .O(N__3896),
            .I(TACK_EN_i_ess));
    IoInMux I__408 (
            .O(N__3893),
            .I(N__3890));
    LocalMux I__407 (
            .O(N__3890),
            .I(N__3887));
    Span12Mux_s5_v I__406 (
            .O(N__3887),
            .I(N__3884));
    Odrv12 I__405 (
            .O(N__3884),
            .I(VBENn_c));
    InMux I__404 (
            .O(N__3881),
            .I(N__3878));
    LocalMux I__403 (
            .O(N__3878),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1 ));
    CascadeMux I__402 (
            .O(N__3875),
            .I(N__3869));
    InMux I__401 (
            .O(N__3874),
            .I(N__3866));
    InMux I__400 (
            .O(N__3873),
            .I(N__3859));
    InMux I__399 (
            .O(N__3872),
            .I(N__3859));
    InMux I__398 (
            .O(N__3869),
            .I(N__3859));
    LocalMux I__397 (
            .O(N__3866),
            .I(N__3856));
    LocalMux I__396 (
            .O(N__3859),
            .I(N__3853));
    Span12Mux_v I__395 (
            .O(N__3856),
            .I(N__3850));
    Span12Mux_h I__394 (
            .O(N__3853),
            .I(N__3847));
    Span12Mux_h I__393 (
            .O(N__3850),
            .I(N__3842));
    Span12Mux_v I__392 (
            .O(N__3847),
            .I(N__3842));
    Odrv12 I__391 (
            .O(N__3842),
            .I(CLK40_PLL_i));
    InMux I__390 (
            .O(N__3839),
            .I(N__3835));
    InMux I__389 (
            .O(N__3838),
            .I(N__3832));
    LocalMux I__388 (
            .O(N__3835),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    LocalMux I__387 (
            .O(N__3832),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__386 (
            .O(N__3827),
            .I(N__3823));
    InMux I__385 (
            .O(N__3826),
            .I(N__3820));
    LocalMux I__384 (
            .O(N__3823),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    LocalMux I__383 (
            .O(N__3820),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__382 (
            .O(N__3815),
            .I(bfn_7_7_0_));
    InMux I__381 (
            .O(N__3812),
            .I(N__3808));
    InMux I__380 (
            .O(N__3811),
            .I(N__3805));
    LocalMux I__379 (
            .O(N__3808),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    LocalMux I__378 (
            .O(N__3805),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    InMux I__377 (
            .O(N__3800),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__376 (
            .O(N__3797),
            .I(N__3793));
    InMux I__375 (
            .O(N__3796),
            .I(N__3790));
    LocalMux I__374 (
            .O(N__3793),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    LocalMux I__373 (
            .O(N__3790),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    InMux I__372 (
            .O(N__3785),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__371 (
            .O(N__3782),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    CascadeMux I__370 (
            .O(N__3779),
            .I(N__3775));
    InMux I__369 (
            .O(N__3778),
            .I(N__3772));
    InMux I__368 (
            .O(N__3775),
            .I(N__3769));
    LocalMux I__367 (
            .O(N__3772),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__366 (
            .O(N__3769),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__365 (
            .O(N__3764),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__364 (
            .O(N__3761),
            .I(N__3757));
    InMux I__363 (
            .O(N__3760),
            .I(N__3754));
    LocalMux I__362 (
            .O(N__3757),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__361 (
            .O(N__3754),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__360 (
            .O(N__3749),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__359 (
            .O(N__3746),
            .I(N__3742));
    InMux I__358 (
            .O(N__3745),
            .I(N__3739));
    LocalMux I__357 (
            .O(N__3742),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__356 (
            .O(N__3739),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__355 (
            .O(N__3734),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__354 (
            .O(N__3731),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    IoInMux I__353 (
            .O(N__3728),
            .I(N__3725));
    LocalMux I__352 (
            .O(N__3725),
            .I(N__3722));
    Span4Mux_s2_v I__351 (
            .O(N__3722),
            .I(N__3719));
    Span4Mux_v I__350 (
            .O(N__3719),
            .I(N__3716));
    Span4Mux_h I__349 (
            .O(N__3716),
            .I(N__3713));
    Odrv4 I__348 (
            .O(N__3713),
            .I(CLK80_PLL_i_i));
    InMux I__347 (
            .O(N__3710),
            .I(N__3707));
    LocalMux I__346 (
            .O(N__3707),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ));
    InMux I__345 (
            .O(N__3704),
            .I(N__3697));
    InMux I__344 (
            .O(N__3703),
            .I(N__3697));
    InMux I__343 (
            .O(N__3702),
            .I(N__3694));
    LocalMux I__342 (
            .O(N__3697),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__341 (
            .O(N__3694),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    IoInMux I__340 (
            .O(N__3689),
            .I(N__3686));
    LocalMux I__339 (
            .O(N__3686),
            .I(N__3683));
    Span4Mux_s3_h I__338 (
            .O(N__3683),
            .I(N__3680));
    Span4Mux_h I__337 (
            .O(N__3680),
            .I(N__3677));
    Sp12to4 I__336 (
            .O(N__3677),
            .I(N__3674));
    Span12Mux_v I__335 (
            .O(N__3674),
            .I(N__3670));
    InMux I__334 (
            .O(N__3673),
            .I(N__3667));
    Odrv12 I__333 (
            .O(N__3670),
            .I(TACK_OUTn));
    LocalMux I__332 (
            .O(N__3667),
            .I(TACK_OUTn));
    InMux I__331 (
            .O(N__3662),
            .I(N__3650));
    InMux I__330 (
            .O(N__3661),
            .I(N__3650));
    InMux I__329 (
            .O(N__3660),
            .I(N__3650));
    InMux I__328 (
            .O(N__3659),
            .I(N__3650));
    LocalMux I__327 (
            .O(N__3650),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    IoInMux I__326 (
            .O(N__3647),
            .I(N__3644));
    LocalMux I__325 (
            .O(N__3644),
            .I(N__3641));
    Odrv12 I__324 (
            .O(N__3641),
            .I(CLK40_PLL_i_i));
    IoInMux I__323 (
            .O(N__3638),
            .I(N__3635));
    LocalMux I__322 (
            .O(N__3635),
            .I(N__3632));
    Span4Mux_s3_h I__321 (
            .O(N__3632),
            .I(N__3629));
    Span4Mux_v I__320 (
            .O(N__3629),
            .I(N__3626));
    Span4Mux_v I__319 (
            .O(N__3626),
            .I(N__3623));
    Odrv4 I__318 (
            .O(N__3623),
            .I(N_981_i));
    IoInMux I__317 (
            .O(N__3620),
            .I(N__3617));
    LocalMux I__316 (
            .O(N__3617),
            .I(N__3614));
    Span4Mux_s0_v I__315 (
            .O(N__3614),
            .I(N__3611));
    Span4Mux_v I__314 (
            .O(N__3611),
            .I(N__3608));
    Sp12to4 I__313 (
            .O(N__3608),
            .I(N__3605));
    Span12Mux_h I__312 (
            .O(N__3605),
            .I(N__3602));
    Span12Mux_v I__311 (
            .O(N__3602),
            .I(N__3599));
    Odrv12 I__310 (
            .O(N__3599),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__8473));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .I(N__8475));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__8476));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__8471));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__8472));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .I(N__8474));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__8354),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__7208),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__7253),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLK40_OUT_obuf_RNO_LC_1_10_2.C_ON=1'b0;
    defparam CLK40_OUT_obuf_RNO_LC_1_10_2.SEQ_MODE=4'b0000;
    defparam CLK40_OUT_obuf_RNO_LC_1_10_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLK40_OUT_obuf_RNO_LC_1_10_2 (
            .in0(N__3874),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_obuft_RNO_LC_3_13_2.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_3_13_2.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_3_13_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 TACKn_obuft_RNO_LC_3_13_2 (
            .in0(N__3905),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_981_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_5_1_0.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_5_1_0.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_5_1_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_5_1_0 (
            .in0(N__8840),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_6_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_6_7_1 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_6_7_1  (
            .in0(N__3796),
            .in1(N__3811),
            .in2(N__3779),
            .in3(N__3826),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_6_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_6_7_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_6_7_6  (
            .in0(_gnd_net_),
            .in1(N__3745),
            .in2(_gnd_net_),
            .in3(N__3760),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_6_10_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_6_10_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__3702),
            .in2(_gnd_net_),
            .in3(N__3838),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_6_11_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_6_11_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_6_11_0 .LUT_INIT=16'b0011001000110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_6_11_0  (
            .in0(N__3710),
            .in1(N__3659),
            .in2(N__6788),
            .in3(N__6540),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8836),
            .ce(),
            .sr(N__9254));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_6_11_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_6_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_6_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3704),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8836),
            .ce(),
            .sr(N__9254));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_6_11_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_6_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_6_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_6_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3839),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8836),
            .ce(),
            .sr(N__9254));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_6_11_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_6_11_5 .LUT_INIT=16'b1010111110001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_6_11_5  (
            .in0(N__3662),
            .in1(N__3872),
            .in2(N__6542),
            .in3(N__6766),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8836),
            .ce(),
            .sr(N__9254));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_6_11_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_6_11_6 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_6_11_6 .LUT_INIT=16'b1111111110100010;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_6_11_6  (
            .in0(N__3673),
            .in1(N__3661),
            .in2(N__3875),
            .in3(N__3703),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8836),
            .ce(),
            .sr(N__9254));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_6_11_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_6_11_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_6_11_7  (
            .in0(N__3660),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3873),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8836),
            .ce(),
            .sr(N__9254));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__3827),
            .in2(_gnd_net_),
            .in3(N__3815),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__8470),
            .ce(),
            .sr(N__4568));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__3812),
            .in2(_gnd_net_),
            .in3(N__3800),
            .lcout(\U712_CHIP_RAM.REFRESH5lto1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__8470),
            .ce(),
            .sr(N__4568));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__3797),
            .in2(_gnd_net_),
            .in3(N__3785),
            .lcout(\U712_CHIP_RAM.REFRESH5lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__8470),
            .ce(),
            .sr(N__4568));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__3962),
            .in2(_gnd_net_),
            .in3(N__3782),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__8470),
            .ce(),
            .sr(N__4568));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__3778),
            .in2(_gnd_net_),
            .in3(N__3764),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__8470),
            .ce(),
            .sr(N__4568));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__3761),
            .in2(_gnd_net_),
            .in3(N__3749),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__8470),
            .ce(),
            .sr(N__4568));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__3746),
            .in2(_gnd_net_),
            .in3(N__3734),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__8470),
            .ce(),
            .sr(N__4568));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(N__3943),
            .in2(_gnd_net_),
            .in3(N__3731),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8470),
            .ce(),
            .sr(N__4568));
    defparam \U712_CHIP_RAM.REFRESH_LC_7_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_7_8_3 .LUT_INIT=16'b1111001111111011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_7_8_3  (
            .in0(N__3961),
            .in1(N__3950),
            .in2(N__3944),
            .in3(N__3929),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8824),
            .ce(),
            .sr(N__9265));
    defparam \U712_CHIP_RAM.DBDIR_LC_7_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_7_9_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_7_9_2 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_7_9_2  (
            .in0(N__6445),
            .in1(N__3916),
            .in2(_gnd_net_),
            .in3(N__4280),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8829),
            .ce(),
            .sr(N__9260));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_11_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_11_4 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_11_4 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_11_4  (
            .in0(N__8429),
            .in1(N__6765),
            .in2(_gnd_net_),
            .in3(N__6541),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8835),
            .ce(N__6743),
            .sr(N__9244));
    defparam \U712_BUFFERS.un1_VBENn_0_a3_LC_8_5_7 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a3_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a3_LC_8_5_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a3_LC_8_5_7  (
            .in0(N__4046),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7896),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_6 .LUT_INIT=16'b0010101000101011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_6  (
            .in0(N__6060),
            .in1(N__6188),
            .in2(N__6323),
            .in3(N__3881),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_8_3 .LUT_INIT=16'b1100111101000111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_8_3  (
            .in0(N__4959),
            .in1(N__5143),
            .in2(N__6728),
            .in3(N__6380),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_8_6 .LUT_INIT=16'b0100110000001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_8_6  (
            .in0(N__6381),
            .in1(N__8433),
            .in2(N__5154),
            .in3(N__4960),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_i_i_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_9_3 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_9_3  (
            .in0(N__4079),
            .in1(N__5315),
            .in2(N__6396),
            .in3(N__4055),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8825),
            .ce(),
            .sr(N__9255));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_8_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_8_9_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_8_9_4  (
            .in0(N__4930),
            .in1(N__6376),
            .in2(_gnd_net_),
            .in3(N__5133),
            .lcout(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_8_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_8_9_5 .LUT_INIT=16'b1111011111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_LC_8_9_5  (
            .in0(N__4310),
            .in1(N__4673),
            .in2(N__4082),
            .in3(N__5316),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8825),
            .ce(),
            .sr(N__9255));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_9_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_9_7  (
            .in0(N__6181),
            .in1(N__6061),
            .in2(N__5153),
            .in3(N__6316),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_2_LC_8_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_2_LC_8_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_2_LC_8_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_2_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4412),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8830),
            .ce(),
            .sr(N__9245));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_8_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_8_10_3 .LUT_INIT=16'b0101000001010100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_8_10_3  (
            .in0(N__7564),
            .in1(N__7021),
            .in2(N__5933),
            .in3(N__7051),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8830),
            .ce(),
            .sr(N__9245));
    defparam \U712_CHIP_RAM.DBENn_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_8_10_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_8_10_5 .LUT_INIT=16'b1110001011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_8_10_5  (
            .in0(N__5619),
            .in1(N__4268),
            .in2(N__6089),
            .in3(N__8534),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8830),
            .ce(),
            .sr(N__9245));
    defparam \U712_REG_SM.REG_CYCLE_LC_8_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_8_11_2 .LUT_INIT=16'b1010110010101110;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_8_11_2  (
            .in0(N__7489),
            .in1(N__4038),
            .in2(N__7022),
            .in3(N__7511),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8833),
            .ce(),
            .sr(N__9235));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_11_7 .LUT_INIT=16'b0011011100000101;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_11_7  (
            .in0(N__4073),
            .in1(N__7824),
            .in2(N__7616),
            .in3(N__4433),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8833),
            .ce(),
            .sr(N__9235));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_12_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__4408),
            .in2(_gnd_net_),
            .in3(N__5021),
            .lcout(\U712_CHIP_RAM.un5_DMA_CYCLE_START_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_LC_8_14_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_LC_8_14_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a3_LC_8_14_5  (
            .in0(N__5325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4045),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_2  (
            .in0(N__4001),
            .in1(N__3983),
            .in2(_gnd_net_),
            .in3(N__7432),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_6_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_6_4  (
            .in0(N__7396),
            .in1(N__4205),
            .in2(_gnd_net_),
            .in3(N__4193),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(N__4363),
            .in2(_gnd_net_),
            .in3(N__6077),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_6_7  (
            .in0(N__4175),
            .in1(N__4157),
            .in2(_gnd_net_),
            .in3(N__7395),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_7_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__5971),
            .in2(_gnd_net_),
            .in3(N__4094),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_7_2 .LUT_INIT=16'b1111101011111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_7_2  (
            .in0(N__4483),
            .in1(N__4465),
            .in2(N__4136),
            .in3(N__6321),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8817),
            .ce(N__4691),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_4  (
            .in0(N__4133),
            .in1(N__4115),
            .in2(_gnd_net_),
            .in3(N__7391),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_9_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_9_7_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_9_7_5  (
            .in0(N__6054),
            .in1(N__4463),
            .in2(_gnd_net_),
            .in3(N__5240),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_7_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_7_6  (
            .in0(N__6320),
            .in1(N__6055),
            .in2(N__4097),
            .in3(N__5156),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_7_7 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_7_7  (
            .in0(N__5972),
            .in1(N__4088),
            .in2(N__4469),
            .in3(N__4484),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8817),
            .ce(N__4691),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_1  (
            .in0(N__4262),
            .in1(N__4929),
            .in2(N__4256),
            .in3(N__4889),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8820),
            .ce(N__4833),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_9_8_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_9_8_2  (
            .in0(N__4763),
            .in1(N__6305),
            .in2(N__5191),
            .in3(N__5057),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_a3_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_9_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_9_0  (
            .in0(N__6267),
            .in1(N__6175),
            .in2(_gnd_net_),
            .in3(N__4457),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_9_1 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_9_1  (
            .in0(N__6611),
            .in1(N__4222),
            .in2(N__4244),
            .in3(N__6044),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CLK_EN_e_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_9_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_9_2 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_9_9_2  (
            .in0(N__5056),
            .in1(N__4331),
            .in2(N__4241),
            .in3(N__6206),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8822),
            .ce(),
            .sr(N__9246));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_9_9_3 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_9_9_3  (
            .in0(N__6691),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5122),
            .lcout(\U712_CHIP_RAM.N_176 ),
            .ltout(\U712_CHIP_RAM.N_176_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_4_0_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_4_0_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_4_0_LC_9_9_4 .LUT_INIT=16'b0000101000111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_4_0_LC_9_9_4  (
            .in0(N__6266),
            .in1(N__5137),
            .in2(N__4211),
            .in3(N__5239),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_9_9_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__6157),
            .in2(_gnd_net_),
            .in3(N__6265),
            .lcout(\U712_CHIP_RAM.N_166 ),
            .ltout(\U712_CHIP_RAM.N_166_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_9_9_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_9_9_6  (
            .in0(N__6043),
            .in1(N__6692),
            .in2(N__4208),
            .in3(N__6610),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIVLD65_0_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIVLD65_0_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIVLD65_0_LC_9_9_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIVLD65_0_LC_9_9_7  (
            .in0(N__4975),
            .in1(N__6375),
            .in2(N__4334),
            .in3(N__5005),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIH7LR1_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIH7LR1_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIH7LR1_LC_9_10_0 .LUT_INIT=16'b1000010010000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIH7LR1_LC_9_10_0  (
            .in0(N__6695),
            .in1(N__4330),
            .in2(N__6297),
            .in3(N__5043),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR9AQ_3_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR9AQ_3_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR9AQ_3_LC_9_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIR9AQ_3_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__5113),
            .in2(_gnd_net_),
            .in3(N__6151),
            .lcout(\U712_CHIP_RAM.N_313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_10_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_10_2  (
            .in0(N__4665),
            .in1(N__4309),
            .in2(N__5141),
            .in3(N__4319),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_10_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_10_3  (
            .in0(N__9286),
            .in1(_gnd_net_),
            .in2(N__4313),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_9_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_9_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_9_10_4 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__6084),
            .in2(N__6627),
            .in3(N__4308),
            .lcout(\U712_CHIP_RAM.N_232 ),
            .ltout(\U712_CHIP_RAM.N_232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_9_10_5 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_9_10_5  (
            .in0(N__4794),
            .in1(N__8443),
            .in2(N__4295),
            .in3(N__4924),
            .lcout(\U712_CHIP_RAM.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_10_6 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_10_6  (
            .in0(N__6696),
            .in1(N__4292),
            .in2(N__6628),
            .in3(N__5140),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8826),
            .ce(),
            .sr(N__9236));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_10_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__4286),
            .in2(_gnd_net_),
            .in3(N__4279),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_9_11_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__4432),
            .in2(_gnd_net_),
            .in3(N__6493),
            .lcout(\U712_CHIP_RAM.N_167 ),
            .ltout(\U712_CHIP_RAM.N_167_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_11_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_11_2  (
            .in0(N__4981),
            .in1(N__6401),
            .in2(N__4421),
            .in3(N__4931),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8831),
            .ce(N__4418),
            .sr(N__9232));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5020),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8834),
            .ce(),
            .sr(N__9228));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_LC_9_14_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_LC_9_14_1 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_LC_9_14_1  (
            .in0(N__7884),
            .in1(N__8276),
            .in2(_gnd_net_),
            .in3(N__4397),
            .lcout(\U712_BYTE_ENABLE.N_265 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_9_14_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_9_14_3 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_9_14_3  (
            .in0(N__8313),
            .in1(N__5452),
            .in2(N__7914),
            .in3(N__4396),
            .lcout(\U712_BYTE_ENABLE.N_268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_9_14_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_9_14_5 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_9_14_5  (
            .in0(N__8312),
            .in1(N__5451),
            .in2(N__7913),
            .in3(N__4395),
            .lcout(\U712_BYTE_ENABLE.N_272 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_10_4_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_4_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_4_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_5_1 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_5_1  (
            .in0(N__7912),
            .in1(N__4346),
            .in2(N__7454),
            .in3(N__8939),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_6_0 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_6_0  (
            .in0(N__7910),
            .in1(N__4340),
            .in2(N__7431),
            .in3(N__8585),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIIGLS1_0_LC_10_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIIGLS1_0_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIIGLS1_0_LC_10_6_1 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIIGLS1_0_LC_10_6_1  (
            .in0(N__8444),
            .in1(N__6078),
            .in2(_gnd_net_),
            .in3(N__5242),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_RNIIGLS1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_6_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_6_2  (
            .in0(N__8050),
            .in1(N__7366),
            .in2(N__8187),
            .in3(N__8132),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_2_LC_10_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_2_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_2_LC_10_6_3 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_2_LC_10_6_3  (
            .in0(N__8133),
            .in1(N__8051),
            .in2(_gnd_net_),
            .in3(N__7386),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_6_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_6_5  (
            .in0(N__4556),
            .in1(_gnd_net_),
            .in2(N__4538),
            .in3(N__7387),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_6_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_6_6  (
            .in0(N__4520),
            .in1(N__4502),
            .in2(_gnd_net_),
            .in3(N__7367),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_6_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_6_7  (
            .in0(N__7368),
            .in1(N__7911),
            .in2(N__4487),
            .in3(N__9038),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_7_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_7_1  (
            .in0(N__6177),
            .in1(N__6056),
            .in2(_gnd_net_),
            .in3(N__6718),
            .lcout(\U712_CHIP_RAM.N_258 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_7_3 .LUT_INIT=16'b1111111110101011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_7_3  (
            .in0(N__4482),
            .in1(N__4464),
            .in2(N__6322),
            .in3(N__4622),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8814),
            .ce(N__4690),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_10_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_10_7_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_10_7_4  (
            .in0(_gnd_net_),
            .in1(N__6041),
            .in2(_gnd_net_),
            .in3(N__6176),
            .lcout(\U712_CHIP_RAM.N_206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_7_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_7_5  (
            .in0(N__6042),
            .in1(N__5241),
            .in2(_gnd_net_),
            .in3(N__5155),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_230_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_7_6 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_7_6  (
            .in0(N__6719),
            .in1(N__5187),
            .in2(N__4628),
            .in3(N__6312),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_7_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_7_7  (
            .in0(N__5964),
            .in1(_gnd_net_),
            .in2(N__4625),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIGGM16_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIGGM16_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIGGM16_LC_10_8_0 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIGGM16_LC_10_8_0  (
            .in0(N__4980),
            .in1(N__4923),
            .in2(N__4592),
            .in3(N__6403),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_1  (
            .in0(N__8436),
            .in1(N__4775),
            .in2(N__4577),
            .in3(N__4796),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_8_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_8_2  (
            .in0(N__4672),
            .in1(N__4616),
            .in2(_gnd_net_),
            .in3(N__8437),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_3 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_3  (
            .in0(N__4610),
            .in1(N__6714),
            .in2(N__4604),
            .in3(N__6629),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_285_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_4  (
            .in0(_gnd_net_),
            .in1(N__4601),
            .in2(N__4595),
            .in3(N__8131),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8818),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHHIB1_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHHIB1_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHHIB1_LC_10_8_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHHIB1_LC_10_8_5  (
            .in0(N__8438),
            .in1(N__5006),
            .in2(_gnd_net_),
            .in3(N__5142),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIGNOI5_LC_10_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIGNOI5_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIGNOI5_LC_10_8_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIGNOI5_LC_10_8_6  (
            .in0(N__4979),
            .in1(N__6402),
            .in2(N__4580),
            .in3(N__6202),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITE99E_3_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITE99E_3_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITE99E_3_LC_10_8_7 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITE99E_3_LC_10_8_7  (
            .in0(N__8439),
            .in1(N__4774),
            .in2(N__4694),
            .in3(N__4795),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_10_9_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_10_9_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__6053),
            .in2(_gnd_net_),
            .in3(N__6615),
            .lcout(\U712_CHIP_RAM.N_314 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_9_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_9_1  (
            .in0(N__4886),
            .in1(N__6707),
            .in2(_gnd_net_),
            .in3(N__4649),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__8821),
            .ce(N__4840),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_9_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__6295),
            .in2(_gnd_net_),
            .in3(N__4646),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_9_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_9_3  (
            .in0(N__4887),
            .in1(N__6185),
            .in2(_gnd_net_),
            .in3(N__4643),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__8821),
            .ce(N__4840),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_9_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_9_4  (
            .in0(N__4883),
            .in1(N__4706),
            .in2(_gnd_net_),
            .in3(N__4640),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__8821),
            .ce(N__4840),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_9_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_9_5  (
            .in0(N__4888),
            .in1(N__4733),
            .in2(_gnd_net_),
            .in3(N__4637),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__8821),
            .ce(N__4840),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_9_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_9_6  (
            .in0(N__4884),
            .in1(N__4720),
            .in2(_gnd_net_),
            .in3(N__4634),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__8821),
            .ce(N__4840),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_9_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_9_7  (
            .in0(N__4745),
            .in1(N__4885),
            .in2(_gnd_net_),
            .in3(N__4631),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8821),
            .ce(N__4840),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIVLD65_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIVLD65_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIVLD65_LC_10_10_0 .LUT_INIT=16'b1100110100000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIVLD65_LC_10_10_0  (
            .in0(N__5001),
            .in1(N__6404),
            .in2(N__4982),
            .in3(N__4925),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_10_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_10_1  (
            .in0(N__4882),
            .in1(N__4850),
            .in2(N__4844),
            .in3(N__4759),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8823),
            .ce(N__4841),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_10_10_2 .LUT_INIT=16'b0001000000001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_10_10_2  (
            .in0(N__5118),
            .in1(N__6694),
            .in2(N__6187),
            .in3(N__6269),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_196_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_10_10_3 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__6079),
            .in2(N__4799),
            .in3(N__6613),
            .lcout(\U712_CHIP_RAM.N_315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_10_10_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__6693),
            .in2(_gnd_net_),
            .in3(N__6268),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_197_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_10_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_10_10_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_10_10_5  (
            .in0(N__6161),
            .in1(N__4758),
            .in2(N__4778),
            .in3(N__6614),
            .lcout(\U712_CHIP_RAM.N_233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_10_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_10_6  (
            .in0(N__5117),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8435),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8RZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_10_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_10_7  (
            .in0(N__4744),
            .in1(N__4732),
            .in2(N__4721),
            .in3(N__4705),
            .lcout(\U712_CHIP_RAM.N_165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_6_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_6_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_6_LC_10_11_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_6_LC_10_11_0  (
            .in0(_gnd_net_),
            .in1(N__5044),
            .in2(_gnd_net_),
            .in3(N__6720),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_219_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_11_1 .LUT_INIT=16'b1101110111010101;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_11_1  (
            .in0(N__5138),
            .in1(N__6186),
            .in2(N__5249),
            .in3(N__6296),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_7_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_11_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_11_2  (
            .in0(N__5246),
            .in1(N__5963),
            .in2(N__5207),
            .in3(N__5204),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_49_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_10_11_3 .LUT_INIT=16'b1100111111001010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_10_11_3  (
            .in0(N__6098),
            .in1(N__6556),
            .in2(N__5195),
            .in3(N__6563),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8827),
            .ce(),
            .sr(N__9229));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_5_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_5_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_5_LC_10_11_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_5_LC_10_11_5  (
            .in0(N__5045),
            .in1(N__5192),
            .in2(N__6298),
            .in3(N__7811),
            .lcout(\U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_10_11_6 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_10_11_6  (
            .in0(N__6332),
            .in1(N__5046),
            .in2(N__5165),
            .in3(N__5139),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8827),
            .ce(),
            .sr(N__9229));
    defparam DBR_SYNC_1_LC_10_12_0.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_10_12_0.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_10_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_10_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6962),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8832),
            .ce(),
            .sr(N__9222));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_12_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_12_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_10_12_6  (
            .in0(N__5526),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5390),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8832),
            .ce(),
            .sr(N__9222));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0_0_LC_10_13_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0_0_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0_0_LC_10_13_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0_0_LC_10_13_2  (
            .in0(N__5334),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5634),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0_0_LC_10_13_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0_0_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0_0_LC_10_13_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0_0_LC_10_13_3  (
            .in0(N__5635),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5335),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_185_i_LC_10_14_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_185_i_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_185_i_LC_10_14_0 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \U712_BYTE_ENABLE.N_185_i_LC_10_14_0  (
            .in0(N__5402),
            .in1(N__5415),
            .in2(N__5539),
            .in3(N__5603),
            .lcout(N_185_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_10_14_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_10_14_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_10_14_2  (
            .in0(N__5458),
            .in1(N__8326),
            .in2(_gnd_net_),
            .in3(N__7885),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_270_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_186_i_LC_10_14_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_186_i_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_186_i_LC_10_14_3 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_186_i_LC_10_14_3  (
            .in0(N__5416),
            .in1(N__5488),
            .in2(N__5573),
            .in3(N__5389),
            .lcout(N_186_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_187_i_LC_10_14_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_187_i_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_187_i_LC_10_14_5 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \U712_BYTE_ENABLE.N_187_i_LC_10_14_5  (
            .in0(N__5417),
            .in1(N__5546),
            .in2(N__5540),
            .in3(N__5489),
            .lcout(N_187_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_10_14_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_10_14_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_10_14_6  (
            .in0(N__5459),
            .in1(N__8327),
            .in2(_gnd_net_),
            .in3(N__7886),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_266_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_184_i_LC_10_14_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_184_i_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_184_i_LC_10_14_7 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_184_i_LC_10_14_7  (
            .in0(N__5414),
            .in1(N__5401),
            .in2(N__5393),
            .in3(N__5388),
            .lcout(N_184_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_10_20_3 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_10_20_3 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_m2_LC_10_20_3  (
            .in0(N__6481),
            .in1(N__6444),
            .in2(_gnd_net_),
            .in3(N__5342),
            .lcout(DRDDIR_i_m2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_5_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_11_5_0  (
            .in0(N__7306),
            .in1(N__8573),
            .in2(N__6884),
            .in3(N__5276),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8806),
            .ce(N__8724),
            .sr(N__9261));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_5_3 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_11_5_3  (
            .in0(N__7307),
            .in1(N__6881),
            .in2(N__9410),
            .in3(N__5747),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8806),
            .ce(N__8724),
            .sr(N__9261));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_6_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_11_6_0  (
            .in0(N__7299),
            .in1(N__7274),
            .in2(N__6882),
            .in3(N__5720),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8808),
            .ce(N__8703),
            .sr(N__9256));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_6_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_6_3  (
            .in0(N__7920),
            .in1(N__5690),
            .in2(N__7464),
            .in3(N__9092),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_6_4 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_11_6_4  (
            .in0(N__7298),
            .in1(N__6871),
            .in2(N__5684),
            .in3(N__7265),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8808),
            .ce(N__8703),
            .sr(N__9256));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_0 .LUT_INIT=16'b1111001110111011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_0  (
            .in0(N__8669),
            .in1(N__7956),
            .in2(N__5915),
            .in3(N__7888),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_7_1 .LUT_INIT=16'b0000000000111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_7_1  (
            .in0(N__8126),
            .in1(N__8064),
            .in2(N__7445),
            .in3(N__8181),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_7_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_7_2  (
            .in0(N__9287),
            .in1(_gnd_net_),
            .in2(N__5657),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_2_LC_11_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_2_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_2_LC_11_7_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_2_LC_11_7_4  (
            .in0(N__8063),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8127),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_7_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_7_5  (
            .in0(N__7890),
            .in1(N__5654),
            .in2(N__7446),
            .in3(N__8630),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_7 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_7  (
            .in0(N__7889),
            .in1(N__5911),
            .in2(N__7965),
            .in3(N__8668),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_8_1 .LUT_INIT=16'b0011001011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_8_1  (
            .in0(N__8978),
            .in1(N__6859),
            .in2(N__7919),
            .in3(N__7449),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_8_2 .LUT_INIT=16'b0101001001010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_8_2  (
            .in0(N__7448),
            .in1(N__7902),
            .in2(N__6877),
            .in3(N__8977),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_8_3  (
            .in0(N__5888),
            .in1(N__5867),
            .in2(_gnd_net_),
            .in3(N__7450),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_8_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_8_4  (
            .in0(N__7451),
            .in1(N__7903),
            .in2(N__5849),
            .in3(N__9026),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_11_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_11_8_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__5846),
            .in2(N__5840),
            .in3(N__5837),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8815),
            .ce(N__8704),
            .sr(N__9237));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_11_8_7  (
            .in0(N__5813),
            .in1(N__5804),
            .in2(_gnd_net_),
            .in3(N__5753),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8815),
            .ce(N__8704),
            .sr(N__9237));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_11_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_11_9_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_11_9_0  (
            .in0(N__5774),
            .in1(N__7898),
            .in2(_gnd_net_),
            .in3(N__8594),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_324_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_9_1 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__6876),
            .in2(N__5756),
            .in3(N__7452),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_11_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_11_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_11_9_2  (
            .in0(N__6482),
            .in1(N__6449),
            .in2(_gnd_net_),
            .in3(N__6397),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_1_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_1_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_1_LC_11_9_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_1_LC_11_9_5  (
            .in0(N__6697),
            .in1(N__6273),
            .in2(N__6088),
            .in3(N__6612),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_9_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__7897),
            .in2(N__6191),
            .in3(N__6171),
            .lcout(\U712_CHIP_RAM.N_248 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_11_10_0 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_11_10_0  (
            .in0(N__6080),
            .in1(N__6701),
            .in2(_gnd_net_),
            .in3(N__6616),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_0_2_LC_11_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_0_2_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_0_2_LC_11_10_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI9DCD1_0_2_LC_11_10_1  (
            .in0(N__7218),
            .in1(N__7088),
            .in2(N__7073),
            .in3(N__7166),
            .lcout(\U712_REG_SM.N_171 ),
            .ltout(\U712_REG_SM.N_171_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_11_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_11_10_2 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_11_10_2  (
            .in0(N__7112),
            .in1(_gnd_net_),
            .in2(N__5939),
            .in3(N__7140),
            .lcout(\U712_REG_SM.N_205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIFFTG1_2_LC_11_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIFFTG1_2_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIFFTG1_2_LC_11_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIFFTG1_2_LC_11_10_3  (
            .in0(N__7220),
            .in1(N__7138),
            .in2(N__7175),
            .in3(N__7110),
            .lcout(),
            .ltout(\U712_REG_SM.DS_EN_0_sqmuxa_0_a2_0_a3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_11_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_11_10_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_11_10_4  (
            .in0(N__7090),
            .in1(N__7071),
            .in2(N__5936),
            .in3(N__5932),
            .lcout(\U712_REG_SM.DS_EN_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_11_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_11_10_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_11_10_6  (
            .in0(N__7089),
            .in1(N__7219),
            .in2(N__7174),
            .in3(N__7070),
            .lcout(\U712_REG_SM.N_199 ),
            .ltout(\U712_REG_SM.N_199_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_11_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_11_10_7 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__7111),
            .in2(N__6791),
            .in3(N__7139),
            .lcout(\U712_REG_SM.N_210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_11_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_11_0 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_11_0  (
            .in0(N__8394),
            .in1(N__6787),
            .in2(N__6770),
            .in3(N__6528),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_208_i_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_11_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_11_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6746),
            .in3(N__9285),
            .lcout(\U712_CYCLE_TERM.N_208_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_11_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_11_11_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_11_11_2  (
            .in0(N__6734),
            .in1(N__6727),
            .in2(_gnd_net_),
            .in3(N__6623),
            .lcout(\U712_CHIP_RAM.N_249 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_11_11_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_11_11_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_11_11_3  (
            .in0(N__6973),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6557),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_11_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_11_11_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_11_11_4  (
            .in0(N__7109),
            .in1(N__7741),
            .in2(N__6515),
            .in3(N__7148),
            .lcout(\U712_REG_SM.STATE_COUNT_RNITQLC2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_11_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_11_11_6 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_11_11_6  (
            .in0(N__7108),
            .in1(N__6503),
            .in2(_gnd_net_),
            .in3(N__7147),
            .lcout(\U712_REG_SM.N_174 ),
            .ltout(\U712_REG_SM.N_174_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIBM0G2_2_LC_11_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIBM0G2_2_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIBM0G2_2_LC_11_11_7 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIBM0G2_2_LC_11_11_7  (
            .in0(N__6961),
            .in1(_gnd_net_),
            .in2(N__6497),
            .in3(N__6494),
            .lcout(\U712_REG_SM.N_202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_12_0 .LUT_INIT=16'b1010111000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_11_12_0  (
            .in0(N__7010),
            .in1(N__7033),
            .in2(N__6992),
            .in3(N__7052),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8828),
            .ce(),
            .sr(N__9217));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_12_1 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_11_12_1  (
            .in0(N__7034),
            .in1(N__6988),
            .in2(N__7490),
            .in3(N__7510),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8828),
            .ce(),
            .sr(N__9217));
    defparam \U712_REG_SM.REG_TACK_LC_11_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_11_12_3 .LUT_INIT=16'b1011100010111010;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_11_12_3  (
            .in0(N__7032),
            .in1(N__7011),
            .in2(N__6977),
            .in3(N__6987),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8828),
            .ce(),
            .sr(N__9217));
    defparam DBR_SYNC_0_LC_11_12_5.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_11_12_5.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_11_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_11_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8517),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8828),
            .ce(),
            .sr(N__9217));
    defparam \U712_CHIP_RAM.CASn_LC_12_3_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_12_3_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_12_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7466),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8802),
            .ce(),
            .sr(N__9264));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_5_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_12_5_6  (
            .in0(N__8071),
            .in1(N__7453),
            .in2(N__8144),
            .in3(N__8194),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8803),
            .ce(N__8725),
            .sr(N__9253));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_6_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_6_3  (
            .in0(N__7921),
            .in1(N__6914),
            .in2(N__7465),
            .in3(N__9050),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_6_4 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_12_6_4  (
            .in0(N__7296),
            .in1(N__6872),
            .in2(N__6905),
            .in3(N__9443),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8805),
            .ce(N__8711),
            .sr(N__9243));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_6_7 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_12_6_7  (
            .in0(N__8675),
            .in1(N__7297),
            .in2(N__6883),
            .in3(N__6821),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8805),
            .ce(N__8711),
            .sr(N__9243));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_12_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_12_7_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(N__7887),
            .in2(_gnd_net_),
            .in3(N__7447),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_8_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_8_3  (
            .in0(N__8618),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9388),
            .ce(N__9351),
            .sr(N__9231));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_6  (
            .in0(N__8657),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9388),
            .ce(N__9351),
            .sr(N__9231));
    defparam \U712_REG_SM.C3_SYNC_0_LC_12_9_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_12_9_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_12_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7252),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8813),
            .ce(),
            .sr(N__9227));
    defparam \U712_REG_SM.C1_SYNC_2_LC_12_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_2_LC_12_10_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_2_LC_12_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_2_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7072),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8816),
            .ce(),
            .sr(N__9221));
    defparam \U712_REG_SM.C1_SYNC_0_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_12_10_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_12_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7207),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8816),
            .ce(),
            .sr(N__9221));
    defparam \U712_REG_SM.C3_SYNC_1_LC_12_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_12_10_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_12_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7173),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8816),
            .ce(),
            .sr(N__9221));
    defparam \U712_REG_SM.C3_SYNC_2_LC_12_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_2_LC_12_10_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_2_LC_12_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_2_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7141),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8816),
            .ce(),
            .sr(N__9221));
    defparam \U712_REG_SM.C1_SYNC_1_LC_12_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_12_10_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_12_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7091),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8816),
            .ce(),
            .sr(N__9221));
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_12_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_12_11_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_GO_LC_12_11_0  (
            .in0(N__7662),
            .in1(N__7578),
            .in2(N__7730),
            .in3(N__7627),
            .lcout(\U712_REG_SM.REG_CYCLE_GOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8819),
            .ce(),
            .sr(N__9216));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_12_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_12_11_1 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_12_11_1  (
            .in0(N__7580),
            .in1(N__7742),
            .in2(N__7729),
            .in3(N__7663),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8819),
            .ce(),
            .sr(N__9216));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_12_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_12_11_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_12_11_2 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_12_11_2  (
            .in0(N__7725),
            .in1(N__7577),
            .in2(_gnd_net_),
            .in3(N__7560),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8819),
            .ce(),
            .sr(N__9216));
    defparam \U712_REG_SM.REGENn_1_LC_12_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_1_LC_12_11_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_1_LC_12_11_3 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \U712_REG_SM.REGENn_1_LC_12_11_3  (
            .in0(N__7559),
            .in1(N__7677),
            .in2(_gnd_net_),
            .in3(N__7661),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8819),
            .ce(),
            .sr(N__9216));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_12_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_12_11_4 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_12_11_4  (
            .in0(N__7664),
            .in1(N__7536),
            .in2(_gnd_net_),
            .in3(N__7524),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8819),
            .ce(),
            .sr(N__9216));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_12_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_12_11_5 .LUT_INIT=16'b0000101000111011;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_12_11_5  (
            .in0(N__7579),
            .in1(N__7649),
            .in2(N__7628),
            .in3(N__7615),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8819),
            .ce(),
            .sr(N__9216));
    defparam \U712_REG_SM.DS_EN_LC_12_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_12_11_6 .LUT_INIT=16'b0000101100001010;
    LogicCell40 \U712_REG_SM.DS_EN_LC_12_11_6  (
            .in0(N__8227),
            .in1(N__7525),
            .in2(N__7565),
            .in3(N__7538),
            .lcout(DS_ENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8819),
            .ce(),
            .sr(N__9216));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_11_7 .LUT_INIT=16'b0100111000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_12_11_7  (
            .in0(N__7537),
            .in1(N__7488),
            .in2(N__7526),
            .in3(N__7506),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8819),
            .ce(),
            .sr(N__9216));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_12_7 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_12_7  (
            .in0(N__8518),
            .in1(N__9283),
            .in2(_gnd_net_),
            .in3(N__8480),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_5.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_5.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_17_5 (
            .in0(N__8434),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_12_19_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_12_19_1 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_12_19_1  (
            .in0(N__8236),
            .in1(N__8324),
            .in2(_gnd_net_),
            .in3(N__8268),
            .lcout(N_118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_12_19_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_12_19_4 .LUT_INIT=16'b1010000011111111;
    LogicCell40 \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_12_19_4  (
            .in0(N__8325),
            .in1(_gnd_net_),
            .in2(N__8275),
            .in3(N__8237),
            .lcout(N_113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CRCSn_LC_13_1_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_1_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_13_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8198),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8801),
            .ce(),
            .sr(N__9267));
    defparam \U712_CHIP_RAM.WEn_LC_13_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_13_4_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_13_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_13_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8140),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8804),
            .ce(),
            .sr(N__9266));
    defparam \U712_CHIP_RAM.RASn_LC_13_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_13_5_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_13_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_13_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8072),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8807),
            .ce(),
            .sr(N__9262));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_6_1 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_13_6_1  (
            .in0(N__8009),
            .in1(N__7967),
            .in2(N__7922),
            .in3(N__8852),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8809),
            .ce(N__8729),
            .sr(N__9257));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_6_6 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_13_6_6  (
            .in0(N__7966),
            .in1(N__7943),
            .in2(N__9017),
            .in3(N__7918),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8809),
            .ce(N__8729),
            .sr(N__9257));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9080),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9387),
            .ce(N__9353),
            .sr(N__9247));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9116),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9387),
            .ce(N__9353),
            .sr(N__9247));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_3  (
            .in0(N__8653),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__8922),
            .sr(N__9238));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_0  (
            .in0(N__8617),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__8920),
            .sr(N__9233));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9002),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__8920),
            .sr(N__9233));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_10_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_10_2  (
            .in0(N__8558),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9385),
            .ce(N__9341),
            .sr(N__9230));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8557),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__8904),
            .sr(N__9223));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_13_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_13_12_7 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_13_12_7  (
            .in0(N__8519),
            .in1(N__9284),
            .in2(_gnd_net_),
            .in3(N__9395),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9112),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__8927),
            .sr(N__9258));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_7_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_7_2  (
            .in0(N__9076),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__8927),
            .sr(N__9258));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9431),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__8923),
            .sr(N__9248));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_8_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_8_7  (
            .in0(N__9470),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__8923),
            .sr(N__9248));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8963),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9386),
            .ce(N__9352),
            .sr(N__9239));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_9_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_9_7  (
            .in0(N__8998),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9386),
            .ce(N__9352),
            .sr(N__9239));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8962),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__8921),
            .sr(N__9234));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_7_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_7_0  (
            .in0(N__8870),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9391),
            .ce(N__9355),
            .sr(N__9263));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9469),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9390),
            .ce(N__9359),
            .sr(N__9259));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_9_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_9_4  (
            .in0(N__9427),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9389),
            .ce(N__9354),
            .sr(N__9249));
endmodule // U712_TOP

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 9 2025 19:17:52

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    DRA,
    CMA,
    DA,
    A,
    DBRn,
    RAMENn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    TCIn,
    TBIn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    input [1:0] SIZ;
    input [9:0] DRA;
    output [10:0] CMA;
    output [2:0] DA;
    input [20:0] A;
    input DBRn;
    output RAMENn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    output TCIn;
    output TBIn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__12127;
    wire N__12126;
    wire N__12125;
    wire N__12118;
    wire N__12117;
    wire N__12116;
    wire N__12109;
    wire N__12108;
    wire N__12107;
    wire N__12100;
    wire N__12099;
    wire N__12098;
    wire N__12091;
    wire N__12090;
    wire N__12089;
    wire N__12082;
    wire N__12081;
    wire N__12080;
    wire N__12073;
    wire N__12072;
    wire N__12071;
    wire N__12064;
    wire N__12063;
    wire N__12062;
    wire N__12055;
    wire N__12054;
    wire N__12053;
    wire N__12046;
    wire N__12045;
    wire N__12044;
    wire N__12037;
    wire N__12036;
    wire N__12035;
    wire N__12028;
    wire N__12027;
    wire N__12026;
    wire N__12019;
    wire N__12018;
    wire N__12017;
    wire N__12010;
    wire N__12009;
    wire N__12008;
    wire N__12001;
    wire N__12000;
    wire N__11999;
    wire N__11992;
    wire N__11991;
    wire N__11990;
    wire N__11983;
    wire N__11982;
    wire N__11981;
    wire N__11974;
    wire N__11973;
    wire N__11972;
    wire N__11965;
    wire N__11964;
    wire N__11963;
    wire N__11956;
    wire N__11955;
    wire N__11954;
    wire N__11947;
    wire N__11946;
    wire N__11945;
    wire N__11938;
    wire N__11937;
    wire N__11936;
    wire N__11929;
    wire N__11928;
    wire N__11927;
    wire N__11920;
    wire N__11919;
    wire N__11918;
    wire N__11911;
    wire N__11910;
    wire N__11909;
    wire N__11902;
    wire N__11901;
    wire N__11900;
    wire N__11893;
    wire N__11892;
    wire N__11891;
    wire N__11884;
    wire N__11883;
    wire N__11882;
    wire N__11875;
    wire N__11874;
    wire N__11873;
    wire N__11866;
    wire N__11865;
    wire N__11864;
    wire N__11857;
    wire N__11856;
    wire N__11855;
    wire N__11848;
    wire N__11847;
    wire N__11846;
    wire N__11839;
    wire N__11838;
    wire N__11837;
    wire N__11830;
    wire N__11829;
    wire N__11828;
    wire N__11821;
    wire N__11820;
    wire N__11819;
    wire N__11812;
    wire N__11811;
    wire N__11810;
    wire N__11803;
    wire N__11802;
    wire N__11801;
    wire N__11794;
    wire N__11793;
    wire N__11792;
    wire N__11785;
    wire N__11784;
    wire N__11783;
    wire N__11776;
    wire N__11775;
    wire N__11774;
    wire N__11767;
    wire N__11766;
    wire N__11765;
    wire N__11758;
    wire N__11757;
    wire N__11756;
    wire N__11749;
    wire N__11748;
    wire N__11747;
    wire N__11740;
    wire N__11739;
    wire N__11738;
    wire N__11731;
    wire N__11730;
    wire N__11729;
    wire N__11722;
    wire N__11721;
    wire N__11720;
    wire N__11713;
    wire N__11712;
    wire N__11711;
    wire N__11704;
    wire N__11703;
    wire N__11702;
    wire N__11695;
    wire N__11694;
    wire N__11693;
    wire N__11686;
    wire N__11685;
    wire N__11684;
    wire N__11677;
    wire N__11676;
    wire N__11675;
    wire N__11668;
    wire N__11667;
    wire N__11666;
    wire N__11659;
    wire N__11658;
    wire N__11657;
    wire N__11650;
    wire N__11649;
    wire N__11648;
    wire N__11641;
    wire N__11640;
    wire N__11639;
    wire N__11632;
    wire N__11631;
    wire N__11630;
    wire N__11623;
    wire N__11622;
    wire N__11621;
    wire N__11614;
    wire N__11613;
    wire N__11612;
    wire N__11605;
    wire N__11604;
    wire N__11603;
    wire N__11596;
    wire N__11595;
    wire N__11594;
    wire N__11587;
    wire N__11586;
    wire N__11585;
    wire N__11578;
    wire N__11577;
    wire N__11576;
    wire N__11569;
    wire N__11568;
    wire N__11567;
    wire N__11560;
    wire N__11559;
    wire N__11558;
    wire N__11551;
    wire N__11550;
    wire N__11549;
    wire N__11542;
    wire N__11541;
    wire N__11540;
    wire N__11533;
    wire N__11532;
    wire N__11531;
    wire N__11524;
    wire N__11523;
    wire N__11522;
    wire N__11515;
    wire N__11514;
    wire N__11513;
    wire N__11506;
    wire N__11505;
    wire N__11504;
    wire N__11497;
    wire N__11496;
    wire N__11495;
    wire N__11488;
    wire N__11487;
    wire N__11486;
    wire N__11479;
    wire N__11478;
    wire N__11477;
    wire N__11470;
    wire N__11469;
    wire N__11468;
    wire N__11461;
    wire N__11460;
    wire N__11459;
    wire N__11452;
    wire N__11451;
    wire N__11450;
    wire N__11443;
    wire N__11442;
    wire N__11441;
    wire N__11434;
    wire N__11433;
    wire N__11432;
    wire N__11425;
    wire N__11424;
    wire N__11423;
    wire N__11416;
    wire N__11415;
    wire N__11414;
    wire N__11407;
    wire N__11406;
    wire N__11405;
    wire N__11398;
    wire N__11397;
    wire N__11396;
    wire N__11389;
    wire N__11388;
    wire N__11387;
    wire N__11380;
    wire N__11379;
    wire N__11378;
    wire N__11371;
    wire N__11370;
    wire N__11369;
    wire N__11362;
    wire N__11361;
    wire N__11360;
    wire N__11353;
    wire N__11352;
    wire N__11351;
    wire N__11344;
    wire N__11343;
    wire N__11342;
    wire N__11335;
    wire N__11334;
    wire N__11333;
    wire N__11326;
    wire N__11325;
    wire N__11324;
    wire N__11317;
    wire N__11316;
    wire N__11315;
    wire N__11308;
    wire N__11307;
    wire N__11306;
    wire N__11299;
    wire N__11298;
    wire N__11297;
    wire N__11290;
    wire N__11289;
    wire N__11288;
    wire N__11281;
    wire N__11280;
    wire N__11279;
    wire N__11262;
    wire N__11259;
    wire N__11256;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11243;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11235;
    wire N__11232;
    wire N__11231;
    wire N__11226;
    wire N__11223;
    wire N__11220;
    wire N__11217;
    wire N__11216;
    wire N__11215;
    wire N__11214;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11202;
    wire N__11199;
    wire N__11196;
    wire N__11191;
    wire N__11178;
    wire N__11175;
    wire N__11174;
    wire N__11171;
    wire N__11170;
    wire N__11169;
    wire N__11166;
    wire N__11163;
    wire N__11160;
    wire N__11157;
    wire N__11156;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11144;
    wire N__11139;
    wire N__11134;
    wire N__11129;
    wire N__11124;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11082;
    wire N__11079;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11058;
    wire N__11055;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11031;
    wire N__11028;
    wire N__11025;
    wire N__11024;
    wire N__11023;
    wire N__11020;
    wire N__11019;
    wire N__11018;
    wire N__11015;
    wire N__11014;
    wire N__11011;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10990;
    wire N__10987;
    wire N__10986;
    wire N__10979;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10950;
    wire N__10949;
    wire N__10948;
    wire N__10947;
    wire N__10940;
    wire N__10937;
    wire N__10936;
    wire N__10935;
    wire N__10934;
    wire N__10933;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10917;
    wire N__10914;
    wire N__10909;
    wire N__10906;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10884;
    wire N__10883;
    wire N__10882;
    wire N__10881;
    wire N__10878;
    wire N__10875;
    wire N__10874;
    wire N__10873;
    wire N__10870;
    wire N__10869;
    wire N__10866;
    wire N__10865;
    wire N__10864;
    wire N__10859;
    wire N__10854;
    wire N__10851;
    wire N__10844;
    wire N__10841;
    wire N__10834;
    wire N__10829;
    wire N__10826;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10812;
    wire N__10811;
    wire N__10808;
    wire N__10807;
    wire N__10806;
    wire N__10803;
    wire N__10802;
    wire N__10799;
    wire N__10792;
    wire N__10789;
    wire N__10782;
    wire N__10781;
    wire N__10780;
    wire N__10779;
    wire N__10776;
    wire N__10773;
    wire N__10770;
    wire N__10767;
    wire N__10764;
    wire N__10757;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10737;
    wire N__10736;
    wire N__10733;
    wire N__10730;
    wire N__10729;
    wire N__10728;
    wire N__10725;
    wire N__10722;
    wire N__10719;
    wire N__10716;
    wire N__10713;
    wire N__10710;
    wire N__10707;
    wire N__10702;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10686;
    wire N__10685;
    wire N__10684;
    wire N__10681;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10668;
    wire N__10663;
    wire N__10660;
    wire N__10657;
    wire N__10654;
    wire N__10647;
    wire N__10644;
    wire N__10641;
    wire N__10638;
    wire N__10635;
    wire N__10632;
    wire N__10629;
    wire N__10628;
    wire N__10625;
    wire N__10624;
    wire N__10623;
    wire N__10620;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10612;
    wire N__10611;
    wire N__10610;
    wire N__10609;
    wire N__10608;
    wire N__10607;
    wire N__10604;
    wire N__10603;
    wire N__10602;
    wire N__10601;
    wire N__10600;
    wire N__10599;
    wire N__10598;
    wire N__10593;
    wire N__10590;
    wire N__10587;
    wire N__10584;
    wire N__10581;
    wire N__10578;
    wire N__10573;
    wire N__10572;
    wire N__10569;
    wire N__10564;
    wire N__10561;
    wire N__10556;
    wire N__10551;
    wire N__10550;
    wire N__10549;
    wire N__10546;
    wire N__10545;
    wire N__10540;
    wire N__10537;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10518;
    wire N__10513;
    wire N__10510;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10488;
    wire N__10483;
    wire N__10478;
    wire N__10471;
    wire N__10468;
    wire N__10465;
    wire N__10462;
    wire N__10457;
    wire N__10454;
    wire N__10449;
    wire N__10446;
    wire N__10443;
    wire N__10440;
    wire N__10437;
    wire N__10434;
    wire N__10433;
    wire N__10430;
    wire N__10429;
    wire N__10426;
    wire N__10423;
    wire N__10420;
    wire N__10417;
    wire N__10416;
    wire N__10411;
    wire N__10408;
    wire N__10405;
    wire N__10402;
    wire N__10399;
    wire N__10396;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10374;
    wire N__10371;
    wire N__10368;
    wire N__10365;
    wire N__10364;
    wire N__10363;
    wire N__10362;
    wire N__10361;
    wire N__10360;
    wire N__10359;
    wire N__10344;
    wire N__10341;
    wire N__10338;
    wire N__10337;
    wire N__10336;
    wire N__10335;
    wire N__10334;
    wire N__10333;
    wire N__10332;
    wire N__10331;
    wire N__10330;
    wire N__10329;
    wire N__10328;
    wire N__10327;
    wire N__10326;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10292;
    wire N__10291;
    wire N__10290;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10273;
    wire N__10272;
    wire N__10271;
    wire N__10270;
    wire N__10269;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10261;
    wire N__10260;
    wire N__10259;
    wire N__10258;
    wire N__10257;
    wire N__10256;
    wire N__10255;
    wire N__10254;
    wire N__10253;
    wire N__10250;
    wire N__10249;
    wire N__10248;
    wire N__10247;
    wire N__10246;
    wire N__10245;
    wire N__10244;
    wire N__10243;
    wire N__10240;
    wire N__10239;
    wire N__10238;
    wire N__10237;
    wire N__10236;
    wire N__10233;
    wire N__10232;
    wire N__10231;
    wire N__10230;
    wire N__10229;
    wire N__10228;
    wire N__10227;
    wire N__10226;
    wire N__10225;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10131;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10117;
    wire N__10114;
    wire N__10111;
    wire N__10108;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10086;
    wire N__10083;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10072;
    wire N__10069;
    wire N__10068;
    wire N__10065;
    wire N__10062;
    wire N__10059;
    wire N__10056;
    wire N__10053;
    wire N__10050;
    wire N__10045;
    wire N__10040;
    wire N__10037;
    wire N__10032;
    wire N__10029;
    wire N__10028;
    wire N__10025;
    wire N__10024;
    wire N__10021;
    wire N__10020;
    wire N__10019;
    wire N__10016;
    wire N__10011;
    wire N__10008;
    wire N__10005;
    wire N__10004;
    wire N__9997;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9975;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9967;
    wire N__9966;
    wire N__9965;
    wire N__9964;
    wire N__9963;
    wire N__9962;
    wire N__9961;
    wire N__9960;
    wire N__9959;
    wire N__9954;
    wire N__9953;
    wire N__9952;
    wire N__9951;
    wire N__9950;
    wire N__9947;
    wire N__9946;
    wire N__9945;
    wire N__9942;
    wire N__9939;
    wire N__9938;
    wire N__9937;
    wire N__9936;
    wire N__9933;
    wire N__9932;
    wire N__9925;
    wire N__9922;
    wire N__9919;
    wire N__9918;
    wire N__9915;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9895;
    wire N__9892;
    wire N__9889;
    wire N__9886;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9863;
    wire N__9854;
    wire N__9849;
    wire N__9846;
    wire N__9839;
    wire N__9836;
    wire N__9831;
    wire N__9822;
    wire N__9819;
    wire N__9814;
    wire N__9805;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9789;
    wire N__9788;
    wire N__9787;
    wire N__9786;
    wire N__9783;
    wire N__9782;
    wire N__9781;
    wire N__9780;
    wire N__9779;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9765;
    wire N__9760;
    wire N__9759;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9745;
    wire N__9744;
    wire N__9743;
    wire N__9742;
    wire N__9741;
    wire N__9740;
    wire N__9739;
    wire N__9738;
    wire N__9733;
    wire N__9726;
    wire N__9721;
    wire N__9718;
    wire N__9717;
    wire N__9714;
    wire N__9711;
    wire N__9706;
    wire N__9699;
    wire N__9698;
    wire N__9697;
    wire N__9696;
    wire N__9695;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9672;
    wire N__9667;
    wire N__9662;
    wire N__9657;
    wire N__9654;
    wire N__9633;
    wire N__9630;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9603;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9591;
    wire N__9588;
    wire N__9587;
    wire N__9586;
    wire N__9583;
    wire N__9582;
    wire N__9579;
    wire N__9576;
    wire N__9573;
    wire N__9570;
    wire N__9565;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9549;
    wire N__9546;
    wire N__9543;
    wire N__9540;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9528;
    wire N__9525;
    wire N__9522;
    wire N__9519;
    wire N__9516;
    wire N__9513;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9501;
    wire N__9498;
    wire N__9495;
    wire N__9494;
    wire N__9493;
    wire N__9490;
    wire N__9487;
    wire N__9486;
    wire N__9483;
    wire N__9478;
    wire N__9475;
    wire N__9472;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9450;
    wire N__9447;
    wire N__9444;
    wire N__9441;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9431;
    wire N__9430;
    wire N__9429;
    wire N__9426;
    wire N__9423;
    wire N__9420;
    wire N__9417;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9395;
    wire N__9390;
    wire N__9387;
    wire N__9386;
    wire N__9383;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9369;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9339;
    wire N__9336;
    wire N__9333;
    wire N__9330;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9309;
    wire N__9306;
    wire N__9303;
    wire N__9300;
    wire N__9297;
    wire N__9296;
    wire N__9295;
    wire N__9294;
    wire N__9291;
    wire N__9286;
    wire N__9283;
    wire N__9278;
    wire N__9275;
    wire N__9270;
    wire N__9267;
    wire N__9264;
    wire N__9261;
    wire N__9258;
    wire N__9255;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9219;
    wire N__9216;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9194;
    wire N__9193;
    wire N__9192;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9174;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9132;
    wire N__9131;
    wire N__9128;
    wire N__9127;
    wire N__9126;
    wire N__9125;
    wire N__9122;
    wire N__9121;
    wire N__9118;
    wire N__9113;
    wire N__9112;
    wire N__9109;
    wire N__9104;
    wire N__9099;
    wire N__9096;
    wire N__9095;
    wire N__9094;
    wire N__9085;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9069;
    wire N__9066;
    wire N__9063;
    wire N__9060;
    wire N__9057;
    wire N__9054;
    wire N__9051;
    wire N__9048;
    wire N__9045;
    wire N__9042;
    wire N__9039;
    wire N__9038;
    wire N__9037;
    wire N__9036;
    wire N__9035;
    wire N__9034;
    wire N__9033;
    wire N__9032;
    wire N__9031;
    wire N__9030;
    wire N__9029;
    wire N__9028;
    wire N__9027;
    wire N__9026;
    wire N__9025;
    wire N__9024;
    wire N__9023;
    wire N__9022;
    wire N__9021;
    wire N__9020;
    wire N__9019;
    wire N__9018;
    wire N__9017;
    wire N__9016;
    wire N__9015;
    wire N__9014;
    wire N__9013;
    wire N__9012;
    wire N__9011;
    wire N__9010;
    wire N__9009;
    wire N__9006;
    wire N__9005;
    wire N__9004;
    wire N__9003;
    wire N__9002;
    wire N__9001;
    wire N__9000;
    wire N__8999;
    wire N__8998;
    wire N__8997;
    wire N__8916;
    wire N__8913;
    wire N__8912;
    wire N__8909;
    wire N__8908;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8898;
    wire N__8895;
    wire N__8892;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8880;
    wire N__8877;
    wire N__8872;
    wire N__8869;
    wire N__8866;
    wire N__8859;
    wire N__8858;
    wire N__8853;
    wire N__8850;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8838;
    wire N__8835;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8823;
    wire N__8820;
    wire N__8817;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8809;
    wire N__8804;
    wire N__8801;
    wire N__8796;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8778;
    wire N__8775;
    wire N__8772;
    wire N__8769;
    wire N__8766;
    wire N__8763;
    wire N__8760;
    wire N__8757;
    wire N__8754;
    wire N__8751;
    wire N__8748;
    wire N__8745;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8715;
    wire N__8712;
    wire N__8709;
    wire N__8708;
    wire N__8707;
    wire N__8706;
    wire N__8703;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8689;
    wire N__8686;
    wire N__8683;
    wire N__8680;
    wire N__8679;
    wire N__8672;
    wire N__8669;
    wire N__8664;
    wire N__8663;
    wire N__8662;
    wire N__8659;
    wire N__8656;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8644;
    wire N__8641;
    wire N__8640;
    wire N__8635;
    wire N__8632;
    wire N__8629;
    wire N__8628;
    wire N__8621;
    wire N__8620;
    wire N__8619;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8604;
    wire N__8601;
    wire N__8592;
    wire N__8589;
    wire N__8586;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8574;
    wire N__8571;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8544;
    wire N__8541;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8531;
    wire N__8526;
    wire N__8523;
    wire N__8522;
    wire N__8521;
    wire N__8520;
    wire N__8519;
    wire N__8518;
    wire N__8517;
    wire N__8516;
    wire N__8515;
    wire N__8512;
    wire N__8507;
    wire N__8506;
    wire N__8505;
    wire N__8504;
    wire N__8503;
    wire N__8498;
    wire N__8497;
    wire N__8496;
    wire N__8495;
    wire N__8494;
    wire N__8493;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8482;
    wire N__8481;
    wire N__8476;
    wire N__8473;
    wire N__8470;
    wire N__8467;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8448;
    wire N__8443;
    wire N__8436;
    wire N__8433;
    wire N__8432;
    wire N__8431;
    wire N__8430;
    wire N__8429;
    wire N__8428;
    wire N__8427;
    wire N__8426;
    wire N__8425;
    wire N__8422;
    wire N__8419;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8397;
    wire N__8392;
    wire N__8385;
    wire N__8378;
    wire N__8373;
    wire N__8370;
    wire N__8365;
    wire N__8358;
    wire N__8349;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8331;
    wire N__8328;
    wire N__8325;
    wire N__8322;
    wire N__8319;
    wire N__8316;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8304;
    wire N__8301;
    wire N__8298;
    wire N__8295;
    wire N__8292;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8272;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8259;
    wire N__8252;
    wire N__8247;
    wire N__8244;
    wire N__8241;
    wire N__8238;
    wire N__8235;
    wire N__8232;
    wire N__8231;
    wire N__8228;
    wire N__8227;
    wire N__8226;
    wire N__8225;
    wire N__8224;
    wire N__8221;
    wire N__8218;
    wire N__8213;
    wire N__8208;
    wire N__8199;
    wire N__8198;
    wire N__8197;
    wire N__8196;
    wire N__8195;
    wire N__8194;
    wire N__8193;
    wire N__8192;
    wire N__8189;
    wire N__8188;
    wire N__8187;
    wire N__8180;
    wire N__8179;
    wire N__8178;
    wire N__8175;
    wire N__8172;
    wire N__8169;
    wire N__8164;
    wire N__8159;
    wire N__8156;
    wire N__8151;
    wire N__8148;
    wire N__8133;
    wire N__8132;
    wire N__8129;
    wire N__8128;
    wire N__8127;
    wire N__8126;
    wire N__8125;
    wire N__8124;
    wire N__8121;
    wire N__8118;
    wire N__8109;
    wire N__8106;
    wire N__8097;
    wire N__8096;
    wire N__8095;
    wire N__8094;
    wire N__8093;
    wire N__8090;
    wire N__8089;
    wire N__8088;
    wire N__8083;
    wire N__8078;
    wire N__8075;
    wire N__8070;
    wire N__8067;
    wire N__8058;
    wire N__8055;
    wire N__8052;
    wire N__8049;
    wire N__8048;
    wire N__8047;
    wire N__8044;
    wire N__8043;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8010;
    wire N__8007;
    wire N__8004;
    wire N__8003;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7962;
    wire N__7959;
    wire N__7956;
    wire N__7953;
    wire N__7950;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7917;
    wire N__7914;
    wire N__7911;
    wire N__7908;
    wire N__7905;
    wire N__7902;
    wire N__7899;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7881;
    wire N__7880;
    wire N__7879;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7863;
    wire N__7860;
    wire N__7857;
    wire N__7854;
    wire N__7851;
    wire N__7848;
    wire N__7845;
    wire N__7842;
    wire N__7839;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7831;
    wire N__7826;
    wire N__7823;
    wire N__7818;
    wire N__7815;
    wire N__7812;
    wire N__7809;
    wire N__7808;
    wire N__7807;
    wire N__7804;
    wire N__7801;
    wire N__7798;
    wire N__7797;
    wire N__7790;
    wire N__7787;
    wire N__7782;
    wire N__7779;
    wire N__7778;
    wire N__7773;
    wire N__7772;
    wire N__7771;
    wire N__7770;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7743;
    wire N__7742;
    wire N__7739;
    wire N__7736;
    wire N__7731;
    wire N__7728;
    wire N__7725;
    wire N__7724;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7716;
    wire N__7713;
    wire N__7712;
    wire N__7709;
    wire N__7702;
    wire N__7701;
    wire N__7700;
    wire N__7697;
    wire N__7696;
    wire N__7695;
    wire N__7690;
    wire N__7689;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7665;
    wire N__7662;
    wire N__7647;
    wire N__7644;
    wire N__7641;
    wire N__7640;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7602;
    wire N__7599;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7581;
    wire N__7578;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7548;
    wire N__7545;
    wire N__7542;
    wire N__7539;
    wire N__7536;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7499;
    wire N__7496;
    wire N__7493;
    wire N__7488;
    wire N__7485;
    wire N__7482;
    wire N__7479;
    wire N__7476;
    wire N__7473;
    wire N__7470;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7455;
    wire N__7452;
    wire N__7449;
    wire N__7446;
    wire N__7443;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7428;
    wire N__7425;
    wire N__7422;
    wire N__7419;
    wire N__7418;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7396;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7384;
    wire N__7379;
    wire N__7376;
    wire N__7373;
    wire N__7372;
    wire N__7369;
    wire N__7366;
    wire N__7363;
    wire N__7356;
    wire N__7353;
    wire N__7350;
    wire N__7347;
    wire N__7344;
    wire N__7341;
    wire N__7338;
    wire N__7335;
    wire N__7332;
    wire N__7329;
    wire N__7326;
    wire N__7323;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7311;
    wire N__7308;
    wire N__7305;
    wire N__7302;
    wire N__7299;
    wire N__7296;
    wire N__7293;
    wire N__7290;
    wire N__7287;
    wire N__7284;
    wire N__7281;
    wire N__7278;
    wire N__7275;
    wire N__7272;
    wire N__7269;
    wire N__7266;
    wire N__7263;
    wire N__7260;
    wire N__7257;
    wire N__7254;
    wire N__7251;
    wire N__7248;
    wire N__7245;
    wire N__7242;
    wire N__7239;
    wire N__7236;
    wire N__7233;
    wire N__7230;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7220;
    wire N__7217;
    wire N__7216;
    wire N__7213;
    wire N__7212;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7191;
    wire N__7186;
    wire N__7179;
    wire N__7176;
    wire N__7173;
    wire N__7170;
    wire N__7167;
    wire N__7164;
    wire N__7161;
    wire N__7158;
    wire N__7155;
    wire N__7152;
    wire N__7149;
    wire N__7146;
    wire N__7143;
    wire N__7140;
    wire N__7137;
    wire N__7134;
    wire N__7131;
    wire N__7128;
    wire N__7125;
    wire N__7122;
    wire N__7121;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7113;
    wire N__7110;
    wire N__7107;
    wire N__7104;
    wire N__7101;
    wire N__7100;
    wire N__7099;
    wire N__7094;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7071;
    wire N__7070;
    wire N__7067;
    wire N__7066;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7052;
    wire N__7049;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7029;
    wire N__7028;
    wire N__7023;
    wire N__7020;
    wire N__7017;
    wire N__7014;
    wire N__7011;
    wire N__7008;
    wire N__7005;
    wire N__7002;
    wire N__6999;
    wire N__6996;
    wire N__6993;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6981;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6963;
    wire N__6962;
    wire N__6959;
    wire N__6956;
    wire N__6953;
    wire N__6950;
    wire N__6947;
    wire N__6944;
    wire N__6941;
    wire N__6938;
    wire N__6935;
    wire N__6932;
    wire N__6927;
    wire N__6924;
    wire N__6921;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6902;
    wire N__6901;
    wire N__6900;
    wire N__6899;
    wire N__6898;
    wire N__6897;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6885;
    wire N__6882;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6862;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6852;
    wire N__6847;
    wire N__6844;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6824;
    wire N__6813;
    wire N__6812;
    wire N__6811;
    wire N__6810;
    wire N__6809;
    wire N__6808;
    wire N__6807;
    wire N__6806;
    wire N__6803;
    wire N__6796;
    wire N__6793;
    wire N__6792;
    wire N__6791;
    wire N__6790;
    wire N__6789;
    wire N__6786;
    wire N__6785;
    wire N__6784;
    wire N__6781;
    wire N__6778;
    wire N__6775;
    wire N__6774;
    wire N__6769;
    wire N__6768;
    wire N__6767;
    wire N__6766;
    wire N__6765;
    wire N__6762;
    wire N__6757;
    wire N__6754;
    wire N__6749;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6721;
    wire N__6714;
    wire N__6693;
    wire N__6692;
    wire N__6691;
    wire N__6690;
    wire N__6689;
    wire N__6688;
    wire N__6687;
    wire N__6684;
    wire N__6681;
    wire N__6680;
    wire N__6679;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6667;
    wire N__6660;
    wire N__6659;
    wire N__6658;
    wire N__6657;
    wire N__6654;
    wire N__6653;
    wire N__6652;
    wire N__6651;
    wire N__6648;
    wire N__6645;
    wire N__6642;
    wire N__6639;
    wire N__6634;
    wire N__6631;
    wire N__6626;
    wire N__6619;
    wire N__6616;
    wire N__6597;
    wire N__6596;
    wire N__6595;
    wire N__6594;
    wire N__6591;
    wire N__6588;
    wire N__6587;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6579;
    wire N__6578;
    wire N__6577;
    wire N__6572;
    wire N__6571;
    wire N__6568;
    wire N__6567;
    wire N__6566;
    wire N__6565;
    wire N__6562;
    wire N__6557;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6547;
    wire N__6546;
    wire N__6543;
    wire N__6540;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6520;
    wire N__6513;
    wire N__6498;
    wire N__6495;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6467;
    wire N__6462;
    wire N__6459;
    wire N__6458;
    wire N__6457;
    wire N__6454;
    wire N__6449;
    wire N__6444;
    wire N__6441;
    wire N__6438;
    wire N__6435;
    wire N__6432;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6422;
    wire N__6419;
    wire N__6416;
    wire N__6413;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6377;
    wire N__6374;
    wire N__6371;
    wire N__6368;
    wire N__6363;
    wire N__6360;
    wire N__6357;
    wire N__6354;
    wire N__6351;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6340;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6324;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6302;
    wire N__6299;
    wire N__6294;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6286;
    wire N__6281;
    wire N__6278;
    wire N__6277;
    wire N__6274;
    wire N__6271;
    wire N__6268;
    wire N__6261;
    wire N__6260;
    wire N__6259;
    wire N__6256;
    wire N__6251;
    wire N__6246;
    wire N__6243;
    wire N__6240;
    wire N__6239;
    wire N__6238;
    wire N__6235;
    wire N__6232;
    wire N__6229;
    wire N__6228;
    wire N__6227;
    wire N__6226;
    wire N__6219;
    wire N__6216;
    wire N__6213;
    wire N__6210;
    wire N__6201;
    wire N__6200;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6186;
    wire N__6185;
    wire N__6182;
    wire N__6179;
    wire N__6178;
    wire N__6177;
    wire N__6174;
    wire N__6171;
    wire N__6168;
    wire N__6165;
    wire N__6164;
    wire N__6163;
    wire N__6160;
    wire N__6157;
    wire N__6154;
    wire N__6151;
    wire N__6148;
    wire N__6147;
    wire N__6146;
    wire N__6145;
    wire N__6144;
    wire N__6141;
    wire N__6136;
    wire N__6129;
    wire N__6126;
    wire N__6123;
    wire N__6120;
    wire N__6117;
    wire N__6102;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6094;
    wire N__6093;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6082;
    wire N__6081;
    wire N__6080;
    wire N__6077;
    wire N__6076;
    wire N__6075;
    wire N__6072;
    wire N__6069;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6047;
    wire N__6030;
    wire N__6029;
    wire N__6028;
    wire N__6023;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6006;
    wire N__6003;
    wire N__6002;
    wire N__5999;
    wire N__5996;
    wire N__5993;
    wire N__5992;
    wire N__5991;
    wire N__5990;
    wire N__5989;
    wire N__5988;
    wire N__5985;
    wire N__5982;
    wire N__5979;
    wire N__5974;
    wire N__5969;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5943;
    wire N__5940;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5922;
    wire N__5919;
    wire N__5916;
    wire N__5913;
    wire N__5910;
    wire N__5907;
    wire N__5904;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5868;
    wire N__5865;
    wire N__5862;
    wire N__5859;
    wire N__5856;
    wire N__5853;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5838;
    wire N__5835;
    wire N__5834;
    wire N__5833;
    wire N__5830;
    wire N__5825;
    wire N__5820;
    wire N__5817;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5792;
    wire N__5791;
    wire N__5786;
    wire N__5783;
    wire N__5778;
    wire N__5777;
    wire N__5774;
    wire N__5773;
    wire N__5772;
    wire N__5769;
    wire N__5766;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5748;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5729;
    wire N__5726;
    wire N__5723;
    wire N__5718;
    wire N__5715;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5703;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5673;
    wire N__5670;
    wire N__5667;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5634;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5622;
    wire N__5619;
    wire N__5616;
    wire N__5613;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5598;
    wire N__5595;
    wire N__5592;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5568;
    wire N__5565;
    wire N__5562;
    wire N__5559;
    wire N__5558;
    wire N__5557;
    wire N__5556;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5548;
    wire N__5545;
    wire N__5540;
    wire N__5535;
    wire N__5532;
    wire N__5523;
    wire N__5522;
    wire N__5519;
    wire N__5518;
    wire N__5517;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5469;
    wire N__5466;
    wire N__5463;
    wire N__5462;
    wire N__5459;
    wire N__5456;
    wire N__5453;
    wire N__5450;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5427;
    wire N__5424;
    wire N__5421;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5400;
    wire N__5397;
    wire N__5396;
    wire N__5395;
    wire N__5394;
    wire N__5393;
    wire N__5390;
    wire N__5387;
    wire N__5386;
    wire N__5381;
    wire N__5380;
    wire N__5379;
    wire N__5378;
    wire N__5377;
    wire N__5376;
    wire N__5373;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5354;
    wire N__5349;
    wire N__5334;
    wire N__5331;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5319;
    wire N__5318;
    wire N__5317;
    wire N__5314;
    wire N__5311;
    wire N__5310;
    wire N__5307;
    wire N__5302;
    wire N__5299;
    wire N__5292;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5187;
    wire N__5184;
    wire N__5183;
    wire N__5182;
    wire N__5181;
    wire N__5180;
    wire N__5177;
    wire N__5172;
    wire N__5169;
    wire N__5166;
    wire N__5157;
    wire N__5154;
    wire N__5153;
    wire N__5152;
    wire N__5149;
    wire N__5146;
    wire N__5145;
    wire N__5142;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5130;
    wire N__5121;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5091;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5079;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5067;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5055;
    wire N__5052;
    wire N__5051;
    wire N__5050;
    wire N__5049;
    wire N__5046;
    wire N__5043;
    wire N__5042;
    wire N__5041;
    wire N__5036;
    wire N__5033;
    wire N__5026;
    wire N__5019;
    wire N__5018;
    wire N__5017;
    wire N__5010;
    wire N__5009;
    wire N__5006;
    wire N__5005;
    wire N__5002;
    wire N__4999;
    wire N__4996;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4977;
    wire N__4974;
    wire N__4973;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4904;
    wire N__4903;
    wire N__4902;
    wire N__4899;
    wire N__4898;
    wire N__4897;
    wire N__4896;
    wire N__4895;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4875;
    wire N__4872;
    wire N__4863;
    wire N__4862;
    wire N__4861;
    wire N__4858;
    wire N__4855;
    wire N__4852;
    wire N__4845;
    wire N__4842;
    wire N__4841;
    wire N__4836;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4821;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4809;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4797;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4764;
    wire N__4761;
    wire N__4758;
    wire N__4755;
    wire N__4752;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4740;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4728;
    wire N__4727;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4713;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4701;
    wire N__4698;
    wire N__4695;
    wire N__4692;
    wire N__4689;
    wire N__4686;
    wire N__4683;
    wire N__4680;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4652;
    wire N__4651;
    wire N__4650;
    wire N__4647;
    wire N__4644;
    wire N__4639;
    wire N__4632;
    wire N__4631;
    wire N__4630;
    wire N__4629;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4611;
    wire N__4608;
    wire N__4607;
    wire N__4606;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4575;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4530;
    wire N__4527;
    wire N__4524;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4494;
    wire N__4491;
    wire N__4488;
    wire N__4485;
    wire N__4482;
    wire N__4479;
    wire N__4476;
    wire N__4473;
    wire N__4470;
    wire N__4467;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4319;
    wire N__4318;
    wire N__4317;
    wire N__4316;
    wire N__4315;
    wire N__4314;
    wire N__4313;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4263;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4248;
    wire N__4245;
    wire N__4242;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4232;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4212;
    wire N__4209;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4197;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4161;
    wire N__4158;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4122;
    wire N__4119;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4107;
    wire N__4104;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4089;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4074;
    wire N__4071;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_PLL_i_i;
    wire DBRn_c_i_cascade_;
    wire DBRn_c_i_0;
    wire DBRn_c_i;
    wire \INVU712_CHIP_RAM.DMA_A20C_net ;
    wire U712_CYCLE_TERM_TCIn_0_i;
    wire \U712_CYCLE_TERM.RAM_CYCLEZ0 ;
    wire \U712_REG_SM.N_486_cascade_ ;
    wire \U712_CHIP_RAM.CLK_EN_6_0_a3_0_a2_1 ;
    wire N_490;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0 ;
    wire \U712_CHIP_RAM.N_554_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_a2_0_cascade_ ;
    wire \U712_CHIP_RAM.N_373 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0 ;
    wire \U712_CHIP_RAM.N_409 ;
    wire \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_2_cascade_ ;
    wire \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1 ;
    wire \U712_CYCLE_TERM.N_565 ;
    wire \U712_CYCLE_TERM.N_407 ;
    wire \U712_CYCLE_TERM.N_534 ;
    wire bfn_9_9_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.N_371_cascade_ ;
    wire \U712_CHIP_RAM.N_375_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_498 ;
    wire \U712_CHIP_RAM.N_547_cascade_ ;
    wire \U712_CHIP_RAM.N_501_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_a2_0_cascade_ ;
    wire bfn_9_12_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.N_666_cascade_ ;
    wire \U712_CHIP_RAM.N_393_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0 ;
    wire \U712_CHIP_RAM.CLK_EN_6_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0_cascade_ ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0 ;
    wire \U712_CHIP_RAM.N_504 ;
    wire \U712_CYCLE_TERM.N_539_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire CPU_TACKm;
    wire \U712_CYCLE_TERM.TACK_STATEZ1Z_2 ;
    wire A_c_6;
    wire A_c_13;
    wire A_c_18;
    wire A_c_16;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_ ;
    wire A_c_5;
    wire A_c_12;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire A_c_14;
    wire A_c_7;
    wire \U712_CHIP_RAM.REFRESH5lto2 ;
    wire \U712_CHIP_RAM.REFRESH5lto1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire A_c_8;
    wire A_c_15;
    wire \U712_CHIP_RAM.N_669_cascade_ ;
    wire \U712_CHIP_RAM.N_520_cascade_ ;
    wire \U712_CHIP_RAM.N_560 ;
    wire \U712_CHIP_RAM.N_501 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1 ;
    wire \U712_CHIP_RAM.N_515 ;
    wire \U712_CHIP_RAM.N_516 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.N_519 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0 ;
    wire CONSTANT_ONE_NET;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_0 ;
    wire \U712_CHIP_RAM.N_78 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.N_559_cascade_ ;
    wire \U712_CHIP_RAM.N_665 ;
    wire \U712_CHIP_RAM.N_665_cascade_ ;
    wire \U712_CHIP_RAM.N_471 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ;
    wire A_c_20;
    wire \U712_CHIP_RAM.N_506_cascade_ ;
    wire \U712_CHIP_RAM.DMA_AZ0Z20 ;
    wire \U712_CHIP_RAM.N_375 ;
    wire \U712_CHIP_RAM.N_547 ;
    wire \U712_CHIP_RAM.N_522 ;
    wire \U712_CHIP_RAM.N_523_cascade_ ;
    wire \U712_CHIP_RAM.BANK0_9 ;
    wire BANK0_c;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.N_545_cascade_ ;
    wire \U712_CHIP_RAM.N_549 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_1 ;
    wire \U712_CHIP_RAM.N_666 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_557 ;
    wire \U712_CHIP_RAM.N_393 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_0_a2_0 ;
    wire \U712_CHIP_RAM.N_557_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_ ;
    wire \U712_CHIP_RAM.N_31 ;
    wire LATCH_CLK_c;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_566 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire TACK_OUTn;
    wire ASn_c;
    wire REG_TACK;
    wire AWEn_c;
    wire \U712_CHIP_RAM.BANK0_0_sqmuxa_1 ;
    wire DBDIR_c;
    wire \U712_REG_SM.N_447 ;
    wire \U712_REG_SM.N_447_cascade_ ;
    wire \U712_REG_SM.REG_TACK_RNOZ0Z_0 ;
    wire \U712_REG_SM.N_478 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire \U712_CHIP_RAM.N_379_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.REFRESH_RST_cascade_ ;
    wire \U712_CHIP_RAM.un1_CMA28_0_i ;
    wire A_c_11;
    wire A_c_4;
    wire \U712_CHIP_RAM.N_517 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_a2_1_0 ;
    wire A_c_9;
    wire A_c_2;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CHIP_RAM.N_567 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_1_cascade_ ;
    wire \U712_CHIP_RAM.N_562 ;
    wire \U712_CHIP_RAM.N_502 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.N_545 ;
    wire \U712_CHIP_RAM.N_572 ;
    wire \U712_CHIP_RAM.N_518_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_a2_0_0 ;
    wire RAMENn_c;
    wire \U712_CHIP_RAM.N_492_cascade_ ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.STATE_COUNT_srsts_i_0_0_a2_0_0_0_cascade_ ;
    wire \U712_REG_SM.N_374 ;
    wire \U712_REG_SM.N_374_cascade_ ;
    wire \U712_REG_SM.N_417 ;
    wire C3_c;
    wire \U712_REG_SM.DS_EN_RNOZ0Z_0 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire RASn_c;
    wire WEn_c;
    wire CRCSn_c;
    wire A_c_19;
    wire CMA_c_9;
    wire A_c_17;
    wire CMA_c_8;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CMA_c_10;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire \U712_CHIP_RAM.CMA_5_i_0_8 ;
    wire TSn_c;
    wire \U712_REG_SM.N_477_cascade_ ;
    wire REGSPACEn_c;
    wire A_c_10;
    wire \U712_CHIP_RAM.N_422 ;
    wire A_c_3;
    wire \U712_CHIP_RAM.N_445 ;
    wire DBRn_c;
    wire DBR_SYNCZ0Z_0;
    wire \U712_REG_SM.START_RSTZ0 ;
    wire \U712_CYCLE_TERM.TACK_EN_RNOZ0Z_0 ;
    wire \U712_CYCLE_TERM.un13_0 ;
    wire TACK_EN;
    wire \U712_REG_SM.N_661 ;
    wire \U712_REG_SM.N_389 ;
    wire \U712_REG_SM.N_475_cascade_ ;
    wire N_57_i;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_0 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_REG_SM.N_449_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.START_RST_0_sqmuxa ;
    wire \U712_REG_SM.N_396_cascade_ ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.un1_STATE_COUNT_4_i_i_0_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_2 ;
    wire \U712_REG_SM.N_479 ;
    wire CLK40_PLL_i;
    wire CLK40_PLL_i_i;
    wire RESETn_c_i;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire \U712_CHIP_RAM.un3_DMA_CYCLE_START ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire RESETn_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire N_295_i;
    wire N_299_i;
    wire DBENn_c;
    wire DMA_CYCLEm;
    wire N_297_i;
    wire \U712_BYTE_ENABLE.N_528 ;
    wire \U712_BYTE_ENABLE.N_377_cascade_ ;
    wire \U712_BYTE_ENABLE.N_508 ;
    wire \U712_BYTE_ENABLE.N_377 ;
    wire \U712_BYTE_ENABLE.N_530 ;
    wire \U712_BYTE_ENABLE.N_532 ;
    wire \U712_BYTE_ENABLE.N_364_i ;
    wire DMA_LATCH_EN_c;
    wire N_403_i;
    wire CASn_c;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ;
    wire \U712_CHIP_RAM.N_379 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire CLK80_PLL;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire CPU_CYCLEm;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ1Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire DRA_c_1;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire N_402_i;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire DRA_c_5;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire N_291;
    wire N_400_i;
    wire DS_ENm;
    wire N_293;
    wire SIZ_c_0;
    wire A_c_1;
    wire A_c_0;
    wire SIZ_c_1;
    wire N_401_i;
    wire DRA_c_8;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire AGNUS_REV_c;
    wire RAS0n_c;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire REG_CYCLEm;
    wire DRDENn_c;
    wire RnW_c;
    wire CASUn_c;
    wire WRITE_CYCLEm;
    wire CASLn_c;
    wire N_450;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__4089),
            .RESETB(N__4938),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__12127),
            .DIN(N__12126),
            .DOUT(N__12125),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__12127),
            .PADOUT(N__12126),
            .PADIN(N__12125),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8718),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__12118),
            .DIN(N__12117),
            .DOUT(N__12116),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__12118),
            .PADOUT(N__12117),
            .PADIN(N__12116),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__12109),
            .DIN(N__12108),
            .DOUT(N__12107),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__12109),
            .PADOUT(N__12108),
            .PADIN(N__12107),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9240),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__12100),
            .DIN(N__12099),
            .DOUT(N__12098),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__12100),
            .PADOUT(N__12099),
            .PADIN(N__12098),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11121),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__12091),
            .DIN(N__12090),
            .DOUT(N__12089),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__12091),
            .PADOUT(N__12090),
            .PADIN(N__12089),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__12082),
            .DIN(N__12081),
            .DOUT(N__12080),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__12082),
            .PADOUT(N__12081),
            .PADIN(N__12080),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__12073),
            .DIN(N__12072),
            .DOUT(N__12071),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__12073),
            .PADOUT(N__12072),
            .PADIN(N__12071),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__12064),
            .DIN(N__12063),
            .DOUT(N__12062),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__12064),
            .PADOUT(N__12063),
            .PADIN(N__12062),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__12055),
            .DIN(N__12054),
            .DOUT(N__12053),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__12055),
            .PADOUT(N__12054),
            .PADIN(N__12053),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__12046),
            .DIN(N__12045),
            .DOUT(N__12044),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__12046),
            .PADOUT(N__12045),
            .PADIN(N__12044),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__12037),
            .DIN(N__12036),
            .DOUT(N__12035),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__12037),
            .PADOUT(N__12036),
            .PADIN(N__12035),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5616),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__12028),
            .DIN(N__12027),
            .DOUT(N__12026),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__12028),
            .PADOUT(N__12027),
            .PADIN(N__12026),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9252),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__12019),
            .DIN(N__12018),
            .DOUT(N__12017),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__12019),
            .PADOUT(N__12018),
            .PADIN(N__12017),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__12010),
            .DIN(N__12009),
            .DOUT(N__12008),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__12010),
            .PADOUT(N__12009),
            .PADIN(N__12008),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6485),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__12001),
            .DIN(N__12000),
            .DOUT(N__11999),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__12001),
            .PADOUT(N__12000),
            .PADIN(N__11999),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__11992),
            .DIN(N__11991),
            .DOUT(N__11990),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__11992),
            .PADOUT(N__11991),
            .PADIN(N__11990),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__11983),
            .DIN(N__11982),
            .DOUT(N__11981),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__11983),
            .PADOUT(N__11982),
            .PADIN(N__11981),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4200),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__11974),
            .DIN(N__11973),
            .DOUT(N__11972),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__11974),
            .PADOUT(N__11973),
            .PADIN(N__11972),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11965),
            .DIN(N__11964),
            .DOUT(N__11963),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11965),
            .PADOUT(N__11964),
            .PADIN(N__11963),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__11956),
            .DIN(N__11955),
            .DOUT(N__11954),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__11956),
            .PADOUT(N__11955),
            .PADIN(N__11954),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8841),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__11947),
            .DIN(N__11946),
            .DOUT(N__11945),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__11947),
            .PADOUT(N__11946),
            .PADIN(N__11945),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__11938),
            .DIN(N__11937),
            .DOUT(N__11936),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__11938),
            .PADOUT(N__11937),
            .PADIN(N__11936),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7332),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11929),
            .DIN(N__11928),
            .DOUT(N__11927),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11929),
            .PADOUT(N__11928),
            .PADIN(N__11927),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__11920),
            .DIN(N__11919),
            .DOUT(N__11918),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__11920),
            .PADOUT(N__11919),
            .PADIN(N__11918),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10746),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__11911),
            .DIN(N__11910),
            .DOUT(N__11909),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__11911),
            .PADOUT(N__11910),
            .PADIN(N__11909),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7425),
            .DIN0(),
            .DOUT0(N__5292),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__11902),
            .DIN(N__11901),
            .DOUT(N__11900),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__11902),
            .PADOUT(N__11901),
            .PADIN(N__11900),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11893),
            .DIN(N__11892),
            .DOUT(N__11891),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11893),
            .PADOUT(N__11892),
            .PADIN(N__11891),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__11884),
            .DIN(N__11883),
            .DOUT(N__11882),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__11884),
            .PADOUT(N__11883),
            .PADIN(N__11882),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11875),
            .DIN(N__11874),
            .DOUT(N__11873),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11875),
            .PADOUT(N__11874),
            .PADIN(N__11873),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__11866),
            .DIN(N__11865),
            .DOUT(N__11864),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__11866),
            .PADOUT(N__11865),
            .PADIN(N__11864),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__11857),
            .DIN(N__11856),
            .DOUT(N__11855),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__11857),
            .PADOUT(N__11856),
            .PADIN(N__11855),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9270),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__11848),
            .DIN(N__11847),
            .DOUT(N__11846),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__11848),
            .PADOUT(N__11847),
            .PADIN(N__11846),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11839),
            .DIN(N__11838),
            .DOUT(N__11837),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11839),
            .PADOUT(N__11838),
            .PADIN(N__11837),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11830),
            .DIN(N__11829),
            .DOUT(N__11828),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11830),
            .PADOUT(N__11829),
            .PADIN(N__11828),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11821),
            .DIN(N__11820),
            .DOUT(N__11819),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11821),
            .PADOUT(N__11820),
            .PADIN(N__11819),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuf_iopad (
            .OE(N__11812),
            .DIN(N__11811),
            .DOUT(N__11810),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TCIn_obuf_preio (
            .PADOEN(N__11812),
            .PADOUT(N__11811),
            .PADIN(N__11810),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4128),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__11803),
            .DIN(N__11802),
            .DOUT(N__11801),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__11803),
            .PADOUT(N__11802),
            .PADIN(N__11801),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__11794),
            .DIN(N__11793),
            .DOUT(N__11792),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__11794),
            .PADOUT(N__11793),
            .PADIN(N__11792),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6921),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__11785),
            .DIN(N__11784),
            .DOUT(N__11783),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__11785),
            .PADOUT(N__11784),
            .PADIN(N__11783),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5112),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__11776),
            .DIN(N__11775),
            .DOUT(N__11774),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__11776),
            .PADOUT(N__11775),
            .PADIN(N__11774),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8003),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11767),
            .DIN(N__11766),
            .DOUT(N__11765),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11767),
            .PADOUT(N__11766),
            .PADIN(N__11765),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4170),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__11758),
            .DIN(N__11757),
            .DOUT(N__11756),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__11758),
            .PADOUT(N__11757),
            .PADIN(N__11756),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__11749),
            .DIN(N__11748),
            .DOUT(N__11747),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__11749),
            .PADOUT(N__11748),
            .PADIN(N__11747),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5820),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_0_iopad (
            .OE(N__11740),
            .DIN(N__11739),
            .DOUT(N__11738),
            .PACKAGEPIN(DA[0]));
    defparam DA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_0_preio (
            .PADOEN(N__11740),
            .PADOUT(N__11739),
            .PADIN(N__11738),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6429),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11731),
            .DIN(N__11730),
            .DOUT(N__11729),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11731),
            .PADOUT(N__11730),
            .PADIN(N__11729),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8301),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11722),
            .DIN(N__11721),
            .DOUT(N__11720),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11722),
            .PADOUT(N__11721),
            .PADIN(N__11720),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11713),
            .DIN(N__11712),
            .DOUT(N__11711),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11713),
            .PADOUT(N__11712),
            .PADIN(N__11711),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11704),
            .DIN(N__11703),
            .DOUT(N__11702),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11704),
            .PADOUT(N__11703),
            .PADIN(N__11702),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__11695),
            .DIN(N__11694),
            .DOUT(N__11693),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__11695),
            .PADOUT(N__11694),
            .PADIN(N__11693),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__11686),
            .DIN(N__11685),
            .DOUT(N__11684),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__11686),
            .PADOUT(N__11685),
            .PADIN(N__11684),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7179),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11677),
            .DIN(N__11676),
            .DOUT(N__11675),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11677),
            .PADOUT(N__11676),
            .PADIN(N__11675),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11668),
            .DIN(N__11667),
            .DOUT(N__11666),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11668),
            .PADOUT(N__11667),
            .PADIN(N__11666),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8002),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__11659),
            .DIN(N__11658),
            .DOUT(N__11657),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__11659),
            .PADOUT(N__11658),
            .PADIN(N__11657),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9219),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11650),
            .DIN(N__11649),
            .DOUT(N__11648),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11650),
            .PADOUT(N__11649),
            .PADIN(N__11648),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10101),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11641),
            .DIN(N__11640),
            .DOUT(N__11639),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11641),
            .PADOUT(N__11640),
            .PADIN(N__11639),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7860),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11632),
            .DIN(N__11631),
            .DOUT(N__11630),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11632),
            .PADOUT(N__11631),
            .PADIN(N__11630),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7296),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__11623),
            .DIN(N__11622),
            .DOUT(N__11621),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__11623),
            .PADOUT(N__11622),
            .PADIN(N__11621),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5816),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11614),
            .DIN(N__11613),
            .DOUT(N__11612),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11614),
            .PADOUT(N__11613),
            .PADIN(N__11612),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__11605),
            .DIN(N__11604),
            .DOUT(N__11603),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__11605),
            .PADOUT(N__11604),
            .PADIN(N__11603),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__11596),
            .DIN(N__11595),
            .DOUT(N__11594),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__11596),
            .PADOUT(N__11595),
            .PADIN(N__11594),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8739),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__11587),
            .DIN(N__11586),
            .DOUT(N__11585),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__11587),
            .PADOUT(N__11586),
            .PADIN(N__11585),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7356),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__11578),
            .DIN(N__11577),
            .DOUT(N__11576),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__11578),
            .PADOUT(N__11577),
            .PADIN(N__11576),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5703),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__11569),
            .DIN(N__11568),
            .DOUT(N__11567),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__11569),
            .PADOUT(N__11568),
            .PADIN(N__11567),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8592),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__11560),
            .DIN(N__11559),
            .DOUT(N__11558),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__11560),
            .PADOUT(N__11559),
            .PADIN(N__11558),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__11551),
            .DIN(N__11550),
            .DOUT(N__11549),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__11551),
            .PADOUT(N__11550),
            .PADIN(N__11549),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_2_iopad (
            .OE(N__11542),
            .DIN(N__11541),
            .DOUT(N__11540),
            .PACKAGEPIN(DA[2]));
    defparam DA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_2_preio (
            .PADOEN(N__11542),
            .PADOUT(N__11541),
            .PADIN(N__11540),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5904),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11533),
            .DIN(N__11532),
            .DOUT(N__11531),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11533),
            .PADOUT(N__11532),
            .PADIN(N__11531),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11524),
            .DIN(N__11523),
            .DOUT(N__11522),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11524),
            .PADOUT(N__11523),
            .PADIN(N__11522),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__11515),
            .DIN(N__11514),
            .DOUT(N__11513),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__11515),
            .PADOUT(N__11514),
            .PADIN(N__11513),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7233),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__11506),
            .DIN(N__11505),
            .DOUT(N__11504),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__11506),
            .PADOUT(N__11505),
            .PADIN(N__11504),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9507),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__11497),
            .DIN(N__11496),
            .DOUT(N__11495),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__11497),
            .PADOUT(N__11496),
            .PADIN(N__11495),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__11488),
            .DIN(N__11487),
            .DOUT(N__11486),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__11488),
            .PADOUT(N__11487),
            .PADIN(N__11486),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8760),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__11479),
            .DIN(N__11478),
            .DOUT(N__11477),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__11479),
            .PADOUT(N__11478),
            .PADIN(N__11477),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7418),
            .DIN0(),
            .DOUT0(N__5291),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__11470),
            .DIN(N__11469),
            .DOUT(N__11468),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__11470),
            .PADOUT(N__11469),
            .PADIN(N__11468),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7158),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__11461),
            .DIN(N__11460),
            .DOUT(N__11459),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__11461),
            .PADOUT(N__11460),
            .PADIN(N__11459),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__11452),
            .DIN(N__11451),
            .DOUT(N__11450),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__11452),
            .PADOUT(N__11451),
            .PADIN(N__11450),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__11443),
            .DIN(N__11442),
            .DOUT(N__11441),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__11443),
            .PADOUT(N__11442),
            .PADIN(N__11441),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7257),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__11434),
            .DIN(N__11433),
            .DOUT(N__11432),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__11434),
            .PADOUT(N__11433),
            .PADIN(N__11432),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__11425),
            .DIN(N__11424),
            .DOUT(N__11423),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__11425),
            .PADOUT(N__11424),
            .PADIN(N__11423),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_1_iopad (
            .OE(N__11416),
            .DIN(N__11415),
            .DOUT(N__11414),
            .PACKAGEPIN(DA[1]));
    defparam DA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_1_preio (
            .PADOEN(N__11416),
            .PADOUT(N__11415),
            .PADIN(N__11414),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7587),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__11407),
            .DIN(N__11406),
            .DOUT(N__11405),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__11407),
            .PADOUT(N__11406),
            .PADIN(N__11405),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__11398),
            .DIN(N__11397),
            .DOUT(N__11396),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__11398),
            .PADOUT(N__11397),
            .PADIN(N__11396),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__11389),
            .DIN(N__11388),
            .DOUT(N__11387),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__11389),
            .PADOUT(N__11388),
            .PADIN(N__11387),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5646),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__11380),
            .DIN(N__11379),
            .DOUT(N__11378),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__11380),
            .PADOUT(N__11379),
            .PADIN(N__11378),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11109),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__11371),
            .DIN(N__11370),
            .DOUT(N__11369),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__11371),
            .PADOUT(N__11370),
            .PADIN(N__11369),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11091),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__11362),
            .DIN(N__11361),
            .DOUT(N__11360),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__11362),
            .PADOUT(N__11361),
            .PADIN(N__11360),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4443),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__11353),
            .DIN(N__11352),
            .DOUT(N__11351),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__11353),
            .PADOUT(N__11352),
            .PADIN(N__11351),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11344),
            .DIN(N__11343),
            .DOUT(N__11342),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11344),
            .PADOUT(N__11343),
            .PADIN(N__11342),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__11335),
            .DIN(N__11334),
            .DOUT(N__11333),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__11335),
            .PADOUT(N__11334),
            .PADIN(N__11333),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9060),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__11326),
            .DIN(N__11325),
            .DOUT(N__11324),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__11326),
            .PADOUT(N__11325),
            .PADIN(N__11324),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__11317),
            .DIN(N__11316),
            .DOUT(N__11315),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__11317),
            .PADOUT(N__11316),
            .PADIN(N__11315),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__11308),
            .DIN(N__11307),
            .DOUT(N__11306),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__11308),
            .PADOUT(N__11307),
            .PADIN(N__11306),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5427),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__11299),
            .DIN(N__11298),
            .DOUT(N__11297),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__11299),
            .PADOUT(N__11298),
            .PADIN(N__11297),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11043),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__11290),
            .DIN(N__11289),
            .DOUT(N__11288),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__11290),
            .PADOUT(N__11289),
            .PADIN(N__11288),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8004),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__11281),
            .DIN(N__11280),
            .DOUT(N__11279),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__11281),
            .PADOUT(N__11280),
            .PADIN(N__11279),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__2749 (
            .O(N__11262),
            .I(N__11259));
    InMux I__2748 (
            .O(N__11259),
            .I(N__11256));
    LocalMux I__2747 (
            .O(N__11256),
            .I(N__11252));
    InMux I__2746 (
            .O(N__11255),
            .I(N__11249));
    Span4Mux_v I__2745 (
            .O(N__11252),
            .I(N__11246));
    LocalMux I__2744 (
            .O(N__11249),
            .I(N__11243));
    Span4Mux_h I__2743 (
            .O(N__11246),
            .I(N__11239));
    Span4Mux_v I__2742 (
            .O(N__11243),
            .I(N__11236));
    InMux I__2741 (
            .O(N__11242),
            .I(N__11232));
    Sp12to4 I__2740 (
            .O(N__11239),
            .I(N__11226));
    Sp12to4 I__2739 (
            .O(N__11236),
            .I(N__11226));
    InMux I__2738 (
            .O(N__11235),
            .I(N__11223));
    LocalMux I__2737 (
            .O(N__11232),
            .I(N__11220));
    InMux I__2736 (
            .O(N__11231),
            .I(N__11217));
    Span12Mux_h I__2735 (
            .O(N__11226),
            .I(N__11210));
    LocalMux I__2734 (
            .O(N__11223),
            .I(N__11207));
    Span4Mux_h I__2733 (
            .O(N__11220),
            .I(N__11202));
    LocalMux I__2732 (
            .O(N__11217),
            .I(N__11202));
    InMux I__2731 (
            .O(N__11216),
            .I(N__11199));
    InMux I__2730 (
            .O(N__11215),
            .I(N__11196));
    InMux I__2729 (
            .O(N__11214),
            .I(N__11191));
    InMux I__2728 (
            .O(N__11213),
            .I(N__11191));
    Odrv12 I__2727 (
            .O(N__11210),
            .I(WRITE_CYCLEm));
    Odrv4 I__2726 (
            .O(N__11207),
            .I(WRITE_CYCLEm));
    Odrv4 I__2725 (
            .O(N__11202),
            .I(WRITE_CYCLEm));
    LocalMux I__2724 (
            .O(N__11199),
            .I(WRITE_CYCLEm));
    LocalMux I__2723 (
            .O(N__11196),
            .I(WRITE_CYCLEm));
    LocalMux I__2722 (
            .O(N__11191),
            .I(WRITE_CYCLEm));
    InMux I__2721 (
            .O(N__11178),
            .I(N__11175));
    LocalMux I__2720 (
            .O(N__11175),
            .I(N__11171));
    InMux I__2719 (
            .O(N__11174),
            .I(N__11166));
    Span4Mux_h I__2718 (
            .O(N__11171),
            .I(N__11163));
    InMux I__2717 (
            .O(N__11170),
            .I(N__11160));
    InMux I__2716 (
            .O(N__11169),
            .I(N__11157));
    LocalMux I__2715 (
            .O(N__11166),
            .I(N__11152));
    Span4Mux_v I__2714 (
            .O(N__11163),
            .I(N__11149));
    LocalMux I__2713 (
            .O(N__11160),
            .I(N__11144));
    LocalMux I__2712 (
            .O(N__11157),
            .I(N__11144));
    InMux I__2711 (
            .O(N__11156),
            .I(N__11139));
    InMux I__2710 (
            .O(N__11155),
            .I(N__11139));
    Span12Mux_v I__2709 (
            .O(N__11152),
            .I(N__11134));
    Sp12to4 I__2708 (
            .O(N__11149),
            .I(N__11134));
    Span12Mux_h I__2707 (
            .O(N__11144),
            .I(N__11129));
    LocalMux I__2706 (
            .O(N__11139),
            .I(N__11129));
    Span12Mux_h I__2705 (
            .O(N__11134),
            .I(N__11124));
    Span12Mux_v I__2704 (
            .O(N__11129),
            .I(N__11124));
    Odrv12 I__2703 (
            .O(N__11124),
            .I(CASLn_c));
    IoInMux I__2702 (
            .O(N__11121),
            .I(N__11118));
    LocalMux I__2701 (
            .O(N__11118),
            .I(N__11115));
    Span12Mux_s4_h I__2700 (
            .O(N__11115),
            .I(N__11112));
    Odrv12 I__2699 (
            .O(N__11112),
            .I(N_450));
    IoInMux I__2698 (
            .O(N__11109),
            .I(N__11106));
    LocalMux I__2697 (
            .O(N__11106),
            .I(N__11103));
    Span4Mux_s3_v I__2696 (
            .O(N__11103),
            .I(N__11100));
    Span4Mux_h I__2695 (
            .O(N__11100),
            .I(N__11097));
    Span4Mux_v I__2694 (
            .O(N__11097),
            .I(N__11094));
    Odrv4 I__2693 (
            .O(N__11094),
            .I(N_291));
    IoInMux I__2692 (
            .O(N__11091),
            .I(N__11088));
    LocalMux I__2691 (
            .O(N__11088),
            .I(N__11085));
    IoSpan4Mux I__2690 (
            .O(N__11085),
            .I(N__11082));
    Span4Mux_s2_v I__2689 (
            .O(N__11082),
            .I(N__11079));
    Span4Mux_v I__2688 (
            .O(N__11079),
            .I(N__11076));
    Odrv4 I__2687 (
            .O(N__11076),
            .I(N_400_i));
    InMux I__2686 (
            .O(N__11073),
            .I(N__11070));
    LocalMux I__2685 (
            .O(N__11070),
            .I(N__11066));
    InMux I__2684 (
            .O(N__11069),
            .I(N__11063));
    Span4Mux_v I__2683 (
            .O(N__11066),
            .I(N__11058));
    LocalMux I__2682 (
            .O(N__11063),
            .I(N__11058));
    Span4Mux_v I__2681 (
            .O(N__11058),
            .I(N__11055));
    Sp12to4 I__2680 (
            .O(N__11055),
            .I(N__11051));
    InMux I__2679 (
            .O(N__11054),
            .I(N__11048));
    Odrv12 I__2678 (
            .O(N__11051),
            .I(DS_ENm));
    LocalMux I__2677 (
            .O(N__11048),
            .I(DS_ENm));
    IoInMux I__2676 (
            .O(N__11043),
            .I(N__11040));
    LocalMux I__2675 (
            .O(N__11040),
            .I(N__11037));
    Span4Mux_s2_v I__2674 (
            .O(N__11037),
            .I(N__11034));
    Span4Mux_h I__2673 (
            .O(N__11034),
            .I(N__11031));
    Span4Mux_v I__2672 (
            .O(N__11031),
            .I(N__11028));
    Odrv4 I__2671 (
            .O(N__11028),
            .I(N_293));
    CascadeMux I__2670 (
            .O(N__11025),
            .I(N__11020));
    CascadeMux I__2669 (
            .O(N__11024),
            .I(N__11015));
    InMux I__2668 (
            .O(N__11023),
            .I(N__11011));
    InMux I__2667 (
            .O(N__11020),
            .I(N__11004));
    InMux I__2666 (
            .O(N__11019),
            .I(N__11004));
    InMux I__2665 (
            .O(N__11018),
            .I(N__11004));
    InMux I__2664 (
            .O(N__11015),
            .I(N__11001));
    CascadeMux I__2663 (
            .O(N__11014),
            .I(N__10998));
    LocalMux I__2662 (
            .O(N__11011),
            .I(N__10995));
    LocalMux I__2661 (
            .O(N__11004),
            .I(N__10990));
    LocalMux I__2660 (
            .O(N__11001),
            .I(N__10990));
    InMux I__2659 (
            .O(N__10998),
            .I(N__10987));
    Span4Mux_v I__2658 (
            .O(N__10995),
            .I(N__10979));
    Span4Mux_h I__2657 (
            .O(N__10990),
            .I(N__10979));
    LocalMux I__2656 (
            .O(N__10987),
            .I(N__10979));
    InMux I__2655 (
            .O(N__10986),
            .I(N__10976));
    Span4Mux_h I__2654 (
            .O(N__10979),
            .I(N__10973));
    LocalMux I__2653 (
            .O(N__10976),
            .I(N__10970));
    Span4Mux_v I__2652 (
            .O(N__10973),
            .I(N__10967));
    Span12Mux_v I__2651 (
            .O(N__10970),
            .I(N__10964));
    Span4Mux_h I__2650 (
            .O(N__10967),
            .I(N__10961));
    Span12Mux_h I__2649 (
            .O(N__10964),
            .I(N__10958));
    Sp12to4 I__2648 (
            .O(N__10961),
            .I(N__10955));
    Odrv12 I__2647 (
            .O(N__10958),
            .I(SIZ_c_0));
    Odrv12 I__2646 (
            .O(N__10955),
            .I(SIZ_c_0));
    InMux I__2645 (
            .O(N__10950),
            .I(N__10940));
    InMux I__2644 (
            .O(N__10949),
            .I(N__10940));
    InMux I__2643 (
            .O(N__10948),
            .I(N__10940));
    InMux I__2642 (
            .O(N__10947),
            .I(N__10937));
    LocalMux I__2641 (
            .O(N__10940),
            .I(N__10928));
    LocalMux I__2640 (
            .O(N__10937),
            .I(N__10928));
    InMux I__2639 (
            .O(N__10936),
            .I(N__10925));
    InMux I__2638 (
            .O(N__10935),
            .I(N__10922));
    InMux I__2637 (
            .O(N__10934),
            .I(N__10917));
    InMux I__2636 (
            .O(N__10933),
            .I(N__10917));
    Span4Mux_v I__2635 (
            .O(N__10928),
            .I(N__10914));
    LocalMux I__2634 (
            .O(N__10925),
            .I(N__10909));
    LocalMux I__2633 (
            .O(N__10922),
            .I(N__10909));
    LocalMux I__2632 (
            .O(N__10917),
            .I(N__10906));
    Span4Mux_v I__2631 (
            .O(N__10914),
            .I(N__10901));
    Span4Mux_v I__2630 (
            .O(N__10909),
            .I(N__10901));
    Span12Mux_s7_v I__2629 (
            .O(N__10906),
            .I(N__10898));
    Sp12to4 I__2628 (
            .O(N__10901),
            .I(N__10895));
    Span12Mux_h I__2627 (
            .O(N__10898),
            .I(N__10892));
    Span12Mux_h I__2626 (
            .O(N__10895),
            .I(N__10889));
    Odrv12 I__2625 (
            .O(N__10892),
            .I(A_c_1));
    Odrv12 I__2624 (
            .O(N__10889),
            .I(A_c_1));
    InMux I__2623 (
            .O(N__10884),
            .I(N__10878));
    InMux I__2622 (
            .O(N__10883),
            .I(N__10875));
    CascadeMux I__2621 (
            .O(N__10882),
            .I(N__10870));
    CascadeMux I__2620 (
            .O(N__10881),
            .I(N__10866));
    LocalMux I__2619 (
            .O(N__10878),
            .I(N__10859));
    LocalMux I__2618 (
            .O(N__10875),
            .I(N__10859));
    InMux I__2617 (
            .O(N__10874),
            .I(N__10854));
    InMux I__2616 (
            .O(N__10873),
            .I(N__10854));
    InMux I__2615 (
            .O(N__10870),
            .I(N__10851));
    InMux I__2614 (
            .O(N__10869),
            .I(N__10844));
    InMux I__2613 (
            .O(N__10866),
            .I(N__10844));
    InMux I__2612 (
            .O(N__10865),
            .I(N__10844));
    InMux I__2611 (
            .O(N__10864),
            .I(N__10841));
    Span4Mux_v I__2610 (
            .O(N__10859),
            .I(N__10834));
    LocalMux I__2609 (
            .O(N__10854),
            .I(N__10834));
    LocalMux I__2608 (
            .O(N__10851),
            .I(N__10834));
    LocalMux I__2607 (
            .O(N__10844),
            .I(N__10829));
    LocalMux I__2606 (
            .O(N__10841),
            .I(N__10829));
    Span4Mux_v I__2605 (
            .O(N__10834),
            .I(N__10826));
    Span12Mux_s10_v I__2604 (
            .O(N__10829),
            .I(N__10821));
    Sp12to4 I__2603 (
            .O(N__10826),
            .I(N__10821));
    Span12Mux_h I__2602 (
            .O(N__10821),
            .I(N__10818));
    Odrv12 I__2601 (
            .O(N__10818),
            .I(A_c_0));
    CascadeMux I__2600 (
            .O(N__10815),
            .I(N__10812));
    InMux I__2599 (
            .O(N__10812),
            .I(N__10808));
    CascadeMux I__2598 (
            .O(N__10811),
            .I(N__10803));
    LocalMux I__2597 (
            .O(N__10808),
            .I(N__10799));
    InMux I__2596 (
            .O(N__10807),
            .I(N__10792));
    InMux I__2595 (
            .O(N__10806),
            .I(N__10792));
    InMux I__2594 (
            .O(N__10803),
            .I(N__10792));
    InMux I__2593 (
            .O(N__10802),
            .I(N__10789));
    Span4Mux_v I__2592 (
            .O(N__10799),
            .I(N__10782));
    LocalMux I__2591 (
            .O(N__10792),
            .I(N__10782));
    LocalMux I__2590 (
            .O(N__10789),
            .I(N__10782));
    Span4Mux_h I__2589 (
            .O(N__10782),
            .I(N__10776));
    InMux I__2588 (
            .O(N__10781),
            .I(N__10773));
    InMux I__2587 (
            .O(N__10780),
            .I(N__10770));
    InMux I__2586 (
            .O(N__10779),
            .I(N__10767));
    Span4Mux_v I__2585 (
            .O(N__10776),
            .I(N__10764));
    LocalMux I__2584 (
            .O(N__10773),
            .I(N__10757));
    LocalMux I__2583 (
            .O(N__10770),
            .I(N__10757));
    LocalMux I__2582 (
            .O(N__10767),
            .I(N__10757));
    Sp12to4 I__2581 (
            .O(N__10764),
            .I(N__10752));
    Span12Mux_v I__2580 (
            .O(N__10757),
            .I(N__10752));
    Span12Mux_h I__2579 (
            .O(N__10752),
            .I(N__10749));
    Odrv12 I__2578 (
            .O(N__10749),
            .I(SIZ_c_1));
    IoInMux I__2577 (
            .O(N__10746),
            .I(N__10743));
    LocalMux I__2576 (
            .O(N__10743),
            .I(N__10740));
    Odrv12 I__2575 (
            .O(N__10740),
            .I(N_401_i));
    InMux I__2574 (
            .O(N__10737),
            .I(N__10733));
    InMux I__2573 (
            .O(N__10736),
            .I(N__10730));
    LocalMux I__2572 (
            .O(N__10733),
            .I(N__10725));
    LocalMux I__2571 (
            .O(N__10730),
            .I(N__10722));
    InMux I__2570 (
            .O(N__10729),
            .I(N__10719));
    InMux I__2569 (
            .O(N__10728),
            .I(N__10716));
    Span4Mux_v I__2568 (
            .O(N__10725),
            .I(N__10713));
    Span4Mux_v I__2567 (
            .O(N__10722),
            .I(N__10710));
    LocalMux I__2566 (
            .O(N__10719),
            .I(N__10707));
    LocalMux I__2565 (
            .O(N__10716),
            .I(N__10702));
    Sp12to4 I__2564 (
            .O(N__10713),
            .I(N__10702));
    Span4Mux_h I__2563 (
            .O(N__10710),
            .I(N__10697));
    Span4Mux_v I__2562 (
            .O(N__10707),
            .I(N__10697));
    Span12Mux_h I__2561 (
            .O(N__10702),
            .I(N__10694));
    Sp12to4 I__2560 (
            .O(N__10697),
            .I(N__10691));
    Odrv12 I__2559 (
            .O(N__10694),
            .I(DRA_c_8));
    Odrv12 I__2558 (
            .O(N__10691),
            .I(DRA_c_8));
    InMux I__2557 (
            .O(N__10686),
            .I(N__10681));
    InMux I__2556 (
            .O(N__10685),
            .I(N__10677));
    InMux I__2555 (
            .O(N__10684),
            .I(N__10674));
    LocalMux I__2554 (
            .O(N__10681),
            .I(N__10671));
    InMux I__2553 (
            .O(N__10680),
            .I(N__10668));
    LocalMux I__2552 (
            .O(N__10677),
            .I(N__10663));
    LocalMux I__2551 (
            .O(N__10674),
            .I(N__10663));
    Span4Mux_v I__2550 (
            .O(N__10671),
            .I(N__10660));
    LocalMux I__2549 (
            .O(N__10668),
            .I(N__10657));
    Span4Mux_v I__2548 (
            .O(N__10663),
            .I(N__10654));
    Sp12to4 I__2547 (
            .O(N__10660),
            .I(N__10647));
    Span12Mux_v I__2546 (
            .O(N__10657),
            .I(N__10647));
    Sp12to4 I__2545 (
            .O(N__10654),
            .I(N__10647));
    Span12Mux_h I__2544 (
            .O(N__10647),
            .I(N__10644));
    Odrv12 I__2543 (
            .O(N__10644),
            .I(DRA_c_7));
    InMux I__2542 (
            .O(N__10641),
            .I(N__10638));
    LocalMux I__2541 (
            .O(N__10638),
            .I(N__10635));
    Span4Mux_h I__2540 (
            .O(N__10635),
            .I(N__10632));
    Odrv4 I__2539 (
            .O(N__10632),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2538 (
            .O(N__10629),
            .I(N__10625));
    CascadeMux I__2537 (
            .O(N__10628),
            .I(N__10620));
    LocalMux I__2536 (
            .O(N__10625),
            .I(N__10616));
    InMux I__2535 (
            .O(N__10624),
            .I(N__10613));
    CascadeMux I__2534 (
            .O(N__10623),
            .I(N__10604));
    InMux I__2533 (
            .O(N__10620),
            .I(N__10593));
    InMux I__2532 (
            .O(N__10619),
            .I(N__10593));
    Span4Mux_v I__2531 (
            .O(N__10616),
            .I(N__10590));
    LocalMux I__2530 (
            .O(N__10613),
            .I(N__10587));
    InMux I__2529 (
            .O(N__10612),
            .I(N__10584));
    InMux I__2528 (
            .O(N__10611),
            .I(N__10581));
    InMux I__2527 (
            .O(N__10610),
            .I(N__10578));
    InMux I__2526 (
            .O(N__10609),
            .I(N__10573));
    InMux I__2525 (
            .O(N__10608),
            .I(N__10573));
    InMux I__2524 (
            .O(N__10607),
            .I(N__10569));
    InMux I__2523 (
            .O(N__10604),
            .I(N__10564));
    InMux I__2522 (
            .O(N__10603),
            .I(N__10564));
    InMux I__2521 (
            .O(N__10602),
            .I(N__10561));
    InMux I__2520 (
            .O(N__10601),
            .I(N__10556));
    InMux I__2519 (
            .O(N__10600),
            .I(N__10556));
    InMux I__2518 (
            .O(N__10599),
            .I(N__10551));
    InMux I__2517 (
            .O(N__10598),
            .I(N__10551));
    LocalMux I__2516 (
            .O(N__10593),
            .I(N__10546));
    Span4Mux_h I__2515 (
            .O(N__10590),
            .I(N__10540));
    Span4Mux_v I__2514 (
            .O(N__10587),
            .I(N__10540));
    LocalMux I__2513 (
            .O(N__10584),
            .I(N__10537));
    LocalMux I__2512 (
            .O(N__10581),
            .I(N__10532));
    LocalMux I__2511 (
            .O(N__10578),
            .I(N__10532));
    LocalMux I__2510 (
            .O(N__10573),
            .I(N__10529));
    InMux I__2509 (
            .O(N__10572),
            .I(N__10526));
    LocalMux I__2508 (
            .O(N__10569),
            .I(N__10523));
    LocalMux I__2507 (
            .O(N__10564),
            .I(N__10518));
    LocalMux I__2506 (
            .O(N__10561),
            .I(N__10518));
    LocalMux I__2505 (
            .O(N__10556),
            .I(N__10513));
    LocalMux I__2504 (
            .O(N__10551),
            .I(N__10513));
    InMux I__2503 (
            .O(N__10550),
            .I(N__10510));
    InMux I__2502 (
            .O(N__10549),
            .I(N__10507));
    Span4Mux_v I__2501 (
            .O(N__10546),
            .I(N__10504));
    InMux I__2500 (
            .O(N__10545),
            .I(N__10501));
    Span4Mux_h I__2499 (
            .O(N__10540),
            .I(N__10488));
    Span4Mux_v I__2498 (
            .O(N__10537),
            .I(N__10488));
    Span4Mux_v I__2497 (
            .O(N__10532),
            .I(N__10488));
    Span4Mux_h I__2496 (
            .O(N__10529),
            .I(N__10488));
    LocalMux I__2495 (
            .O(N__10526),
            .I(N__10488));
    Span4Mux_v I__2494 (
            .O(N__10523),
            .I(N__10488));
    Sp12to4 I__2493 (
            .O(N__10518),
            .I(N__10483));
    Sp12to4 I__2492 (
            .O(N__10513),
            .I(N__10483));
    LocalMux I__2491 (
            .O(N__10510),
            .I(N__10478));
    LocalMux I__2490 (
            .O(N__10507),
            .I(N__10478));
    Sp12to4 I__2489 (
            .O(N__10504),
            .I(N__10471));
    LocalMux I__2488 (
            .O(N__10501),
            .I(N__10471));
    Sp12to4 I__2487 (
            .O(N__10488),
            .I(N__10471));
    Span12Mux_v I__2486 (
            .O(N__10483),
            .I(N__10468));
    Span12Mux_h I__2485 (
            .O(N__10478),
            .I(N__10465));
    Span12Mux_h I__2484 (
            .O(N__10471),
            .I(N__10462));
    Span12Mux_h I__2483 (
            .O(N__10468),
            .I(N__10457));
    Span12Mux_v I__2482 (
            .O(N__10465),
            .I(N__10457));
    Span12Mux_v I__2481 (
            .O(N__10462),
            .I(N__10454));
    Odrv12 I__2480 (
            .O(N__10457),
            .I(AGNUS_REV_c));
    Odrv12 I__2479 (
            .O(N__10454),
            .I(AGNUS_REV_c));
    InMux I__2478 (
            .O(N__10449),
            .I(N__10446));
    LocalMux I__2477 (
            .O(N__10446),
            .I(N__10443));
    Span4Mux_v I__2476 (
            .O(N__10443),
            .I(N__10440));
    Sp12to4 I__2475 (
            .O(N__10440),
            .I(N__10437));
    Odrv12 I__2474 (
            .O(N__10437),
            .I(RAS0n_c));
    InMux I__2473 (
            .O(N__10434),
            .I(N__10430));
    InMux I__2472 (
            .O(N__10433),
            .I(N__10426));
    LocalMux I__2471 (
            .O(N__10430),
            .I(N__10423));
    InMux I__2470 (
            .O(N__10429),
            .I(N__10420));
    LocalMux I__2469 (
            .O(N__10426),
            .I(N__10417));
    Span4Mux_v I__2468 (
            .O(N__10423),
            .I(N__10411));
    LocalMux I__2467 (
            .O(N__10420),
            .I(N__10411));
    Span4Mux_v I__2466 (
            .O(N__10417),
            .I(N__10408));
    InMux I__2465 (
            .O(N__10416),
            .I(N__10405));
    Span4Mux_v I__2464 (
            .O(N__10411),
            .I(N__10402));
    Span4Mux_v I__2463 (
            .O(N__10408),
            .I(N__10399));
    LocalMux I__2462 (
            .O(N__10405),
            .I(N__10396));
    Sp12to4 I__2461 (
            .O(N__10402),
            .I(N__10391));
    Sp12to4 I__2460 (
            .O(N__10399),
            .I(N__10391));
    Span12Mux_h I__2459 (
            .O(N__10396),
            .I(N__10388));
    Span12Mux_h I__2458 (
            .O(N__10391),
            .I(N__10385));
    Span12Mux_v I__2457 (
            .O(N__10388),
            .I(N__10382));
    Span12Mux_v I__2456 (
            .O(N__10385),
            .I(N__10379));
    Odrv12 I__2455 (
            .O(N__10382),
            .I(DRA_c_9));
    Odrv12 I__2454 (
            .O(N__10379),
            .I(DRA_c_9));
    InMux I__2453 (
            .O(N__10374),
            .I(N__10371));
    LocalMux I__2452 (
            .O(N__10371),
            .I(N__10368));
    Odrv12 I__2451 (
            .O(N__10368),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    ClkMux I__2450 (
            .O(N__10365),
            .I(N__10344));
    ClkMux I__2449 (
            .O(N__10364),
            .I(N__10344));
    ClkMux I__2448 (
            .O(N__10363),
            .I(N__10344));
    ClkMux I__2447 (
            .O(N__10362),
            .I(N__10344));
    ClkMux I__2446 (
            .O(N__10361),
            .I(N__10344));
    ClkMux I__2445 (
            .O(N__10360),
            .I(N__10344));
    ClkMux I__2444 (
            .O(N__10359),
            .I(N__10344));
    GlobalMux I__2443 (
            .O(N__10344),
            .I(N__10341));
    gio2CtrlBuf I__2442 (
            .O(N__10341),
            .I(C3_c_g));
    CEMux I__2441 (
            .O(N__10338),
            .I(N__10299));
    CEMux I__2440 (
            .O(N__10337),
            .I(N__10299));
    CEMux I__2439 (
            .O(N__10336),
            .I(N__10299));
    CEMux I__2438 (
            .O(N__10335),
            .I(N__10299));
    CEMux I__2437 (
            .O(N__10334),
            .I(N__10299));
    CEMux I__2436 (
            .O(N__10333),
            .I(N__10299));
    CEMux I__2435 (
            .O(N__10332),
            .I(N__10299));
    CEMux I__2434 (
            .O(N__10331),
            .I(N__10299));
    CEMux I__2433 (
            .O(N__10330),
            .I(N__10299));
    CEMux I__2432 (
            .O(N__10329),
            .I(N__10299));
    CEMux I__2431 (
            .O(N__10328),
            .I(N__10299));
    CEMux I__2430 (
            .O(N__10327),
            .I(N__10299));
    CEMux I__2429 (
            .O(N__10326),
            .I(N__10299));
    GlobalMux I__2428 (
            .O(N__10299),
            .I(N__10296));
    gio2CtrlBuf I__2427 (
            .O(N__10296),
            .I(DBRn_c_i_0_g));
    InMux I__2426 (
            .O(N__10293),
            .I(N__10286));
    InMux I__2425 (
            .O(N__10292),
            .I(N__10283));
    InMux I__2424 (
            .O(N__10291),
            .I(N__10280));
    InMux I__2423 (
            .O(N__10290),
            .I(N__10277));
    InMux I__2422 (
            .O(N__10289),
            .I(N__10274));
    LocalMux I__2421 (
            .O(N__10286),
            .I(N__10265));
    LocalMux I__2420 (
            .O(N__10283),
            .I(N__10262));
    LocalMux I__2419 (
            .O(N__10280),
            .I(N__10250));
    LocalMux I__2418 (
            .O(N__10277),
            .I(N__10240));
    LocalMux I__2417 (
            .O(N__10274),
            .I(N__10233));
    SRMux I__2416 (
            .O(N__10273),
            .I(N__10146));
    SRMux I__2415 (
            .O(N__10272),
            .I(N__10146));
    SRMux I__2414 (
            .O(N__10271),
            .I(N__10146));
    SRMux I__2413 (
            .O(N__10270),
            .I(N__10146));
    SRMux I__2412 (
            .O(N__10269),
            .I(N__10146));
    SRMux I__2411 (
            .O(N__10268),
            .I(N__10146));
    Glb2LocalMux I__2410 (
            .O(N__10265),
            .I(N__10146));
    Glb2LocalMux I__2409 (
            .O(N__10262),
            .I(N__10146));
    SRMux I__2408 (
            .O(N__10261),
            .I(N__10146));
    SRMux I__2407 (
            .O(N__10260),
            .I(N__10146));
    SRMux I__2406 (
            .O(N__10259),
            .I(N__10146));
    SRMux I__2405 (
            .O(N__10258),
            .I(N__10146));
    SRMux I__2404 (
            .O(N__10257),
            .I(N__10146));
    SRMux I__2403 (
            .O(N__10256),
            .I(N__10146));
    SRMux I__2402 (
            .O(N__10255),
            .I(N__10146));
    SRMux I__2401 (
            .O(N__10254),
            .I(N__10146));
    SRMux I__2400 (
            .O(N__10253),
            .I(N__10146));
    Glb2LocalMux I__2399 (
            .O(N__10250),
            .I(N__10146));
    SRMux I__2398 (
            .O(N__10249),
            .I(N__10146));
    SRMux I__2397 (
            .O(N__10248),
            .I(N__10146));
    SRMux I__2396 (
            .O(N__10247),
            .I(N__10146));
    SRMux I__2395 (
            .O(N__10246),
            .I(N__10146));
    SRMux I__2394 (
            .O(N__10245),
            .I(N__10146));
    SRMux I__2393 (
            .O(N__10244),
            .I(N__10146));
    SRMux I__2392 (
            .O(N__10243),
            .I(N__10146));
    Glb2LocalMux I__2391 (
            .O(N__10240),
            .I(N__10146));
    SRMux I__2390 (
            .O(N__10239),
            .I(N__10146));
    SRMux I__2389 (
            .O(N__10238),
            .I(N__10146));
    SRMux I__2388 (
            .O(N__10237),
            .I(N__10146));
    SRMux I__2387 (
            .O(N__10236),
            .I(N__10146));
    Glb2LocalMux I__2386 (
            .O(N__10233),
            .I(N__10146));
    SRMux I__2385 (
            .O(N__10232),
            .I(N__10146));
    SRMux I__2384 (
            .O(N__10231),
            .I(N__10146));
    SRMux I__2383 (
            .O(N__10230),
            .I(N__10146));
    SRMux I__2382 (
            .O(N__10229),
            .I(N__10146));
    SRMux I__2381 (
            .O(N__10228),
            .I(N__10146));
    SRMux I__2380 (
            .O(N__10227),
            .I(N__10146));
    SRMux I__2379 (
            .O(N__10226),
            .I(N__10146));
    SRMux I__2378 (
            .O(N__10225),
            .I(N__10146));
    GlobalMux I__2377 (
            .O(N__10146),
            .I(N__10143));
    gio2CtrlBuf I__2376 (
            .O(N__10143),
            .I(RESETn_c_i_g));
    InMux I__2375 (
            .O(N__10140),
            .I(N__10137));
    LocalMux I__2374 (
            .O(N__10137),
            .I(N__10134));
    Span4Mux_v I__2373 (
            .O(N__10134),
            .I(N__10131));
    Span4Mux_h I__2372 (
            .O(N__10131),
            .I(N__10127));
    InMux I__2371 (
            .O(N__10130),
            .I(N__10124));
    Sp12to4 I__2370 (
            .O(N__10127),
            .I(N__10121));
    LocalMux I__2369 (
            .O(N__10124),
            .I(N__10118));
    Span12Mux_h I__2368 (
            .O(N__10121),
            .I(N__10114));
    Span4Mux_v I__2367 (
            .O(N__10118),
            .I(N__10111));
    InMux I__2366 (
            .O(N__10117),
            .I(N__10108));
    Odrv12 I__2365 (
            .O(N__10114),
            .I(REG_CYCLEm));
    Odrv4 I__2364 (
            .O(N__10111),
            .I(REG_CYCLEm));
    LocalMux I__2363 (
            .O(N__10108),
            .I(REG_CYCLEm));
    IoInMux I__2362 (
            .O(N__10101),
            .I(N__10098));
    LocalMux I__2361 (
            .O(N__10098),
            .I(N__10095));
    Span4Mux_s2_v I__2360 (
            .O(N__10095),
            .I(N__10092));
    Span4Mux_v I__2359 (
            .O(N__10092),
            .I(N__10089));
    Odrv4 I__2358 (
            .O(N__10089),
            .I(DRDENn_c));
    InMux I__2357 (
            .O(N__10086),
            .I(N__10083));
    LocalMux I__2356 (
            .O(N__10083),
            .I(N__10079));
    InMux I__2355 (
            .O(N__10082),
            .I(N__10076));
    Span4Mux_v I__2354 (
            .O(N__10079),
            .I(N__10073));
    LocalMux I__2353 (
            .O(N__10076),
            .I(N__10069));
    Span4Mux_v I__2352 (
            .O(N__10073),
            .I(N__10065));
    InMux I__2351 (
            .O(N__10072),
            .I(N__10062));
    Span4Mux_v I__2350 (
            .O(N__10069),
            .I(N__10059));
    InMux I__2349 (
            .O(N__10068),
            .I(N__10056));
    Sp12to4 I__2348 (
            .O(N__10065),
            .I(N__10053));
    LocalMux I__2347 (
            .O(N__10062),
            .I(N__10050));
    Sp12to4 I__2346 (
            .O(N__10059),
            .I(N__10045));
    LocalMux I__2345 (
            .O(N__10056),
            .I(N__10045));
    Span12Mux_h I__2344 (
            .O(N__10053),
            .I(N__10040));
    Span12Mux_v I__2343 (
            .O(N__10050),
            .I(N__10040));
    Span12Mux_h I__2342 (
            .O(N__10045),
            .I(N__10037));
    Span12Mux_h I__2341 (
            .O(N__10040),
            .I(N__10032));
    Span12Mux_v I__2340 (
            .O(N__10037),
            .I(N__10032));
    Odrv12 I__2339 (
            .O(N__10032),
            .I(RnW_c));
    InMux I__2338 (
            .O(N__10029),
            .I(N__10025));
    CascadeMux I__2337 (
            .O(N__10028),
            .I(N__10021));
    LocalMux I__2336 (
            .O(N__10025),
            .I(N__10016));
    InMux I__2335 (
            .O(N__10024),
            .I(N__10011));
    InMux I__2334 (
            .O(N__10021),
            .I(N__10011));
    InMux I__2333 (
            .O(N__10020),
            .I(N__10008));
    CascadeMux I__2332 (
            .O(N__10019),
            .I(N__10005));
    Sp12to4 I__2331 (
            .O(N__10016),
            .I(N__9997));
    LocalMux I__2330 (
            .O(N__10011),
            .I(N__9997));
    LocalMux I__2329 (
            .O(N__10008),
            .I(N__9997));
    InMux I__2328 (
            .O(N__10005),
            .I(N__9992));
    InMux I__2327 (
            .O(N__10004),
            .I(N__9992));
    Span12Mux_v I__2326 (
            .O(N__9997),
            .I(N__9989));
    LocalMux I__2325 (
            .O(N__9992),
            .I(N__9986));
    Span12Mux_h I__2324 (
            .O(N__9989),
            .I(N__9983));
    Span4Mux_v I__2323 (
            .O(N__9986),
            .I(N__9980));
    Odrv12 I__2322 (
            .O(N__9983),
            .I(CASUn_c));
    Odrv4 I__2321 (
            .O(N__9980),
            .I(CASUn_c));
    CascadeMux I__2320 (
            .O(N__9975),
            .I(N__9971));
    CascadeMux I__2319 (
            .O(N__9974),
            .I(N__9968));
    InMux I__2318 (
            .O(N__9971),
            .I(N__9954));
    InMux I__2317 (
            .O(N__9968),
            .I(N__9954));
    CascadeMux I__2316 (
            .O(N__9967),
            .I(N__9947));
    InMux I__2315 (
            .O(N__9966),
            .I(N__9942));
    InMux I__2314 (
            .O(N__9965),
            .I(N__9939));
    InMux I__2313 (
            .O(N__9964),
            .I(N__9933));
    InMux I__2312 (
            .O(N__9963),
            .I(N__9925));
    InMux I__2311 (
            .O(N__9962),
            .I(N__9925));
    InMux I__2310 (
            .O(N__9961),
            .I(N__9925));
    InMux I__2309 (
            .O(N__9960),
            .I(N__9922));
    CascadeMux I__2308 (
            .O(N__9959),
            .I(N__9919));
    LocalMux I__2307 (
            .O(N__9954),
            .I(N__9915));
    InMux I__2306 (
            .O(N__9953),
            .I(N__9908));
    InMux I__2305 (
            .O(N__9952),
            .I(N__9908));
    InMux I__2304 (
            .O(N__9951),
            .I(N__9908));
    InMux I__2303 (
            .O(N__9950),
            .I(N__9905));
    InMux I__2302 (
            .O(N__9947),
            .I(N__9902));
    InMux I__2301 (
            .O(N__9946),
            .I(N__9899));
    InMux I__2300 (
            .O(N__9945),
            .I(N__9896));
    LocalMux I__2299 (
            .O(N__9942),
            .I(N__9892));
    LocalMux I__2298 (
            .O(N__9939),
            .I(N__9889));
    InMux I__2297 (
            .O(N__9938),
            .I(N__9886));
    InMux I__2296 (
            .O(N__9937),
            .I(N__9881));
    InMux I__2295 (
            .O(N__9936),
            .I(N__9881));
    LocalMux I__2294 (
            .O(N__9933),
            .I(N__9878));
    InMux I__2293 (
            .O(N__9932),
            .I(N__9875));
    LocalMux I__2292 (
            .O(N__9925),
            .I(N__9872));
    LocalMux I__2291 (
            .O(N__9922),
            .I(N__9869));
    InMux I__2290 (
            .O(N__9919),
            .I(N__9866));
    InMux I__2289 (
            .O(N__9918),
            .I(N__9863));
    Span4Mux_v I__2288 (
            .O(N__9915),
            .I(N__9854));
    LocalMux I__2287 (
            .O(N__9908),
            .I(N__9854));
    LocalMux I__2286 (
            .O(N__9905),
            .I(N__9854));
    LocalMux I__2285 (
            .O(N__9902),
            .I(N__9854));
    LocalMux I__2284 (
            .O(N__9899),
            .I(N__9849));
    LocalMux I__2283 (
            .O(N__9896),
            .I(N__9849));
    InMux I__2282 (
            .O(N__9895),
            .I(N__9846));
    Span4Mux_h I__2281 (
            .O(N__9892),
            .I(N__9839));
    Span4Mux_v I__2280 (
            .O(N__9889),
            .I(N__9839));
    LocalMux I__2279 (
            .O(N__9886),
            .I(N__9839));
    LocalMux I__2278 (
            .O(N__9881),
            .I(N__9836));
    Span4Mux_h I__2277 (
            .O(N__9878),
            .I(N__9831));
    LocalMux I__2276 (
            .O(N__9875),
            .I(N__9831));
    Span4Mux_v I__2275 (
            .O(N__9872),
            .I(N__9822));
    Span4Mux_v I__2274 (
            .O(N__9869),
            .I(N__9822));
    LocalMux I__2273 (
            .O(N__9866),
            .I(N__9822));
    LocalMux I__2272 (
            .O(N__9863),
            .I(N__9822));
    Span4Mux_h I__2271 (
            .O(N__9854),
            .I(N__9819));
    Span12Mux_h I__2270 (
            .O(N__9849),
            .I(N__9814));
    LocalMux I__2269 (
            .O(N__9846),
            .I(N__9814));
    Span4Mux_v I__2268 (
            .O(N__9839),
            .I(N__9805));
    Span4Mux_h I__2267 (
            .O(N__9836),
            .I(N__9805));
    Span4Mux_v I__2266 (
            .O(N__9831),
            .I(N__9805));
    Span4Mux_h I__2265 (
            .O(N__9822),
            .I(N__9805));
    Odrv4 I__2264 (
            .O(N__9819),
            .I(CPU_CYCLEm));
    Odrv12 I__2263 (
            .O(N__9814),
            .I(CPU_CYCLEm));
    Odrv4 I__2262 (
            .O(N__9805),
            .I(CPU_CYCLEm));
    InMux I__2261 (
            .O(N__9798),
            .I(N__9795));
    LocalMux I__2260 (
            .O(N__9795),
            .I(N__9792));
    Odrv12 I__2259 (
            .O(N__9792),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    CascadeMux I__2258 (
            .O(N__9789),
            .I(N__9783));
    InMux I__2257 (
            .O(N__9788),
            .I(N__9776));
    CascadeMux I__2256 (
            .O(N__9787),
            .I(N__9773));
    CascadeMux I__2255 (
            .O(N__9786),
            .I(N__9770));
    InMux I__2254 (
            .O(N__9783),
            .I(N__9765));
    InMux I__2253 (
            .O(N__9782),
            .I(N__9765));
    InMux I__2252 (
            .O(N__9781),
            .I(N__9760));
    InMux I__2251 (
            .O(N__9780),
            .I(N__9760));
    CascadeMux I__2250 (
            .O(N__9779),
            .I(N__9755));
    LocalMux I__2249 (
            .O(N__9776),
            .I(N__9752));
    InMux I__2248 (
            .O(N__9773),
            .I(N__9749));
    InMux I__2247 (
            .O(N__9770),
            .I(N__9746));
    LocalMux I__2246 (
            .O(N__9765),
            .I(N__9733));
    LocalMux I__2245 (
            .O(N__9760),
            .I(N__9733));
    InMux I__2244 (
            .O(N__9759),
            .I(N__9726));
    InMux I__2243 (
            .O(N__9758),
            .I(N__9726));
    InMux I__2242 (
            .O(N__9755),
            .I(N__9726));
    Span4Mux_v I__2241 (
            .O(N__9752),
            .I(N__9721));
    LocalMux I__2240 (
            .O(N__9749),
            .I(N__9721));
    LocalMux I__2239 (
            .O(N__9746),
            .I(N__9718));
    InMux I__2238 (
            .O(N__9745),
            .I(N__9714));
    InMux I__2237 (
            .O(N__9744),
            .I(N__9711));
    InMux I__2236 (
            .O(N__9743),
            .I(N__9706));
    InMux I__2235 (
            .O(N__9742),
            .I(N__9706));
    InMux I__2234 (
            .O(N__9741),
            .I(N__9699));
    InMux I__2233 (
            .O(N__9740),
            .I(N__9699));
    InMux I__2232 (
            .O(N__9739),
            .I(N__9699));
    InMux I__2231 (
            .O(N__9738),
            .I(N__9691));
    Span4Mux_v I__2230 (
            .O(N__9733),
            .I(N__9688));
    LocalMux I__2229 (
            .O(N__9726),
            .I(N__9683));
    Span4Mux_h I__2228 (
            .O(N__9721),
            .I(N__9683));
    Span12Mux_v I__2227 (
            .O(N__9718),
            .I(N__9680));
    InMux I__2226 (
            .O(N__9717),
            .I(N__9677));
    LocalMux I__2225 (
            .O(N__9714),
            .I(N__9672));
    LocalMux I__2224 (
            .O(N__9711),
            .I(N__9672));
    LocalMux I__2223 (
            .O(N__9706),
            .I(N__9667));
    LocalMux I__2222 (
            .O(N__9699),
            .I(N__9667));
    InMux I__2221 (
            .O(N__9698),
            .I(N__9662));
    InMux I__2220 (
            .O(N__9697),
            .I(N__9662));
    InMux I__2219 (
            .O(N__9696),
            .I(N__9657));
    InMux I__2218 (
            .O(N__9695),
            .I(N__9657));
    InMux I__2217 (
            .O(N__9694),
            .I(N__9654));
    LocalMux I__2216 (
            .O(N__9691),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_1 ));
    Odrv4 I__2215 (
            .O(N__9688),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_1 ));
    Odrv4 I__2214 (
            .O(N__9683),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_1 ));
    Odrv12 I__2213 (
            .O(N__9680),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_1 ));
    LocalMux I__2212 (
            .O(N__9677),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_1 ));
    Odrv4 I__2211 (
            .O(N__9672),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_1 ));
    Odrv4 I__2210 (
            .O(N__9667),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_1 ));
    LocalMux I__2209 (
            .O(N__9662),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_1 ));
    LocalMux I__2208 (
            .O(N__9657),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_1 ));
    LocalMux I__2207 (
            .O(N__9654),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_1 ));
    InMux I__2206 (
            .O(N__9633),
            .I(N__9630));
    LocalMux I__2205 (
            .O(N__9630),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    InMux I__2204 (
            .O(N__9627),
            .I(N__9624));
    LocalMux I__2203 (
            .O(N__9624),
            .I(N__9621));
    Odrv4 I__2202 (
            .O(N__9621),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2201 (
            .O(N__9618),
            .I(N__9615));
    LocalMux I__2200 (
            .O(N__9615),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    CascadeMux I__2199 (
            .O(N__9612),
            .I(N__9609));
    InMux I__2198 (
            .O(N__9609),
            .I(N__9606));
    LocalMux I__2197 (
            .O(N__9606),
            .I(N__9603));
    Span4Mux_h I__2196 (
            .O(N__9603),
            .I(N__9600));
    Odrv4 I__2195 (
            .O(N__9600),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2194 (
            .O(N__9597),
            .I(N__9594));
    LocalMux I__2193 (
            .O(N__9594),
            .I(N__9591));
    Odrv4 I__2192 (
            .O(N__9591),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__2191 (
            .O(N__9588),
            .I(N__9583));
    InMux I__2190 (
            .O(N__9587),
            .I(N__9579));
    InMux I__2189 (
            .O(N__9586),
            .I(N__9576));
    LocalMux I__2188 (
            .O(N__9583),
            .I(N__9573));
    InMux I__2187 (
            .O(N__9582),
            .I(N__9570));
    LocalMux I__2186 (
            .O(N__9579),
            .I(N__9565));
    LocalMux I__2185 (
            .O(N__9576),
            .I(N__9565));
    Span4Mux_v I__2184 (
            .O(N__9573),
            .I(N__9560));
    LocalMux I__2183 (
            .O(N__9570),
            .I(N__9560));
    Span4Mux_h I__2182 (
            .O(N__9565),
            .I(N__9557));
    Span4Mux_h I__2181 (
            .O(N__9560),
            .I(N__9554));
    Sp12to4 I__2180 (
            .O(N__9557),
            .I(N__9549));
    Sp12to4 I__2179 (
            .O(N__9554),
            .I(N__9549));
    Span12Mux_v I__2178 (
            .O(N__9549),
            .I(N__9546));
    Odrv12 I__2177 (
            .O(N__9546),
            .I(DRA_c_1));
    InMux I__2176 (
            .O(N__9543),
            .I(N__9540));
    LocalMux I__2175 (
            .O(N__9540),
            .I(N__9536));
    InMux I__2174 (
            .O(N__9539),
            .I(N__9533));
    Span4Mux_v I__2173 (
            .O(N__9536),
            .I(N__9528));
    LocalMux I__2172 (
            .O(N__9533),
            .I(N__9528));
    Sp12to4 I__2171 (
            .O(N__9528),
            .I(N__9525));
    Span12Mux_v I__2170 (
            .O(N__9525),
            .I(N__9522));
    Span12Mux_h I__2169 (
            .O(N__9522),
            .I(N__9519));
    Odrv12 I__2168 (
            .O(N__9519),
            .I(DRA_c_0));
    InMux I__2167 (
            .O(N__9516),
            .I(N__9513));
    LocalMux I__2166 (
            .O(N__9513),
            .I(N__9510));
    Odrv12 I__2165 (
            .O(N__9510),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    IoInMux I__2164 (
            .O(N__9507),
            .I(N__9504));
    LocalMux I__2163 (
            .O(N__9504),
            .I(N__9501));
    Span4Mux_s3_v I__2162 (
            .O(N__9501),
            .I(N__9498));
    Odrv4 I__2161 (
            .O(N__9498),
            .I(N_402_i));
    InMux I__2160 (
            .O(N__9495),
            .I(N__9490));
    InMux I__2159 (
            .O(N__9494),
            .I(N__9487));
    InMux I__2158 (
            .O(N__9493),
            .I(N__9483));
    LocalMux I__2157 (
            .O(N__9490),
            .I(N__9478));
    LocalMux I__2156 (
            .O(N__9487),
            .I(N__9478));
    InMux I__2155 (
            .O(N__9486),
            .I(N__9475));
    LocalMux I__2154 (
            .O(N__9483),
            .I(N__9472));
    Span4Mux_v I__2153 (
            .O(N__9478),
            .I(N__9467));
    LocalMux I__2152 (
            .O(N__9475),
            .I(N__9467));
    Span4Mux_v I__2151 (
            .O(N__9472),
            .I(N__9464));
    Span4Mux_h I__2150 (
            .O(N__9467),
            .I(N__9461));
    Span4Mux_v I__2149 (
            .O(N__9464),
            .I(N__9458));
    Span4Mux_v I__2148 (
            .O(N__9461),
            .I(N__9455));
    Sp12to4 I__2147 (
            .O(N__9458),
            .I(N__9450));
    Sp12to4 I__2146 (
            .O(N__9455),
            .I(N__9450));
    Odrv12 I__2145 (
            .O(N__9450),
            .I(DRA_c_6));
    CascadeMux I__2144 (
            .O(N__9447),
            .I(N__9444));
    InMux I__2143 (
            .O(N__9444),
            .I(N__9441));
    LocalMux I__2142 (
            .O(N__9441),
            .I(N__9438));
    Odrv4 I__2141 (
            .O(N__9438),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2140 (
            .O(N__9435),
            .I(N__9432));
    LocalMux I__2139 (
            .O(N__9432),
            .I(N__9426));
    InMux I__2138 (
            .O(N__9431),
            .I(N__9423));
    InMux I__2137 (
            .O(N__9430),
            .I(N__9420));
    InMux I__2136 (
            .O(N__9429),
            .I(N__9417));
    Span4Mux_h I__2135 (
            .O(N__9426),
            .I(N__9410));
    LocalMux I__2134 (
            .O(N__9423),
            .I(N__9410));
    LocalMux I__2133 (
            .O(N__9420),
            .I(N__9410));
    LocalMux I__2132 (
            .O(N__9417),
            .I(N__9407));
    Span4Mux_h I__2131 (
            .O(N__9410),
            .I(N__9404));
    Span4Mux_v I__2130 (
            .O(N__9407),
            .I(N__9401));
    Sp12to4 I__2129 (
            .O(N__9404),
            .I(N__9398));
    Span4Mux_v I__2128 (
            .O(N__9401),
            .I(N__9395));
    Span12Mux_v I__2127 (
            .O(N__9398),
            .I(N__9390));
    Sp12to4 I__2126 (
            .O(N__9395),
            .I(N__9390));
    Odrv12 I__2125 (
            .O(N__9390),
            .I(DRA_c_5));
    InMux I__2124 (
            .O(N__9387),
            .I(N__9383));
    InMux I__2123 (
            .O(N__9386),
            .I(N__9379));
    LocalMux I__2122 (
            .O(N__9383),
            .I(N__9376));
    InMux I__2121 (
            .O(N__9382),
            .I(N__9373));
    LocalMux I__2120 (
            .O(N__9379),
            .I(N__9370));
    Span4Mux_v I__2119 (
            .O(N__9376),
            .I(N__9364));
    LocalMux I__2118 (
            .O(N__9373),
            .I(N__9364));
    Span4Mux_v I__2117 (
            .O(N__9370),
            .I(N__9361));
    InMux I__2116 (
            .O(N__9369),
            .I(N__9358));
    Span4Mux_h I__2115 (
            .O(N__9364),
            .I(N__9355));
    Span4Mux_v I__2114 (
            .O(N__9361),
            .I(N__9352));
    LocalMux I__2113 (
            .O(N__9358),
            .I(N__9349));
    Span4Mux_v I__2112 (
            .O(N__9355),
            .I(N__9346));
    Sp12to4 I__2111 (
            .O(N__9352),
            .I(N__9339));
    Span12Mux_v I__2110 (
            .O(N__9349),
            .I(N__9339));
    Sp12to4 I__2109 (
            .O(N__9346),
            .I(N__9339));
    Span12Mux_h I__2108 (
            .O(N__9339),
            .I(N__9336));
    Odrv12 I__2107 (
            .O(N__9336),
            .I(DRA_c_4));
    InMux I__2106 (
            .O(N__9333),
            .I(N__9330));
    LocalMux I__2105 (
            .O(N__9330),
            .I(N__9327));
    Odrv4 I__2104 (
            .O(N__9327),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    CascadeMux I__2103 (
            .O(N__9324),
            .I(N__9321));
    InMux I__2102 (
            .O(N__9321),
            .I(N__9318));
    LocalMux I__2101 (
            .O(N__9318),
            .I(\U712_BYTE_ENABLE.N_377 ));
    InMux I__2100 (
            .O(N__9315),
            .I(N__9312));
    LocalMux I__2099 (
            .O(N__9312),
            .I(\U712_BYTE_ENABLE.N_530 ));
    InMux I__2098 (
            .O(N__9309),
            .I(N__9306));
    LocalMux I__2097 (
            .O(N__9306),
            .I(N__9303));
    Odrv4 I__2096 (
            .O(N__9303),
            .I(\U712_BYTE_ENABLE.N_532 ));
    CascadeMux I__2095 (
            .O(N__9300),
            .I(N__9297));
    InMux I__2094 (
            .O(N__9297),
            .I(N__9291));
    InMux I__2093 (
            .O(N__9296),
            .I(N__9286));
    InMux I__2092 (
            .O(N__9295),
            .I(N__9286));
    InMux I__2091 (
            .O(N__9294),
            .I(N__9283));
    LocalMux I__2090 (
            .O(N__9291),
            .I(N__9278));
    LocalMux I__2089 (
            .O(N__9286),
            .I(N__9278));
    LocalMux I__2088 (
            .O(N__9283),
            .I(N__9275));
    Odrv12 I__2087 (
            .O(N__9278),
            .I(\U712_BYTE_ENABLE.N_364_i ));
    Odrv4 I__2086 (
            .O(N__9275),
            .I(\U712_BYTE_ENABLE.N_364_i ));
    IoInMux I__2085 (
            .O(N__9270),
            .I(N__9267));
    LocalMux I__2084 (
            .O(N__9267),
            .I(N__9264));
    Span4Mux_s1_v I__2083 (
            .O(N__9264),
            .I(N__9261));
    Sp12to4 I__2082 (
            .O(N__9261),
            .I(N__9258));
    Span12Mux_h I__2081 (
            .O(N__9258),
            .I(N__9255));
    Odrv12 I__2080 (
            .O(N__9255),
            .I(DMA_LATCH_EN_c));
    IoInMux I__2079 (
            .O(N__9252),
            .I(N__9249));
    LocalMux I__2078 (
            .O(N__9249),
            .I(N__9246));
    Span4Mux_s3_v I__2077 (
            .O(N__9246),
            .I(N__9243));
    Odrv4 I__2076 (
            .O(N__9243),
            .I(N_403_i));
    IoInMux I__2075 (
            .O(N__9240),
            .I(N__9237));
    LocalMux I__2074 (
            .O(N__9237),
            .I(N__9234));
    Span4Mux_s1_v I__2073 (
            .O(N__9234),
            .I(N__9231));
    Span4Mux_v I__2072 (
            .O(N__9231),
            .I(N__9228));
    Span4Mux_v I__2071 (
            .O(N__9228),
            .I(N__9225));
    Sp12to4 I__2070 (
            .O(N__9225),
            .I(N__9222));
    Odrv12 I__2069 (
            .O(N__9222),
            .I(CASn_c));
    IoInMux I__2068 (
            .O(N__9219),
            .I(N__9216));
    LocalMux I__2067 (
            .O(N__9216),
            .I(N__9213));
    IoSpan4Mux I__2066 (
            .O(N__9213),
            .I(N__9210));
    Span4Mux_s3_v I__2065 (
            .O(N__9210),
            .I(N__9207));
    Span4Mux_v I__2064 (
            .O(N__9207),
            .I(N__9204));
    Sp12to4 I__2063 (
            .O(N__9204),
            .I(N__9201));
    Span12Mux_h I__2062 (
            .O(N__9201),
            .I(N__9198));
    Odrv12 I__2061 (
            .O(N__9198),
            .I(CMA_c_4));
    CascadeMux I__2060 (
            .O(N__9195),
            .I(N__9188));
    CascadeMux I__2059 (
            .O(N__9194),
            .I(N__9185));
    CascadeMux I__2058 (
            .O(N__9193),
            .I(N__9182));
    CascadeMux I__2057 (
            .O(N__9192),
            .I(N__9179));
    InMux I__2056 (
            .O(N__9191),
            .I(N__9174));
    InMux I__2055 (
            .O(N__9188),
            .I(N__9174));
    InMux I__2054 (
            .O(N__9185),
            .I(N__9170));
    InMux I__2053 (
            .O(N__9182),
            .I(N__9167));
    InMux I__2052 (
            .O(N__9179),
            .I(N__9164));
    LocalMux I__2051 (
            .O(N__9174),
            .I(N__9161));
    CascadeMux I__2050 (
            .O(N__9173),
            .I(N__9158));
    LocalMux I__2049 (
            .O(N__9170),
            .I(N__9155));
    LocalMux I__2048 (
            .O(N__9167),
            .I(N__9148));
    LocalMux I__2047 (
            .O(N__9164),
            .I(N__9148));
    Span4Mux_h I__2046 (
            .O(N__9161),
            .I(N__9148));
    InMux I__2045 (
            .O(N__9158),
            .I(N__9145));
    Span4Mux_h I__2044 (
            .O(N__9155),
            .I(N__9142));
    Span4Mux_v I__2043 (
            .O(N__9148),
            .I(N__9139));
    LocalMux I__2042 (
            .O(N__9145),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    Odrv4 I__2041 (
            .O(N__9142),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    Odrv4 I__2040 (
            .O(N__9139),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    InMux I__2039 (
            .O(N__9132),
            .I(N__9128));
    CascadeMux I__2038 (
            .O(N__9131),
            .I(N__9122));
    LocalMux I__2037 (
            .O(N__9128),
            .I(N__9118));
    InMux I__2036 (
            .O(N__9127),
            .I(N__9113));
    InMux I__2035 (
            .O(N__9126),
            .I(N__9113));
    InMux I__2034 (
            .O(N__9125),
            .I(N__9109));
    InMux I__2033 (
            .O(N__9122),
            .I(N__9104));
    InMux I__2032 (
            .O(N__9121),
            .I(N__9104));
    Span4Mux_v I__2031 (
            .O(N__9118),
            .I(N__9099));
    LocalMux I__2030 (
            .O(N__9113),
            .I(N__9099));
    InMux I__2029 (
            .O(N__9112),
            .I(N__9096));
    LocalMux I__2028 (
            .O(N__9109),
            .I(N__9085));
    LocalMux I__2027 (
            .O(N__9104),
            .I(N__9085));
    Span4Mux_v I__2026 (
            .O(N__9099),
            .I(N__9085));
    LocalMux I__2025 (
            .O(N__9096),
            .I(N__9085));
    InMux I__2024 (
            .O(N__9095),
            .I(N__9082));
    InMux I__2023 (
            .O(N__9094),
            .I(N__9079));
    Span4Mux_h I__2022 (
            .O(N__9085),
            .I(N__9076));
    LocalMux I__2021 (
            .O(N__9082),
            .I(\U712_CHIP_RAM.N_379 ));
    LocalMux I__2020 (
            .O(N__9079),
            .I(\U712_CHIP_RAM.N_379 ));
    Odrv4 I__2019 (
            .O(N__9076),
            .I(\U712_CHIP_RAM.N_379 ));
    InMux I__2018 (
            .O(N__9069),
            .I(N__9066));
    LocalMux I__2017 (
            .O(N__9066),
            .I(N__9063));
    Odrv4 I__2016 (
            .O(N__9063),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__2015 (
            .O(N__9060),
            .I(N__9057));
    LocalMux I__2014 (
            .O(N__9057),
            .I(N__9054));
    Span4Mux_s3_h I__2013 (
            .O(N__9054),
            .I(N__9051));
    Sp12to4 I__2012 (
            .O(N__9051),
            .I(N__9048));
    Span12Mux_s11_v I__2011 (
            .O(N__9048),
            .I(N__9045));
    Odrv12 I__2010 (
            .O(N__9045),
            .I(CMA_c_6));
    InMux I__2009 (
            .O(N__9042),
            .I(N__9039));
    LocalMux I__2008 (
            .O(N__9039),
            .I(N__9006));
    ClkMux I__2007 (
            .O(N__9038),
            .I(N__8916));
    ClkMux I__2006 (
            .O(N__9037),
            .I(N__8916));
    ClkMux I__2005 (
            .O(N__9036),
            .I(N__8916));
    ClkMux I__2004 (
            .O(N__9035),
            .I(N__8916));
    ClkMux I__2003 (
            .O(N__9034),
            .I(N__8916));
    ClkMux I__2002 (
            .O(N__9033),
            .I(N__8916));
    ClkMux I__2001 (
            .O(N__9032),
            .I(N__8916));
    ClkMux I__2000 (
            .O(N__9031),
            .I(N__8916));
    ClkMux I__1999 (
            .O(N__9030),
            .I(N__8916));
    ClkMux I__1998 (
            .O(N__9029),
            .I(N__8916));
    ClkMux I__1997 (
            .O(N__9028),
            .I(N__8916));
    ClkMux I__1996 (
            .O(N__9027),
            .I(N__8916));
    ClkMux I__1995 (
            .O(N__9026),
            .I(N__8916));
    ClkMux I__1994 (
            .O(N__9025),
            .I(N__8916));
    ClkMux I__1993 (
            .O(N__9024),
            .I(N__8916));
    ClkMux I__1992 (
            .O(N__9023),
            .I(N__8916));
    ClkMux I__1991 (
            .O(N__9022),
            .I(N__8916));
    ClkMux I__1990 (
            .O(N__9021),
            .I(N__8916));
    ClkMux I__1989 (
            .O(N__9020),
            .I(N__8916));
    ClkMux I__1988 (
            .O(N__9019),
            .I(N__8916));
    ClkMux I__1987 (
            .O(N__9018),
            .I(N__8916));
    ClkMux I__1986 (
            .O(N__9017),
            .I(N__8916));
    ClkMux I__1985 (
            .O(N__9016),
            .I(N__8916));
    ClkMux I__1984 (
            .O(N__9015),
            .I(N__8916));
    ClkMux I__1983 (
            .O(N__9014),
            .I(N__8916));
    ClkMux I__1982 (
            .O(N__9013),
            .I(N__8916));
    ClkMux I__1981 (
            .O(N__9012),
            .I(N__8916));
    ClkMux I__1980 (
            .O(N__9011),
            .I(N__8916));
    ClkMux I__1979 (
            .O(N__9010),
            .I(N__8916));
    ClkMux I__1978 (
            .O(N__9009),
            .I(N__8916));
    Glb2LocalMux I__1977 (
            .O(N__9006),
            .I(N__8916));
    ClkMux I__1976 (
            .O(N__9005),
            .I(N__8916));
    ClkMux I__1975 (
            .O(N__9004),
            .I(N__8916));
    ClkMux I__1974 (
            .O(N__9003),
            .I(N__8916));
    ClkMux I__1973 (
            .O(N__9002),
            .I(N__8916));
    ClkMux I__1972 (
            .O(N__9001),
            .I(N__8916));
    ClkMux I__1971 (
            .O(N__9000),
            .I(N__8916));
    ClkMux I__1970 (
            .O(N__8999),
            .I(N__8916));
    ClkMux I__1969 (
            .O(N__8998),
            .I(N__8916));
    ClkMux I__1968 (
            .O(N__8997),
            .I(N__8916));
    GlobalMux I__1967 (
            .O(N__8916),
            .I(CLK80_PLL));
    CEMux I__1966 (
            .O(N__8913),
            .I(N__8909));
    CEMux I__1965 (
            .O(N__8912),
            .I(N__8904));
    LocalMux I__1964 (
            .O(N__8909),
            .I(N__8901));
    CEMux I__1963 (
            .O(N__8908),
            .I(N__8898));
    CEMux I__1962 (
            .O(N__8907),
            .I(N__8895));
    LocalMux I__1961 (
            .O(N__8904),
            .I(N__8892));
    Span4Mux_v I__1960 (
            .O(N__8901),
            .I(N__8888));
    LocalMux I__1959 (
            .O(N__8898),
            .I(N__8885));
    LocalMux I__1958 (
            .O(N__8895),
            .I(N__8880));
    Span4Mux_v I__1957 (
            .O(N__8892),
            .I(N__8880));
    CEMux I__1956 (
            .O(N__8891),
            .I(N__8877));
    Span4Mux_h I__1955 (
            .O(N__8888),
            .I(N__8872));
    Span4Mux_v I__1954 (
            .O(N__8885),
            .I(N__8872));
    Span4Mux_h I__1953 (
            .O(N__8880),
            .I(N__8869));
    LocalMux I__1952 (
            .O(N__8877),
            .I(N__8866));
    Odrv4 I__1951 (
            .O(N__8872),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__1950 (
            .O(N__8869),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv12 I__1949 (
            .O(N__8866),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    InMux I__1948 (
            .O(N__8859),
            .I(N__8853));
    InMux I__1947 (
            .O(N__8858),
            .I(N__8853));
    LocalMux I__1946 (
            .O(N__8853),
            .I(N__8850));
    Odrv12 I__1945 (
            .O(N__8850),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1944 (
            .O(N__8847),
            .I(N__8844));
    LocalMux I__1943 (
            .O(N__8844),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__1942 (
            .O(N__8841),
            .I(N__8838));
    LocalMux I__1941 (
            .O(N__8838),
            .I(N__8835));
    Span4Mux_s3_v I__1940 (
            .O(N__8835),
            .I(N__8832));
    Span4Mux_v I__1939 (
            .O(N__8832),
            .I(N__8829));
    Span4Mux_v I__1938 (
            .O(N__8829),
            .I(N__8826));
    Span4Mux_h I__1937 (
            .O(N__8826),
            .I(N__8823));
    Odrv4 I__1936 (
            .O(N__8823),
            .I(CMA_c_0));
    InMux I__1935 (
            .O(N__8820),
            .I(N__8817));
    LocalMux I__1934 (
            .O(N__8817),
            .I(N__8813));
    InMux I__1933 (
            .O(N__8816),
            .I(N__8810));
    Span4Mux_v I__1932 (
            .O(N__8813),
            .I(N__8804));
    LocalMux I__1931 (
            .O(N__8810),
            .I(N__8804));
    InMux I__1930 (
            .O(N__8809),
            .I(N__8801));
    Span4Mux_h I__1929 (
            .O(N__8804),
            .I(N__8796));
    LocalMux I__1928 (
            .O(N__8801),
            .I(N__8796));
    Span4Mux_v I__1927 (
            .O(N__8796),
            .I(N__8792));
    InMux I__1926 (
            .O(N__8795),
            .I(N__8789));
    Span4Mux_v I__1925 (
            .O(N__8792),
            .I(N__8786));
    LocalMux I__1924 (
            .O(N__8789),
            .I(N__8783));
    Sp12to4 I__1923 (
            .O(N__8786),
            .I(N__8778));
    Span12Mux_v I__1922 (
            .O(N__8783),
            .I(N__8778));
    Span12Mux_h I__1921 (
            .O(N__8778),
            .I(N__8775));
    Odrv12 I__1920 (
            .O(N__8775),
            .I(DRA_c_2));
    InMux I__1919 (
            .O(N__8772),
            .I(N__8769));
    LocalMux I__1918 (
            .O(N__8769),
            .I(N__8766));
    Span4Mux_v I__1917 (
            .O(N__8766),
            .I(N__8763));
    Odrv4 I__1916 (
            .O(N__8763),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    IoInMux I__1915 (
            .O(N__8760),
            .I(N__8757));
    LocalMux I__1914 (
            .O(N__8757),
            .I(N__8754));
    Span4Mux_s2_h I__1913 (
            .O(N__8754),
            .I(N__8751));
    Sp12to4 I__1912 (
            .O(N__8751),
            .I(N__8748));
    Span12Mux_v I__1911 (
            .O(N__8748),
            .I(N__8745));
    Span12Mux_h I__1910 (
            .O(N__8745),
            .I(N__8742));
    Odrv12 I__1909 (
            .O(N__8742),
            .I(N_295_i));
    IoInMux I__1908 (
            .O(N__8739),
            .I(N__8736));
    LocalMux I__1907 (
            .O(N__8736),
            .I(N__8733));
    Span4Mux_s2_h I__1906 (
            .O(N__8733),
            .I(N__8730));
    Sp12to4 I__1905 (
            .O(N__8730),
            .I(N__8727));
    Span12Mux_s11_v I__1904 (
            .O(N__8727),
            .I(N__8724));
    Span12Mux_h I__1903 (
            .O(N__8724),
            .I(N__8721));
    Odrv12 I__1902 (
            .O(N__8721),
            .I(N_299_i));
    IoInMux I__1901 (
            .O(N__8718),
            .I(N__8715));
    LocalMux I__1900 (
            .O(N__8715),
            .I(N__8712));
    IoSpan4Mux I__1899 (
            .O(N__8712),
            .I(N__8709));
    Span4Mux_s3_v I__1898 (
            .O(N__8709),
            .I(N__8703));
    InMux I__1897 (
            .O(N__8708),
            .I(N__8696));
    InMux I__1896 (
            .O(N__8707),
            .I(N__8696));
    InMux I__1895 (
            .O(N__8706),
            .I(N__8696));
    Span4Mux_v I__1894 (
            .O(N__8703),
            .I(N__8693));
    LocalMux I__1893 (
            .O(N__8696),
            .I(N__8690));
    Sp12to4 I__1892 (
            .O(N__8693),
            .I(N__8686));
    Span4Mux_v I__1891 (
            .O(N__8690),
            .I(N__8683));
    InMux I__1890 (
            .O(N__8689),
            .I(N__8680));
    Span12Mux_v I__1889 (
            .O(N__8686),
            .I(N__8672));
    Sp12to4 I__1888 (
            .O(N__8683),
            .I(N__8672));
    LocalMux I__1887 (
            .O(N__8680),
            .I(N__8672));
    InMux I__1886 (
            .O(N__8679),
            .I(N__8669));
    Odrv12 I__1885 (
            .O(N__8672),
            .I(DBENn_c));
    LocalMux I__1884 (
            .O(N__8669),
            .I(DBENn_c));
    CascadeMux I__1883 (
            .O(N__8664),
            .I(N__8659));
    CascadeMux I__1882 (
            .O(N__8663),
            .I(N__8656));
    CascadeMux I__1881 (
            .O(N__8662),
            .I(N__8652));
    InMux I__1880 (
            .O(N__8659),
            .I(N__8649));
    InMux I__1879 (
            .O(N__8656),
            .I(N__8644));
    InMux I__1878 (
            .O(N__8655),
            .I(N__8644));
    InMux I__1877 (
            .O(N__8652),
            .I(N__8641));
    LocalMux I__1876 (
            .O(N__8649),
            .I(N__8635));
    LocalMux I__1875 (
            .O(N__8644),
            .I(N__8635));
    LocalMux I__1874 (
            .O(N__8641),
            .I(N__8632));
    InMux I__1873 (
            .O(N__8640),
            .I(N__8629));
    Span4Mux_h I__1872 (
            .O(N__8635),
            .I(N__8621));
    Span4Mux_v I__1871 (
            .O(N__8632),
            .I(N__8621));
    LocalMux I__1870 (
            .O(N__8629),
            .I(N__8621));
    InMux I__1869 (
            .O(N__8628),
            .I(N__8615));
    Span4Mux_h I__1868 (
            .O(N__8621),
            .I(N__8612));
    InMux I__1867 (
            .O(N__8620),
            .I(N__8609));
    InMux I__1866 (
            .O(N__8619),
            .I(N__8604));
    InMux I__1865 (
            .O(N__8618),
            .I(N__8604));
    LocalMux I__1864 (
            .O(N__8615),
            .I(N__8601));
    Odrv4 I__1863 (
            .O(N__8612),
            .I(DMA_CYCLEm));
    LocalMux I__1862 (
            .O(N__8609),
            .I(DMA_CYCLEm));
    LocalMux I__1861 (
            .O(N__8604),
            .I(DMA_CYCLEm));
    Odrv4 I__1860 (
            .O(N__8601),
            .I(DMA_CYCLEm));
    IoInMux I__1859 (
            .O(N__8592),
            .I(N__8589));
    LocalMux I__1858 (
            .O(N__8589),
            .I(N__8586));
    Span12Mux_s2_h I__1857 (
            .O(N__8586),
            .I(N__8583));
    Span12Mux_h I__1856 (
            .O(N__8583),
            .I(N__8580));
    Span12Mux_v I__1855 (
            .O(N__8580),
            .I(N__8577));
    Odrv12 I__1854 (
            .O(N__8577),
            .I(N_297_i));
    InMux I__1853 (
            .O(N__8574),
            .I(N__8571));
    LocalMux I__1852 (
            .O(N__8571),
            .I(\U712_BYTE_ENABLE.N_528 ));
    CascadeMux I__1851 (
            .O(N__8568),
            .I(\U712_BYTE_ENABLE.N_377_cascade_ ));
    InMux I__1850 (
            .O(N__8565),
            .I(N__8562));
    LocalMux I__1849 (
            .O(N__8562),
            .I(N__8559));
    Odrv4 I__1848 (
            .O(N__8559),
            .I(\U712_BYTE_ENABLE.N_508 ));
    InMux I__1847 (
            .O(N__8556),
            .I(N__8553));
    LocalMux I__1846 (
            .O(N__8553),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1845 (
            .O(N__8550),
            .I(N__8547));
    LocalMux I__1844 (
            .O(N__8547),
            .I(N__8544));
    Odrv4 I__1843 (
            .O(N__8544),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__1842 (
            .O(N__8541),
            .I(N__8538));
    LocalMux I__1841 (
            .O(N__8538),
            .I(N__8535));
    Odrv4 I__1840 (
            .O(N__8535),
            .I(\U712_CHIP_RAM.un3_DMA_CYCLE_START ));
    InMux I__1839 (
            .O(N__8532),
            .I(N__8526));
    InMux I__1838 (
            .O(N__8531),
            .I(N__8526));
    LocalMux I__1837 (
            .O(N__8526),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    CascadeMux I__1836 (
            .O(N__8523),
            .I(N__8512));
    InMux I__1835 (
            .O(N__8522),
            .I(N__8507));
    InMux I__1834 (
            .O(N__8521),
            .I(N__8507));
    InMux I__1833 (
            .O(N__8520),
            .I(N__8498));
    InMux I__1832 (
            .O(N__8519),
            .I(N__8498));
    InMux I__1831 (
            .O(N__8518),
            .I(N__8489));
    InMux I__1830 (
            .O(N__8517),
            .I(N__8486));
    InMux I__1829 (
            .O(N__8516),
            .I(N__8483));
    InMux I__1828 (
            .O(N__8515),
            .I(N__8476));
    InMux I__1827 (
            .O(N__8512),
            .I(N__8476));
    LocalMux I__1826 (
            .O(N__8507),
            .I(N__8473));
    InMux I__1825 (
            .O(N__8506),
            .I(N__8470));
    InMux I__1824 (
            .O(N__8505),
            .I(N__8467));
    InMux I__1823 (
            .O(N__8504),
            .I(N__8462));
    InMux I__1822 (
            .O(N__8503),
            .I(N__8462));
    LocalMux I__1821 (
            .O(N__8498),
            .I(N__8459));
    InMux I__1820 (
            .O(N__8497),
            .I(N__8456));
    InMux I__1819 (
            .O(N__8496),
            .I(N__8453));
    InMux I__1818 (
            .O(N__8495),
            .I(N__8448));
    InMux I__1817 (
            .O(N__8494),
            .I(N__8448));
    InMux I__1816 (
            .O(N__8493),
            .I(N__8443));
    InMux I__1815 (
            .O(N__8492),
            .I(N__8443));
    LocalMux I__1814 (
            .O(N__8489),
            .I(N__8436));
    LocalMux I__1813 (
            .O(N__8486),
            .I(N__8436));
    LocalMux I__1812 (
            .O(N__8483),
            .I(N__8436));
    InMux I__1811 (
            .O(N__8482),
            .I(N__8433));
    InMux I__1810 (
            .O(N__8481),
            .I(N__8422));
    LocalMux I__1809 (
            .O(N__8476),
            .I(N__8419));
    Span4Mux_h I__1808 (
            .O(N__8473),
            .I(N__8410));
    LocalMux I__1807 (
            .O(N__8470),
            .I(N__8410));
    LocalMux I__1806 (
            .O(N__8467),
            .I(N__8410));
    LocalMux I__1805 (
            .O(N__8462),
            .I(N__8410));
    Span4Mux_v I__1804 (
            .O(N__8459),
            .I(N__8407));
    LocalMux I__1803 (
            .O(N__8456),
            .I(N__8404));
    LocalMux I__1802 (
            .O(N__8453),
            .I(N__8397));
    LocalMux I__1801 (
            .O(N__8448),
            .I(N__8397));
    LocalMux I__1800 (
            .O(N__8443),
            .I(N__8397));
    Sp12to4 I__1799 (
            .O(N__8436),
            .I(N__8392));
    LocalMux I__1798 (
            .O(N__8433),
            .I(N__8392));
    InMux I__1797 (
            .O(N__8432),
            .I(N__8385));
    InMux I__1796 (
            .O(N__8431),
            .I(N__8385));
    InMux I__1795 (
            .O(N__8430),
            .I(N__8385));
    InMux I__1794 (
            .O(N__8429),
            .I(N__8378));
    InMux I__1793 (
            .O(N__8428),
            .I(N__8378));
    InMux I__1792 (
            .O(N__8427),
            .I(N__8378));
    InMux I__1791 (
            .O(N__8426),
            .I(N__8373));
    InMux I__1790 (
            .O(N__8425),
            .I(N__8373));
    LocalMux I__1789 (
            .O(N__8422),
            .I(N__8370));
    Span4Mux_v I__1788 (
            .O(N__8419),
            .I(N__8365));
    Span4Mux_v I__1787 (
            .O(N__8410),
            .I(N__8365));
    Span4Mux_h I__1786 (
            .O(N__8407),
            .I(N__8358));
    Span4Mux_v I__1785 (
            .O(N__8404),
            .I(N__8358));
    Span4Mux_v I__1784 (
            .O(N__8397),
            .I(N__8358));
    Span12Mux_v I__1783 (
            .O(N__8392),
            .I(N__8349));
    LocalMux I__1782 (
            .O(N__8385),
            .I(N__8349));
    LocalMux I__1781 (
            .O(N__8378),
            .I(N__8349));
    LocalMux I__1780 (
            .O(N__8373),
            .I(N__8349));
    Span12Mux_v I__1779 (
            .O(N__8370),
            .I(N__8342));
    Sp12to4 I__1778 (
            .O(N__8365),
            .I(N__8342));
    Sp12to4 I__1777 (
            .O(N__8358),
            .I(N__8342));
    Span12Mux_h I__1776 (
            .O(N__8349),
            .I(N__8339));
    Span12Mux_h I__1775 (
            .O(N__8342),
            .I(N__8336));
    Odrv12 I__1774 (
            .O(N__8339),
            .I(RESETn_c));
    Odrv12 I__1773 (
            .O(N__8336),
            .I(RESETn_c));
    InMux I__1772 (
            .O(N__8331),
            .I(N__8328));
    LocalMux I__1771 (
            .O(N__8328),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__1770 (
            .O(N__8325),
            .I(N__8322));
    LocalMux I__1769 (
            .O(N__8322),
            .I(N__8319));
    Span4Mux_v I__1768 (
            .O(N__8319),
            .I(N__8316));
    Odrv4 I__1767 (
            .O(N__8316),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    InMux I__1766 (
            .O(N__8313),
            .I(N__8310));
    LocalMux I__1765 (
            .O(N__8310),
            .I(N__8307));
    Span4Mux_h I__1764 (
            .O(N__8307),
            .I(N__8304));
    Odrv4 I__1763 (
            .O(N__8304),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__1762 (
            .O(N__8301),
            .I(N__8298));
    LocalMux I__1761 (
            .O(N__8298),
            .I(N__8295));
    IoSpan4Mux I__1760 (
            .O(N__8295),
            .I(N__8292));
    Span4Mux_s3_h I__1759 (
            .O(N__8292),
            .I(N__8289));
    Sp12to4 I__1758 (
            .O(N__8289),
            .I(N__8286));
    Span12Mux_h I__1757 (
            .O(N__8286),
            .I(N__8283));
    Odrv12 I__1756 (
            .O(N__8283),
            .I(CMA_c_3));
    InMux I__1755 (
            .O(N__8280),
            .I(N__8276));
    InMux I__1754 (
            .O(N__8279),
            .I(N__8273));
    LocalMux I__1753 (
            .O(N__8276),
            .I(N__8268));
    LocalMux I__1752 (
            .O(N__8273),
            .I(N__8265));
    InMux I__1751 (
            .O(N__8272),
            .I(N__8262));
    InMux I__1750 (
            .O(N__8271),
            .I(N__8259));
    Span4Mux_v I__1749 (
            .O(N__8268),
            .I(N__8252));
    Span4Mux_h I__1748 (
            .O(N__8265),
            .I(N__8252));
    LocalMux I__1747 (
            .O(N__8262),
            .I(N__8252));
    LocalMux I__1746 (
            .O(N__8259),
            .I(N__8247));
    Sp12to4 I__1745 (
            .O(N__8252),
            .I(N__8247));
    Span12Mux_v I__1744 (
            .O(N__8247),
            .I(N__8244));
    Span12Mux_h I__1743 (
            .O(N__8244),
            .I(N__8241));
    Odrv12 I__1742 (
            .O(N__8241),
            .I(DRA_c_3));
    InMux I__1741 (
            .O(N__8238),
            .I(N__8235));
    LocalMux I__1740 (
            .O(N__8235),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__1739 (
            .O(N__8232),
            .I(N__8228));
    InMux I__1738 (
            .O(N__8231),
            .I(N__8221));
    LocalMux I__1737 (
            .O(N__8228),
            .I(N__8218));
    InMux I__1736 (
            .O(N__8227),
            .I(N__8213));
    InMux I__1735 (
            .O(N__8226),
            .I(N__8213));
    InMux I__1734 (
            .O(N__8225),
            .I(N__8208));
    InMux I__1733 (
            .O(N__8224),
            .I(N__8208));
    LocalMux I__1732 (
            .O(N__8221),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    Odrv4 I__1731 (
            .O(N__8218),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1730 (
            .O(N__8213),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1729 (
            .O(N__8208),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    CascadeMux I__1728 (
            .O(N__8199),
            .I(N__8189));
    InMux I__1727 (
            .O(N__8198),
            .I(N__8180));
    InMux I__1726 (
            .O(N__8197),
            .I(N__8180));
    InMux I__1725 (
            .O(N__8196),
            .I(N__8180));
    InMux I__1724 (
            .O(N__8195),
            .I(N__8175));
    InMux I__1723 (
            .O(N__8194),
            .I(N__8172));
    InMux I__1722 (
            .O(N__8193),
            .I(N__8169));
    InMux I__1721 (
            .O(N__8192),
            .I(N__8164));
    InMux I__1720 (
            .O(N__8189),
            .I(N__8164));
    InMux I__1719 (
            .O(N__8188),
            .I(N__8159));
    InMux I__1718 (
            .O(N__8187),
            .I(N__8159));
    LocalMux I__1717 (
            .O(N__8180),
            .I(N__8156));
    InMux I__1716 (
            .O(N__8179),
            .I(N__8151));
    InMux I__1715 (
            .O(N__8178),
            .I(N__8151));
    LocalMux I__1714 (
            .O(N__8175),
            .I(N__8148));
    LocalMux I__1713 (
            .O(N__8172),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1712 (
            .O(N__8169),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1711 (
            .O(N__8164),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1710 (
            .O(N__8159),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1709 (
            .O(N__8156),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1708 (
            .O(N__8151),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1707 (
            .O(N__8148),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    CascadeMux I__1706 (
            .O(N__8133),
            .I(N__8129));
    InMux I__1705 (
            .O(N__8132),
            .I(N__8121));
    InMux I__1704 (
            .O(N__8129),
            .I(N__8118));
    InMux I__1703 (
            .O(N__8128),
            .I(N__8109));
    InMux I__1702 (
            .O(N__8127),
            .I(N__8109));
    InMux I__1701 (
            .O(N__8126),
            .I(N__8109));
    InMux I__1700 (
            .O(N__8125),
            .I(N__8109));
    InMux I__1699 (
            .O(N__8124),
            .I(N__8106));
    LocalMux I__1698 (
            .O(N__8121),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1697 (
            .O(N__8118),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1696 (
            .O(N__8109),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1695 (
            .O(N__8106),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    InMux I__1694 (
            .O(N__8097),
            .I(N__8090));
    InMux I__1693 (
            .O(N__8096),
            .I(N__8083));
    InMux I__1692 (
            .O(N__8095),
            .I(N__8083));
    InMux I__1691 (
            .O(N__8094),
            .I(N__8078));
    InMux I__1690 (
            .O(N__8093),
            .I(N__8078));
    LocalMux I__1689 (
            .O(N__8090),
            .I(N__8075));
    InMux I__1688 (
            .O(N__8089),
            .I(N__8070));
    InMux I__1687 (
            .O(N__8088),
            .I(N__8070));
    LocalMux I__1686 (
            .O(N__8083),
            .I(N__8067));
    LocalMux I__1685 (
            .O(N__8078),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    Odrv12 I__1684 (
            .O(N__8075),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    LocalMux I__1683 (
            .O(N__8070),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    Odrv4 I__1682 (
            .O(N__8067),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    CascadeMux I__1681 (
            .O(N__8058),
            .I(N__8055));
    InMux I__1680 (
            .O(N__8055),
            .I(N__8052));
    LocalMux I__1679 (
            .O(N__8052),
            .I(\U712_REG_SM.N_479 ));
    CascadeMux I__1678 (
            .O(N__8049),
            .I(N__8044));
    InMux I__1677 (
            .O(N__8048),
            .I(N__8038));
    InMux I__1676 (
            .O(N__8047),
            .I(N__8038));
    InMux I__1675 (
            .O(N__8044),
            .I(N__8035));
    InMux I__1674 (
            .O(N__8043),
            .I(N__8032));
    LocalMux I__1673 (
            .O(N__8038),
            .I(N__8027));
    LocalMux I__1672 (
            .O(N__8035),
            .I(N__8027));
    LocalMux I__1671 (
            .O(N__8032),
            .I(N__8024));
    Span4Mux_v I__1670 (
            .O(N__8027),
            .I(N__8021));
    Sp12to4 I__1669 (
            .O(N__8024),
            .I(N__8018));
    Sp12to4 I__1668 (
            .O(N__8021),
            .I(N__8015));
    Span12Mux_v I__1667 (
            .O(N__8018),
            .I(N__8010));
    Span12Mux_h I__1666 (
            .O(N__8015),
            .I(N__8010));
    Span12Mux_v I__1665 (
            .O(N__8010),
            .I(N__8007));
    Odrv12 I__1664 (
            .O(N__8007),
            .I(CLK40_PLL_i));
    IoInMux I__1663 (
            .O(N__8004),
            .I(N__7999));
    IoInMux I__1662 (
            .O(N__8003),
            .I(N__7996));
    IoInMux I__1661 (
            .O(N__8002),
            .I(N__7993));
    LocalMux I__1660 (
            .O(N__7999),
            .I(N__7988));
    LocalMux I__1659 (
            .O(N__7996),
            .I(N__7988));
    LocalMux I__1658 (
            .O(N__7993),
            .I(N__7985));
    IoSpan4Mux I__1657 (
            .O(N__7988),
            .I(N__7982));
    Span4Mux_s3_h I__1656 (
            .O(N__7985),
            .I(N__7979));
    Span4Mux_s1_v I__1655 (
            .O(N__7982),
            .I(N__7976));
    Sp12to4 I__1654 (
            .O(N__7979),
            .I(N__7973));
    Sp12to4 I__1653 (
            .O(N__7976),
            .I(N__7970));
    Span12Mux_v I__1652 (
            .O(N__7973),
            .I(N__7967));
    Span12Mux_h I__1651 (
            .O(N__7970),
            .I(N__7962));
    Span12Mux_h I__1650 (
            .O(N__7967),
            .I(N__7962));
    Odrv12 I__1649 (
            .O(N__7962),
            .I(CLK40_PLL_i_i));
    IoInMux I__1648 (
            .O(N__7959),
            .I(N__7956));
    LocalMux I__1647 (
            .O(N__7956),
            .I(N__7953));
    Span12Mux_s5_v I__1646 (
            .O(N__7953),
            .I(N__7950));
    Odrv12 I__1645 (
            .O(N__7950),
            .I(RESETn_c_i));
    InMux I__1644 (
            .O(N__7947),
            .I(N__7944));
    LocalMux I__1643 (
            .O(N__7944),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__1642 (
            .O(N__7941),
            .I(N__7938));
    LocalMux I__1641 (
            .O(N__7938),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__1640 (
            .O(N__7935),
            .I(N__7932));
    LocalMux I__1639 (
            .O(N__7932),
            .I(N__7929));
    Odrv4 I__1638 (
            .O(N__7929),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1637 (
            .O(N__7926),
            .I(N__7923));
    LocalMux I__1636 (
            .O(N__7923),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1635 (
            .O(N__7920),
            .I(N__7917));
    LocalMux I__1634 (
            .O(N__7917),
            .I(N__7914));
    Span4Mux_h I__1633 (
            .O(N__7914),
            .I(N__7911));
    Odrv4 I__1632 (
            .O(N__7911),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__1631 (
            .O(N__7908),
            .I(N__7905));
    LocalMux I__1630 (
            .O(N__7905),
            .I(N__7902));
    Odrv4 I__1629 (
            .O(N__7902),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    InMux I__1628 (
            .O(N__7899),
            .I(N__7895));
    InMux I__1627 (
            .O(N__7898),
            .I(N__7892));
    LocalMux I__1626 (
            .O(N__7895),
            .I(N__7889));
    LocalMux I__1625 (
            .O(N__7892),
            .I(N__7886));
    Odrv4 I__1624 (
            .O(N__7889),
            .I(\U712_REG_SM.N_661 ));
    Odrv12 I__1623 (
            .O(N__7886),
            .I(\U712_REG_SM.N_661 ));
    InMux I__1622 (
            .O(N__7881),
            .I(N__7876));
    InMux I__1621 (
            .O(N__7880),
            .I(N__7873));
    InMux I__1620 (
            .O(N__7879),
            .I(N__7870));
    LocalMux I__1619 (
            .O(N__7876),
            .I(\U712_REG_SM.N_389 ));
    LocalMux I__1618 (
            .O(N__7873),
            .I(\U712_REG_SM.N_389 ));
    LocalMux I__1617 (
            .O(N__7870),
            .I(\U712_REG_SM.N_389 ));
    CascadeMux I__1616 (
            .O(N__7863),
            .I(\U712_REG_SM.N_475_cascade_ ));
    IoInMux I__1615 (
            .O(N__7860),
            .I(N__7857));
    LocalMux I__1614 (
            .O(N__7857),
            .I(N__7854));
    Span4Mux_s2_v I__1613 (
            .O(N__7854),
            .I(N__7851));
    Span4Mux_h I__1612 (
            .O(N__7851),
            .I(N__7848));
    Sp12to4 I__1611 (
            .O(N__7848),
            .I(N__7845));
    Span12Mux_s9_v I__1610 (
            .O(N__7845),
            .I(N__7842));
    Odrv12 I__1609 (
            .O(N__7842),
            .I(N_57_i));
    InMux I__1608 (
            .O(N__7839),
            .I(N__7835));
    InMux I__1607 (
            .O(N__7838),
            .I(N__7832));
    LocalMux I__1606 (
            .O(N__7835),
            .I(N__7826));
    LocalMux I__1605 (
            .O(N__7832),
            .I(N__7826));
    InMux I__1604 (
            .O(N__7831),
            .I(N__7823));
    Odrv4 I__1603 (
            .O(N__7826),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1602 (
            .O(N__7823),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__1601 (
            .O(N__7818),
            .I(N__7815));
    LocalMux I__1600 (
            .O(N__7815),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    CascadeMux I__1599 (
            .O(N__7812),
            .I(N__7809));
    InMux I__1598 (
            .O(N__7809),
            .I(N__7804));
    InMux I__1597 (
            .O(N__7808),
            .I(N__7801));
    InMux I__1596 (
            .O(N__7807),
            .I(N__7798));
    LocalMux I__1595 (
            .O(N__7804),
            .I(N__7790));
    LocalMux I__1594 (
            .O(N__7801),
            .I(N__7790));
    LocalMux I__1593 (
            .O(N__7798),
            .I(N__7790));
    InMux I__1592 (
            .O(N__7797),
            .I(N__7787));
    Odrv4 I__1591 (
            .O(N__7790),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1590 (
            .O(N__7787),
            .I(DBR_SYNCZ0Z_1));
    CascadeMux I__1589 (
            .O(N__7782),
            .I(\U712_REG_SM.N_449_cascade_ ));
    InMux I__1588 (
            .O(N__7779),
            .I(N__7773));
    InMux I__1587 (
            .O(N__7778),
            .I(N__7773));
    LocalMux I__1586 (
            .O(N__7773),
            .I(N__7766));
    InMux I__1585 (
            .O(N__7772),
            .I(N__7763));
    InMux I__1584 (
            .O(N__7771),
            .I(N__7758));
    InMux I__1583 (
            .O(N__7770),
            .I(N__7758));
    InMux I__1582 (
            .O(N__7769),
            .I(N__7755));
    Span4Mux_h I__1581 (
            .O(N__7766),
            .I(N__7752));
    LocalMux I__1580 (
            .O(N__7763),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1579 (
            .O(N__7758),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1578 (
            .O(N__7755),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv4 I__1577 (
            .O(N__7752),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    InMux I__1576 (
            .O(N__7743),
            .I(N__7739));
    InMux I__1575 (
            .O(N__7742),
            .I(N__7736));
    LocalMux I__1574 (
            .O(N__7739),
            .I(\U712_REG_SM.START_RST_0_sqmuxa ));
    LocalMux I__1573 (
            .O(N__7736),
            .I(\U712_REG_SM.START_RST_0_sqmuxa ));
    CascadeMux I__1572 (
            .O(N__7731),
            .I(\U712_REG_SM.N_396_cascade_ ));
    CascadeMux I__1571 (
            .O(N__7728),
            .I(N__7725));
    InMux I__1570 (
            .O(N__7725),
            .I(N__7720));
    CascadeMux I__1569 (
            .O(N__7724),
            .I(N__7717));
    CascadeMux I__1568 (
            .O(N__7723),
            .I(N__7713));
    LocalMux I__1567 (
            .O(N__7720),
            .I(N__7709));
    InMux I__1566 (
            .O(N__7717),
            .I(N__7702));
    InMux I__1565 (
            .O(N__7716),
            .I(N__7702));
    InMux I__1564 (
            .O(N__7713),
            .I(N__7702));
    InMux I__1563 (
            .O(N__7712),
            .I(N__7697));
    Span4Mux_v I__1562 (
            .O(N__7709),
            .I(N__7690));
    LocalMux I__1561 (
            .O(N__7702),
            .I(N__7690));
    InMux I__1560 (
            .O(N__7701),
            .I(N__7685));
    InMux I__1559 (
            .O(N__7700),
            .I(N__7682));
    LocalMux I__1558 (
            .O(N__7697),
            .I(N__7679));
    InMux I__1557 (
            .O(N__7696),
            .I(N__7676));
    InMux I__1556 (
            .O(N__7695),
            .I(N__7673));
    Span4Mux_h I__1555 (
            .O(N__7690),
            .I(N__7670));
    InMux I__1554 (
            .O(N__7689),
            .I(N__7665));
    InMux I__1553 (
            .O(N__7688),
            .I(N__7665));
    LocalMux I__1552 (
            .O(N__7685),
            .I(N__7662));
    LocalMux I__1551 (
            .O(N__7682),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1550 (
            .O(N__7679),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1549 (
            .O(N__7676),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1548 (
            .O(N__7673),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1547 (
            .O(N__7670),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1546 (
            .O(N__7665),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1545 (
            .O(N__7662),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__1544 (
            .O(N__7647),
            .I(N__7644));
    LocalMux I__1543 (
            .O(N__7644),
            .I(\U712_REG_SM.un1_STATE_COUNT_4_i_i_0_0 ));
    InMux I__1542 (
            .O(N__7641),
            .I(N__7637));
    InMux I__1541 (
            .O(N__7640),
            .I(N__7634));
    LocalMux I__1540 (
            .O(N__7637),
            .I(N__7631));
    LocalMux I__1539 (
            .O(N__7634),
            .I(N__7628));
    Span4Mux_v I__1538 (
            .O(N__7631),
            .I(N__7623));
    Span4Mux_v I__1537 (
            .O(N__7628),
            .I(N__7623));
    Span4Mux_v I__1536 (
            .O(N__7623),
            .I(N__7620));
    Sp12to4 I__1535 (
            .O(N__7620),
            .I(N__7617));
    Span12Mux_h I__1534 (
            .O(N__7617),
            .I(N__7614));
    Odrv12 I__1533 (
            .O(N__7614),
            .I(TSn_c));
    CascadeMux I__1532 (
            .O(N__7611),
            .I(\U712_REG_SM.N_477_cascade_ ));
    InMux I__1531 (
            .O(N__7608),
            .I(N__7605));
    LocalMux I__1530 (
            .O(N__7605),
            .I(N__7602));
    Span4Mux_v I__1529 (
            .O(N__7602),
            .I(N__7599));
    Sp12to4 I__1528 (
            .O(N__7599),
            .I(N__7596));
    Span12Mux_h I__1527 (
            .O(N__7596),
            .I(N__7593));
    Span12Mux_v I__1526 (
            .O(N__7593),
            .I(N__7590));
    Odrv12 I__1525 (
            .O(N__7590),
            .I(REGSPACEn_c));
    IoInMux I__1524 (
            .O(N__7587),
            .I(N__7584));
    LocalMux I__1523 (
            .O(N__7584),
            .I(N__7581));
    Span4Mux_s0_v I__1522 (
            .O(N__7581),
            .I(N__7578));
    Span4Mux_v I__1521 (
            .O(N__7578),
            .I(N__7574));
    InMux I__1520 (
            .O(N__7577),
            .I(N__7571));
    Span4Mux_v I__1519 (
            .O(N__7574),
            .I(N__7568));
    LocalMux I__1518 (
            .O(N__7571),
            .I(N__7565));
    Sp12to4 I__1517 (
            .O(N__7568),
            .I(N__7562));
    Span4Mux_v I__1516 (
            .O(N__7565),
            .I(N__7559));
    Span12Mux_h I__1515 (
            .O(N__7562),
            .I(N__7556));
    Sp12to4 I__1514 (
            .O(N__7559),
            .I(N__7553));
    Span12Mux_v I__1513 (
            .O(N__7556),
            .I(N__7548));
    Span12Mux_h I__1512 (
            .O(N__7553),
            .I(N__7548));
    Odrv12 I__1511 (
            .O(N__7548),
            .I(A_c_10));
    InMux I__1510 (
            .O(N__7545),
            .I(N__7542));
    LocalMux I__1509 (
            .O(N__7542),
            .I(N__7539));
    Odrv4 I__1508 (
            .O(N__7539),
            .I(\U712_CHIP_RAM.N_422 ));
    InMux I__1507 (
            .O(N__7536),
            .I(N__7533));
    LocalMux I__1506 (
            .O(N__7533),
            .I(N__7530));
    Span4Mux_v I__1505 (
            .O(N__7530),
            .I(N__7527));
    Sp12to4 I__1504 (
            .O(N__7527),
            .I(N__7524));
    Span12Mux_h I__1503 (
            .O(N__7524),
            .I(N__7521));
    Span12Mux_v I__1502 (
            .O(N__7521),
            .I(N__7518));
    Odrv12 I__1501 (
            .O(N__7518),
            .I(A_c_3));
    InMux I__1500 (
            .O(N__7515),
            .I(N__7512));
    LocalMux I__1499 (
            .O(N__7512),
            .I(N__7509));
    Odrv4 I__1498 (
            .O(N__7509),
            .I(\U712_CHIP_RAM.N_445 ));
    InMux I__1497 (
            .O(N__7506),
            .I(N__7503));
    LocalMux I__1496 (
            .O(N__7503),
            .I(N__7500));
    Span4Mux_h I__1495 (
            .O(N__7500),
            .I(N__7496));
    InMux I__1494 (
            .O(N__7499),
            .I(N__7493));
    Span4Mux_h I__1493 (
            .O(N__7496),
            .I(N__7488));
    LocalMux I__1492 (
            .O(N__7493),
            .I(N__7488));
    Span4Mux_v I__1491 (
            .O(N__7488),
            .I(N__7485));
    Span4Mux_h I__1490 (
            .O(N__7485),
            .I(N__7482));
    Sp12to4 I__1489 (
            .O(N__7482),
            .I(N__7479));
    Odrv12 I__1488 (
            .O(N__7479),
            .I(DBRn_c));
    InMux I__1487 (
            .O(N__7476),
            .I(N__7473));
    LocalMux I__1486 (
            .O(N__7473),
            .I(DBR_SYNCZ0Z_0));
    InMux I__1485 (
            .O(N__7470),
            .I(N__7466));
    InMux I__1484 (
            .O(N__7469),
            .I(N__7463));
    LocalMux I__1483 (
            .O(N__7466),
            .I(N__7460));
    LocalMux I__1482 (
            .O(N__7463),
            .I(\U712_REG_SM.START_RSTZ0 ));
    Odrv4 I__1481 (
            .O(N__7460),
            .I(\U712_REG_SM.START_RSTZ0 ));
    InMux I__1480 (
            .O(N__7455),
            .I(N__7452));
    LocalMux I__1479 (
            .O(N__7452),
            .I(N__7449));
    Span4Mux_h I__1478 (
            .O(N__7449),
            .I(N__7446));
    Odrv4 I__1477 (
            .O(N__7446),
            .I(\U712_CYCLE_TERM.TACK_EN_RNOZ0Z_0 ));
    InMux I__1476 (
            .O(N__7443),
            .I(N__7439));
    InMux I__1475 (
            .O(N__7442),
            .I(N__7436));
    LocalMux I__1474 (
            .O(N__7439),
            .I(N__7433));
    LocalMux I__1473 (
            .O(N__7436),
            .I(N__7428));
    Span4Mux_h I__1472 (
            .O(N__7433),
            .I(N__7428));
    Odrv4 I__1471 (
            .O(N__7428),
            .I(\U712_CYCLE_TERM.un13_0 ));
    IoInMux I__1470 (
            .O(N__7425),
            .I(N__7422));
    LocalMux I__1469 (
            .O(N__7422),
            .I(N__7419));
    IoSpan4Mux I__1468 (
            .O(N__7419),
            .I(N__7415));
    IoInMux I__1467 (
            .O(N__7418),
            .I(N__7412));
    Span4Mux_s1_v I__1466 (
            .O(N__7415),
            .I(N__7409));
    LocalMux I__1465 (
            .O(N__7412),
            .I(N__7406));
    Span4Mux_v I__1464 (
            .O(N__7409),
            .I(N__7403));
    IoSpan4Mux I__1463 (
            .O(N__7406),
            .I(N__7400));
    Span4Mux_v I__1462 (
            .O(N__7403),
            .I(N__7397));
    Span4Mux_s2_h I__1461 (
            .O(N__7400),
            .I(N__7393));
    Span4Mux_v I__1460 (
            .O(N__7397),
            .I(N__7390));
    InMux I__1459 (
            .O(N__7396),
            .I(N__7387));
    Sp12to4 I__1458 (
            .O(N__7393),
            .I(N__7384));
    Span4Mux_h I__1457 (
            .O(N__7390),
            .I(N__7379));
    LocalMux I__1456 (
            .O(N__7387),
            .I(N__7379));
    Span12Mux_h I__1455 (
            .O(N__7384),
            .I(N__7376));
    Span4Mux_v I__1454 (
            .O(N__7379),
            .I(N__7373));
    Span12Mux_v I__1453 (
            .O(N__7376),
            .I(N__7369));
    Span4Mux_h I__1452 (
            .O(N__7373),
            .I(N__7366));
    InMux I__1451 (
            .O(N__7372),
            .I(N__7363));
    Odrv12 I__1450 (
            .O(N__7369),
            .I(TACK_EN));
    Odrv4 I__1449 (
            .O(N__7366),
            .I(TACK_EN));
    LocalMux I__1448 (
            .O(N__7363),
            .I(TACK_EN));
    IoInMux I__1447 (
            .O(N__7356),
            .I(N__7353));
    LocalMux I__1446 (
            .O(N__7353),
            .I(N__7350));
    IoSpan4Mux I__1445 (
            .O(N__7350),
            .I(N__7347));
    IoSpan4Mux I__1444 (
            .O(N__7347),
            .I(N__7344));
    Sp12to4 I__1443 (
            .O(N__7344),
            .I(N__7341));
    Span12Mux_s7_v I__1442 (
            .O(N__7341),
            .I(N__7338));
    Span12Mux_h I__1441 (
            .O(N__7338),
            .I(N__7335));
    Odrv12 I__1440 (
            .O(N__7335),
            .I(WEn_c));
    IoInMux I__1439 (
            .O(N__7332),
            .I(N__7329));
    LocalMux I__1438 (
            .O(N__7329),
            .I(N__7326));
    Span4Mux_s0_v I__1437 (
            .O(N__7326),
            .I(N__7323));
    Sp12to4 I__1436 (
            .O(N__7323),
            .I(N__7320));
    Span12Mux_h I__1435 (
            .O(N__7320),
            .I(N__7317));
    Odrv12 I__1434 (
            .O(N__7317),
            .I(CRCSn_c));
    InMux I__1433 (
            .O(N__7314),
            .I(N__7311));
    LocalMux I__1432 (
            .O(N__7311),
            .I(N__7308));
    Sp12to4 I__1431 (
            .O(N__7308),
            .I(N__7305));
    Span12Mux_v I__1430 (
            .O(N__7305),
            .I(N__7302));
    Span12Mux_h I__1429 (
            .O(N__7302),
            .I(N__7299));
    Odrv12 I__1428 (
            .O(N__7299),
            .I(A_c_19));
    IoInMux I__1427 (
            .O(N__7296),
            .I(N__7293));
    LocalMux I__1426 (
            .O(N__7293),
            .I(N__7290));
    IoSpan4Mux I__1425 (
            .O(N__7290),
            .I(N__7287));
    Span4Mux_s3_h I__1424 (
            .O(N__7287),
            .I(N__7284));
    Span4Mux_v I__1423 (
            .O(N__7284),
            .I(N__7281));
    Span4Mux_h I__1422 (
            .O(N__7281),
            .I(N__7278));
    Sp12to4 I__1421 (
            .O(N__7278),
            .I(N__7275));
    Odrv12 I__1420 (
            .O(N__7275),
            .I(CMA_c_9));
    InMux I__1419 (
            .O(N__7272),
            .I(N__7269));
    LocalMux I__1418 (
            .O(N__7269),
            .I(N__7266));
    Span12Mux_v I__1417 (
            .O(N__7266),
            .I(N__7263));
    Span12Mux_h I__1416 (
            .O(N__7263),
            .I(N__7260));
    Odrv12 I__1415 (
            .O(N__7260),
            .I(A_c_17));
    IoInMux I__1414 (
            .O(N__7257),
            .I(N__7254));
    LocalMux I__1413 (
            .O(N__7254),
            .I(N__7251));
    Span4Mux_s0_h I__1412 (
            .O(N__7251),
            .I(N__7248));
    Span4Mux_h I__1411 (
            .O(N__7248),
            .I(N__7245));
    Sp12to4 I__1410 (
            .O(N__7245),
            .I(N__7242));
    Span12Mux_s10_v I__1409 (
            .O(N__7242),
            .I(N__7239));
    Span12Mux_h I__1408 (
            .O(N__7239),
            .I(N__7236));
    Odrv12 I__1407 (
            .O(N__7236),
            .I(CMA_c_8));
    IoInMux I__1406 (
            .O(N__7233),
            .I(N__7230));
    LocalMux I__1405 (
            .O(N__7230),
            .I(N__7227));
    Span12Mux_s11_v I__1404 (
            .O(N__7227),
            .I(N__7224));
    Odrv12 I__1403 (
            .O(N__7224),
            .I(CMA_c_1));
    InMux I__1402 (
            .O(N__7221),
            .I(N__7217));
    InMux I__1401 (
            .O(N__7220),
            .I(N__7213));
    LocalMux I__1400 (
            .O(N__7217),
            .I(N__7209));
    InMux I__1399 (
            .O(N__7216),
            .I(N__7206));
    LocalMux I__1398 (
            .O(N__7213),
            .I(N__7203));
    CascadeMux I__1397 (
            .O(N__7212),
            .I(N__7199));
    Span4Mux_h I__1396 (
            .O(N__7209),
            .I(N__7196));
    LocalMux I__1395 (
            .O(N__7206),
            .I(N__7191));
    Span4Mux_h I__1394 (
            .O(N__7203),
            .I(N__7191));
    InMux I__1393 (
            .O(N__7202),
            .I(N__7186));
    InMux I__1392 (
            .O(N__7199),
            .I(N__7186));
    Odrv4 I__1391 (
            .O(N__7196),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1390 (
            .O(N__7191),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1389 (
            .O(N__7186),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1388 (
            .O(N__7179),
            .I(N__7176));
    LocalMux I__1387 (
            .O(N__7176),
            .I(N__7173));
    Span4Mux_s1_v I__1386 (
            .O(N__7173),
            .I(N__7170));
    Span4Mux_v I__1385 (
            .O(N__7170),
            .I(N__7167));
    Sp12to4 I__1384 (
            .O(N__7167),
            .I(N__7164));
    Span12Mux_h I__1383 (
            .O(N__7164),
            .I(N__7161));
    Odrv12 I__1382 (
            .O(N__7161),
            .I(CMA_c_10));
    IoInMux I__1381 (
            .O(N__7158),
            .I(N__7155));
    LocalMux I__1380 (
            .O(N__7155),
            .I(N__7152));
    IoSpan4Mux I__1379 (
            .O(N__7152),
            .I(N__7149));
    Sp12to4 I__1378 (
            .O(N__7149),
            .I(N__7146));
    Span12Mux_s7_v I__1377 (
            .O(N__7146),
            .I(N__7143));
    Odrv12 I__1376 (
            .O(N__7143),
            .I(CMA_c_2));
    InMux I__1375 (
            .O(N__7140),
            .I(N__7137));
    LocalMux I__1374 (
            .O(N__7137),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    InMux I__1373 (
            .O(N__7134),
            .I(N__7131));
    LocalMux I__1372 (
            .O(N__7131),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    InMux I__1371 (
            .O(N__7128),
            .I(N__7125));
    LocalMux I__1370 (
            .O(N__7125),
            .I(N__7122));
    Span4Mux_h I__1369 (
            .O(N__7122),
            .I(N__7117));
    InMux I__1368 (
            .O(N__7121),
            .I(N__7114));
    InMux I__1367 (
            .O(N__7120),
            .I(N__7110));
    Span4Mux_v I__1366 (
            .O(N__7117),
            .I(N__7107));
    LocalMux I__1365 (
            .O(N__7114),
            .I(N__7104));
    InMux I__1364 (
            .O(N__7113),
            .I(N__7101));
    LocalMux I__1363 (
            .O(N__7110),
            .I(N__7094));
    Span4Mux_v I__1362 (
            .O(N__7107),
            .I(N__7094));
    Span4Mux_h I__1361 (
            .O(N__7104),
            .I(N__7091));
    LocalMux I__1360 (
            .O(N__7101),
            .I(N__7088));
    InMux I__1359 (
            .O(N__7100),
            .I(N__7085));
    InMux I__1358 (
            .O(N__7099),
            .I(N__7082));
    Odrv4 I__1357 (
            .O(N__7094),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1356 (
            .O(N__7091),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1355 (
            .O(N__7088),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1354 (
            .O(N__7085),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1353 (
            .O(N__7082),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    InMux I__1352 (
            .O(N__7071),
            .I(N__7067));
    CascadeMux I__1351 (
            .O(N__7070),
            .I(N__7062));
    LocalMux I__1350 (
            .O(N__7067),
            .I(N__7059));
    InMux I__1349 (
            .O(N__7066),
            .I(N__7056));
    InMux I__1348 (
            .O(N__7065),
            .I(N__7053));
    InMux I__1347 (
            .O(N__7062),
            .I(N__7049));
    Span4Mux_v I__1346 (
            .O(N__7059),
            .I(N__7044));
    LocalMux I__1345 (
            .O(N__7056),
            .I(N__7044));
    LocalMux I__1344 (
            .O(N__7053),
            .I(N__7041));
    InMux I__1343 (
            .O(N__7052),
            .I(N__7038));
    LocalMux I__1342 (
            .O(N__7049),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1341 (
            .O(N__7044),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1340 (
            .O(N__7041),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1339 (
            .O(N__7038),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    InMux I__1338 (
            .O(N__7029),
            .I(N__7023));
    InMux I__1337 (
            .O(N__7028),
            .I(N__7023));
    LocalMux I__1336 (
            .O(N__7023),
            .I(\U712_CHIP_RAM.CMA_5_i_0_8 ));
    CascadeMux I__1335 (
            .O(N__7020),
            .I(\U712_REG_SM.N_374_cascade_ ));
    InMux I__1334 (
            .O(N__7017),
            .I(N__7014));
    LocalMux I__1333 (
            .O(N__7014),
            .I(\U712_REG_SM.N_417 ));
    IoInMux I__1332 (
            .O(N__7011),
            .I(N__7008));
    LocalMux I__1331 (
            .O(N__7008),
            .I(N__7005));
    IoSpan4Mux I__1330 (
            .O(N__7005),
            .I(N__7002));
    Span4Mux_s3_h I__1329 (
            .O(N__7002),
            .I(N__6999));
    Span4Mux_v I__1328 (
            .O(N__6999),
            .I(N__6996));
    Span4Mux_h I__1327 (
            .O(N__6996),
            .I(N__6993));
    Sp12to4 I__1326 (
            .O(N__6993),
            .I(N__6989));
    InMux I__1325 (
            .O(N__6992),
            .I(N__6986));
    Span12Mux_h I__1324 (
            .O(N__6989),
            .I(N__6981));
    LocalMux I__1323 (
            .O(N__6986),
            .I(N__6981));
    Span12Mux_h I__1322 (
            .O(N__6981),
            .I(N__6978));
    Odrv12 I__1321 (
            .O(N__6978),
            .I(C3_c));
    InMux I__1320 (
            .O(N__6975),
            .I(N__6972));
    LocalMux I__1319 (
            .O(N__6972),
            .I(\U712_REG_SM.DS_EN_RNOZ0Z_0 ));
    InMux I__1318 (
            .O(N__6969),
            .I(N__6966));
    LocalMux I__1317 (
            .O(N__6966),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__1316 (
            .O(N__6963),
            .I(N__6959));
    IoInMux I__1315 (
            .O(N__6962),
            .I(N__6956));
    LocalMux I__1314 (
            .O(N__6959),
            .I(N__6953));
    LocalMux I__1313 (
            .O(N__6956),
            .I(N__6950));
    Sp12to4 I__1312 (
            .O(N__6953),
            .I(N__6947));
    IoSpan4Mux I__1311 (
            .O(N__6950),
            .I(N__6944));
    Span12Mux_v I__1310 (
            .O(N__6947),
            .I(N__6941));
    IoSpan4Mux I__1309 (
            .O(N__6944),
            .I(N__6938));
    Span12Mux_h I__1308 (
            .O(N__6941),
            .I(N__6935));
    IoSpan4Mux I__1307 (
            .O(N__6938),
            .I(N__6932));
    Odrv12 I__1306 (
            .O(N__6935),
            .I(C1_c));
    Odrv4 I__1305 (
            .O(N__6932),
            .I(C1_c));
    InMux I__1304 (
            .O(N__6927),
            .I(N__6924));
    LocalMux I__1303 (
            .O(N__6924),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    IoInMux I__1302 (
            .O(N__6921),
            .I(N__6918));
    LocalMux I__1301 (
            .O(N__6918),
            .I(N__6915));
    Span4Mux_s3_v I__1300 (
            .O(N__6915),
            .I(N__6912));
    Span4Mux_v I__1299 (
            .O(N__6912),
            .I(N__6909));
    Sp12to4 I__1298 (
            .O(N__6909),
            .I(N__6906));
    Odrv12 I__1297 (
            .O(N__6906),
            .I(RASn_c));
    InMux I__1296 (
            .O(N__6903),
            .I(N__6893));
    CascadeMux I__1295 (
            .O(N__6902),
            .I(N__6890));
    InMux I__1294 (
            .O(N__6901),
            .I(N__6885));
    InMux I__1293 (
            .O(N__6900),
            .I(N__6885));
    CascadeMux I__1292 (
            .O(N__6899),
            .I(N__6882));
    InMux I__1291 (
            .O(N__6898),
            .I(N__6878));
    InMux I__1290 (
            .O(N__6897),
            .I(N__6875));
    InMux I__1289 (
            .O(N__6896),
            .I(N__6872));
    LocalMux I__1288 (
            .O(N__6893),
            .I(N__6869));
    InMux I__1287 (
            .O(N__6890),
            .I(N__6866));
    LocalMux I__1286 (
            .O(N__6885),
            .I(N__6863));
    InMux I__1285 (
            .O(N__6882),
            .I(N__6858));
    InMux I__1284 (
            .O(N__6881),
            .I(N__6855));
    LocalMux I__1283 (
            .O(N__6878),
            .I(N__6852));
    LocalMux I__1282 (
            .O(N__6875),
            .I(N__6847));
    LocalMux I__1281 (
            .O(N__6872),
            .I(N__6847));
    Span4Mux_h I__1280 (
            .O(N__6869),
            .I(N__6844));
    LocalMux I__1279 (
            .O(N__6866),
            .I(N__6839));
    Span4Mux_h I__1278 (
            .O(N__6863),
            .I(N__6839));
    InMux I__1277 (
            .O(N__6862),
            .I(N__6836));
    InMux I__1276 (
            .O(N__6861),
            .I(N__6833));
    LocalMux I__1275 (
            .O(N__6858),
            .I(N__6824));
    LocalMux I__1274 (
            .O(N__6855),
            .I(N__6824));
    Span4Mux_v I__1273 (
            .O(N__6852),
            .I(N__6824));
    Span4Mux_v I__1272 (
            .O(N__6847),
            .I(N__6824));
    Odrv4 I__1271 (
            .O(N__6844),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1270 (
            .O(N__6839),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1269 (
            .O(N__6836),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1268 (
            .O(N__6833),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1267 (
            .O(N__6824),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1266 (
            .O(N__6813),
            .I(N__6803));
    InMux I__1265 (
            .O(N__6812),
            .I(N__6796));
    InMux I__1264 (
            .O(N__6811),
            .I(N__6796));
    InMux I__1263 (
            .O(N__6810),
            .I(N__6796));
    InMux I__1262 (
            .O(N__6809),
            .I(N__6793));
    CascadeMux I__1261 (
            .O(N__6808),
            .I(N__6786));
    InMux I__1260 (
            .O(N__6807),
            .I(N__6781));
    InMux I__1259 (
            .O(N__6806),
            .I(N__6778));
    LocalMux I__1258 (
            .O(N__6803),
            .I(N__6775));
    LocalMux I__1257 (
            .O(N__6796),
            .I(N__6769));
    LocalMux I__1256 (
            .O(N__6793),
            .I(N__6769));
    InMux I__1255 (
            .O(N__6792),
            .I(N__6762));
    InMux I__1254 (
            .O(N__6791),
            .I(N__6757));
    InMux I__1253 (
            .O(N__6790),
            .I(N__6757));
    InMux I__1252 (
            .O(N__6789),
            .I(N__6754));
    InMux I__1251 (
            .O(N__6786),
            .I(N__6749));
    InMux I__1250 (
            .O(N__6785),
            .I(N__6749));
    InMux I__1249 (
            .O(N__6784),
            .I(N__6746));
    LocalMux I__1248 (
            .O(N__6781),
            .I(N__6743));
    LocalMux I__1247 (
            .O(N__6778),
            .I(N__6740));
    Span4Mux_v I__1246 (
            .O(N__6775),
            .I(N__6737));
    InMux I__1245 (
            .O(N__6774),
            .I(N__6734));
    Span4Mux_h I__1244 (
            .O(N__6769),
            .I(N__6731));
    InMux I__1243 (
            .O(N__6768),
            .I(N__6728));
    InMux I__1242 (
            .O(N__6767),
            .I(N__6721));
    InMux I__1241 (
            .O(N__6766),
            .I(N__6721));
    InMux I__1240 (
            .O(N__6765),
            .I(N__6721));
    LocalMux I__1239 (
            .O(N__6762),
            .I(N__6714));
    LocalMux I__1238 (
            .O(N__6757),
            .I(N__6714));
    LocalMux I__1237 (
            .O(N__6754),
            .I(N__6714));
    LocalMux I__1236 (
            .O(N__6749),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1235 (
            .O(N__6746),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1234 (
            .O(N__6743),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1233 (
            .O(N__6740),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1232 (
            .O(N__6737),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1231 (
            .O(N__6734),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1230 (
            .O(N__6731),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1229 (
            .O(N__6728),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1228 (
            .O(N__6721),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv12 I__1227 (
            .O(N__6714),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    CascadeMux I__1226 (
            .O(N__6693),
            .I(N__6684));
    CascadeMux I__1225 (
            .O(N__6692),
            .I(N__6681));
    InMux I__1224 (
            .O(N__6691),
            .I(N__6675));
    InMux I__1223 (
            .O(N__6690),
            .I(N__6672));
    InMux I__1222 (
            .O(N__6689),
            .I(N__6667));
    InMux I__1221 (
            .O(N__6688),
            .I(N__6667));
    InMux I__1220 (
            .O(N__6687),
            .I(N__6660));
    InMux I__1219 (
            .O(N__6684),
            .I(N__6660));
    InMux I__1218 (
            .O(N__6681),
            .I(N__6660));
    CascadeMux I__1217 (
            .O(N__6680),
            .I(N__6654));
    InMux I__1216 (
            .O(N__6679),
            .I(N__6648));
    InMux I__1215 (
            .O(N__6678),
            .I(N__6645));
    LocalMux I__1214 (
            .O(N__6675),
            .I(N__6642));
    LocalMux I__1213 (
            .O(N__6672),
            .I(N__6639));
    LocalMux I__1212 (
            .O(N__6667),
            .I(N__6634));
    LocalMux I__1211 (
            .O(N__6660),
            .I(N__6634));
    InMux I__1210 (
            .O(N__6659),
            .I(N__6631));
    InMux I__1209 (
            .O(N__6658),
            .I(N__6626));
    InMux I__1208 (
            .O(N__6657),
            .I(N__6626));
    InMux I__1207 (
            .O(N__6654),
            .I(N__6619));
    InMux I__1206 (
            .O(N__6653),
            .I(N__6619));
    InMux I__1205 (
            .O(N__6652),
            .I(N__6619));
    InMux I__1204 (
            .O(N__6651),
            .I(N__6616));
    LocalMux I__1203 (
            .O(N__6648),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1202 (
            .O(N__6645),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1201 (
            .O(N__6642),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1200 (
            .O(N__6639),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1199 (
            .O(N__6634),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1198 (
            .O(N__6631),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1197 (
            .O(N__6626),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1196 (
            .O(N__6619),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1195 (
            .O(N__6616),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__1194 (
            .O(N__6597),
            .I(N__6591));
    CascadeMux I__1193 (
            .O(N__6596),
            .I(N__6588));
    InMux I__1192 (
            .O(N__6595),
            .I(N__6583));
    InMux I__1191 (
            .O(N__6594),
            .I(N__6580));
    InMux I__1190 (
            .O(N__6591),
            .I(N__6572));
    InMux I__1189 (
            .O(N__6588),
            .I(N__6572));
    CascadeMux I__1188 (
            .O(N__6587),
            .I(N__6568));
    InMux I__1187 (
            .O(N__6586),
            .I(N__6562));
    LocalMux I__1186 (
            .O(N__6583),
            .I(N__6557));
    LocalMux I__1185 (
            .O(N__6580),
            .I(N__6557));
    InMux I__1184 (
            .O(N__6579),
            .I(N__6554));
    InMux I__1183 (
            .O(N__6578),
            .I(N__6551));
    CascadeMux I__1182 (
            .O(N__6577),
            .I(N__6548));
    LocalMux I__1181 (
            .O(N__6572),
            .I(N__6543));
    InMux I__1180 (
            .O(N__6571),
            .I(N__6540));
    InMux I__1179 (
            .O(N__6568),
            .I(N__6533));
    InMux I__1178 (
            .O(N__6567),
            .I(N__6533));
    InMux I__1177 (
            .O(N__6566),
            .I(N__6533));
    InMux I__1176 (
            .O(N__6565),
            .I(N__6530));
    LocalMux I__1175 (
            .O(N__6562),
            .I(N__6527));
    Span4Mux_v I__1174 (
            .O(N__6557),
            .I(N__6520));
    LocalMux I__1173 (
            .O(N__6554),
            .I(N__6520));
    LocalMux I__1172 (
            .O(N__6551),
            .I(N__6520));
    InMux I__1171 (
            .O(N__6548),
            .I(N__6513));
    InMux I__1170 (
            .O(N__6547),
            .I(N__6513));
    InMux I__1169 (
            .O(N__6546),
            .I(N__6513));
    Odrv4 I__1168 (
            .O(N__6543),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1167 (
            .O(N__6540),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1166 (
            .O(N__6533),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1165 (
            .O(N__6530),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1164 (
            .O(N__6527),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1163 (
            .O(N__6520),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1162 (
            .O(N__6513),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1161 (
            .O(N__6498),
            .I(N__6495));
    LocalMux I__1160 (
            .O(N__6495),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_a2_0_0 ));
    InMux I__1159 (
            .O(N__6492),
            .I(N__6489));
    LocalMux I__1158 (
            .O(N__6489),
            .I(N__6486));
    Span4Mux_v I__1157 (
            .O(N__6486),
            .I(N__6482));
    IoInMux I__1156 (
            .O(N__6485),
            .I(N__6479));
    Span4Mux_h I__1155 (
            .O(N__6482),
            .I(N__6476));
    LocalMux I__1154 (
            .O(N__6479),
            .I(N__6473));
    Sp12to4 I__1153 (
            .O(N__6476),
            .I(N__6470));
    IoSpan4Mux I__1152 (
            .O(N__6473),
            .I(N__6467));
    Odrv12 I__1151 (
            .O(N__6470),
            .I(RAMENn_c));
    Odrv4 I__1150 (
            .O(N__6467),
            .I(RAMENn_c));
    CascadeMux I__1149 (
            .O(N__6462),
            .I(\U712_CHIP_RAM.N_492_cascade_ ));
    InMux I__1148 (
            .O(N__6459),
            .I(N__6454));
    InMux I__1147 (
            .O(N__6458),
            .I(N__6449));
    InMux I__1146 (
            .O(N__6457),
            .I(N__6449));
    LocalMux I__1145 (
            .O(N__6454),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__1144 (
            .O(N__6449),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__1143 (
            .O(N__6444),
            .I(\U712_REG_SM.STATE_COUNT_srsts_i_0_0_a2_0_0_0_cascade_ ));
    InMux I__1142 (
            .O(N__6441),
            .I(N__6438));
    LocalMux I__1141 (
            .O(N__6438),
            .I(\U712_REG_SM.N_374 ));
    InMux I__1140 (
            .O(N__6435),
            .I(N__6432));
    LocalMux I__1139 (
            .O(N__6432),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_a2_1_0 ));
    IoInMux I__1138 (
            .O(N__6429),
            .I(N__6426));
    LocalMux I__1137 (
            .O(N__6426),
            .I(N__6423));
    Span12Mux_s4_v I__1136 (
            .O(N__6423),
            .I(N__6419));
    InMux I__1135 (
            .O(N__6422),
            .I(N__6416));
    Span12Mux_h I__1134 (
            .O(N__6419),
            .I(N__6413));
    LocalMux I__1133 (
            .O(N__6416),
            .I(N__6410));
    Span12Mux_v I__1132 (
            .O(N__6413),
            .I(N__6407));
    Span12Mux_h I__1131 (
            .O(N__6410),
            .I(N__6404));
    Odrv12 I__1130 (
            .O(N__6407),
            .I(A_c_9));
    Odrv12 I__1129 (
            .O(N__6404),
            .I(A_c_9));
    InMux I__1128 (
            .O(N__6399),
            .I(N__6396));
    LocalMux I__1127 (
            .O(N__6396),
            .I(N__6393));
    Sp12to4 I__1126 (
            .O(N__6393),
            .I(N__6390));
    Span12Mux_v I__1125 (
            .O(N__6390),
            .I(N__6387));
    Span12Mux_h I__1124 (
            .O(N__6387),
            .I(N__6384));
    Odrv12 I__1123 (
            .O(N__6384),
            .I(A_c_2));
    InMux I__1122 (
            .O(N__6381),
            .I(N__6378));
    LocalMux I__1121 (
            .O(N__6378),
            .I(N__6374));
    InMux I__1120 (
            .O(N__6377),
            .I(N__6371));
    Span4Mux_h I__1119 (
            .O(N__6374),
            .I(N__6368));
    LocalMux I__1118 (
            .O(N__6371),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    Odrv4 I__1117 (
            .O(N__6368),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__1116 (
            .O(N__6363),
            .I(N__6360));
    LocalMux I__1115 (
            .O(N__6360),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ));
    InMux I__1114 (
            .O(N__6357),
            .I(N__6354));
    LocalMux I__1113 (
            .O(N__6354),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    InMux I__1112 (
            .O(N__6351),
            .I(N__6347));
    InMux I__1111 (
            .O(N__6350),
            .I(N__6344));
    LocalMux I__1110 (
            .O(N__6347),
            .I(N__6341));
    LocalMux I__1109 (
            .O(N__6344),
            .I(N__6337));
    Span4Mux_h I__1108 (
            .O(N__6341),
            .I(N__6334));
    InMux I__1107 (
            .O(N__6340),
            .I(N__6331));
    Odrv4 I__1106 (
            .O(N__6337),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    Odrv4 I__1105 (
            .O(N__6334),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__1104 (
            .O(N__6331),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    CascadeMux I__1103 (
            .O(N__6324),
            .I(N__6320));
    CascadeMux I__1102 (
            .O(N__6323),
            .I(N__6317));
    InMux I__1101 (
            .O(N__6320),
            .I(N__6314));
    InMux I__1100 (
            .O(N__6317),
            .I(N__6311));
    LocalMux I__1099 (
            .O(N__6314),
            .I(N__6308));
    LocalMux I__1098 (
            .O(N__6311),
            .I(N__6305));
    Span4Mux_v I__1097 (
            .O(N__6308),
            .I(N__6302));
    Span4Mux_h I__1096 (
            .O(N__6305),
            .I(N__6299));
    Odrv4 I__1095 (
            .O(N__6302),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    Odrv4 I__1094 (
            .O(N__6299),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    InMux I__1093 (
            .O(N__6294),
            .I(N__6290));
    InMux I__1092 (
            .O(N__6293),
            .I(N__6287));
    LocalMux I__1091 (
            .O(N__6290),
            .I(N__6281));
    LocalMux I__1090 (
            .O(N__6287),
            .I(N__6281));
    InMux I__1089 (
            .O(N__6286),
            .I(N__6278));
    Span4Mux_h I__1088 (
            .O(N__6281),
            .I(N__6274));
    LocalMux I__1087 (
            .O(N__6278),
            .I(N__6271));
    InMux I__1086 (
            .O(N__6277),
            .I(N__6268));
    Odrv4 I__1085 (
            .O(N__6274),
            .I(\U712_CHIP_RAM.N_567 ));
    Odrv4 I__1084 (
            .O(N__6271),
            .I(\U712_CHIP_RAM.N_567 ));
    LocalMux I__1083 (
            .O(N__6268),
            .I(\U712_CHIP_RAM.N_567 ));
    InMux I__1082 (
            .O(N__6261),
            .I(N__6256));
    InMux I__1081 (
            .O(N__6260),
            .I(N__6251));
    InMux I__1080 (
            .O(N__6259),
            .I(N__6251));
    LocalMux I__1079 (
            .O(N__6256),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1078 (
            .O(N__6251),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    CascadeMux I__1077 (
            .O(N__6246),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_1_cascade_ ));
    InMux I__1076 (
            .O(N__6243),
            .I(N__6240));
    LocalMux I__1075 (
            .O(N__6240),
            .I(N__6235));
    InMux I__1074 (
            .O(N__6239),
            .I(N__6232));
    InMux I__1073 (
            .O(N__6238),
            .I(N__6229));
    Span4Mux_h I__1072 (
            .O(N__6235),
            .I(N__6219));
    LocalMux I__1071 (
            .O(N__6232),
            .I(N__6219));
    LocalMux I__1070 (
            .O(N__6229),
            .I(N__6219));
    InMux I__1069 (
            .O(N__6228),
            .I(N__6216));
    InMux I__1068 (
            .O(N__6227),
            .I(N__6213));
    InMux I__1067 (
            .O(N__6226),
            .I(N__6210));
    Odrv4 I__1066 (
            .O(N__6219),
            .I(\U712_CHIP_RAM.N_562 ));
    LocalMux I__1065 (
            .O(N__6216),
            .I(\U712_CHIP_RAM.N_562 ));
    LocalMux I__1064 (
            .O(N__6213),
            .I(\U712_CHIP_RAM.N_562 ));
    LocalMux I__1063 (
            .O(N__6210),
            .I(\U712_CHIP_RAM.N_562 ));
    InMux I__1062 (
            .O(N__6201),
            .I(N__6197));
    InMux I__1061 (
            .O(N__6200),
            .I(N__6194));
    LocalMux I__1060 (
            .O(N__6197),
            .I(N__6191));
    LocalMux I__1059 (
            .O(N__6194),
            .I(\U712_CHIP_RAM.N_502 ));
    Odrv4 I__1058 (
            .O(N__6191),
            .I(\U712_CHIP_RAM.N_502 ));
    CascadeMux I__1057 (
            .O(N__6186),
            .I(N__6182));
    CascadeMux I__1056 (
            .O(N__6185),
            .I(N__6179));
    InMux I__1055 (
            .O(N__6182),
            .I(N__6174));
    InMux I__1054 (
            .O(N__6179),
            .I(N__6171));
    CascadeMux I__1053 (
            .O(N__6178),
            .I(N__6168));
    InMux I__1052 (
            .O(N__6177),
            .I(N__6165));
    LocalMux I__1051 (
            .O(N__6174),
            .I(N__6160));
    LocalMux I__1050 (
            .O(N__6171),
            .I(N__6157));
    InMux I__1049 (
            .O(N__6168),
            .I(N__6154));
    LocalMux I__1048 (
            .O(N__6165),
            .I(N__6151));
    InMux I__1047 (
            .O(N__6164),
            .I(N__6148));
    InMux I__1046 (
            .O(N__6163),
            .I(N__6141));
    Span4Mux_v I__1045 (
            .O(N__6160),
            .I(N__6136));
    Span4Mux_v I__1044 (
            .O(N__6157),
            .I(N__6136));
    LocalMux I__1043 (
            .O(N__6154),
            .I(N__6129));
    Span4Mux_v I__1042 (
            .O(N__6151),
            .I(N__6129));
    LocalMux I__1041 (
            .O(N__6148),
            .I(N__6129));
    InMux I__1040 (
            .O(N__6147),
            .I(N__6126));
    InMux I__1039 (
            .O(N__6146),
            .I(N__6123));
    InMux I__1038 (
            .O(N__6145),
            .I(N__6120));
    InMux I__1037 (
            .O(N__6144),
            .I(N__6117));
    LocalMux I__1036 (
            .O(N__6141),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    Odrv4 I__1035 (
            .O(N__6136),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    Odrv4 I__1034 (
            .O(N__6129),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1033 (
            .O(N__6126),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1032 (
            .O(N__6123),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1031 (
            .O(N__6120),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1030 (
            .O(N__6117),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__1029 (
            .O(N__6102),
            .I(N__6098));
    InMux I__1028 (
            .O(N__6101),
            .I(N__6095));
    LocalMux I__1027 (
            .O(N__6098),
            .I(N__6089));
    LocalMux I__1026 (
            .O(N__6095),
            .I(N__6086));
    InMux I__1025 (
            .O(N__6094),
            .I(N__6083));
    CascadeMux I__1024 (
            .O(N__6093),
            .I(N__6077));
    InMux I__1023 (
            .O(N__6092),
            .I(N__6072));
    Span4Mux_h I__1022 (
            .O(N__6089),
            .I(N__6069));
    Span4Mux_h I__1021 (
            .O(N__6086),
            .I(N__6064));
    LocalMux I__1020 (
            .O(N__6083),
            .I(N__6064));
    InMux I__1019 (
            .O(N__6082),
            .I(N__6061));
    InMux I__1018 (
            .O(N__6081),
            .I(N__6058));
    InMux I__1017 (
            .O(N__6080),
            .I(N__6055));
    InMux I__1016 (
            .O(N__6077),
            .I(N__6052));
    InMux I__1015 (
            .O(N__6076),
            .I(N__6047));
    InMux I__1014 (
            .O(N__6075),
            .I(N__6047));
    LocalMux I__1013 (
            .O(N__6072),
            .I(\U712_CHIP_RAM.N_545 ));
    Odrv4 I__1012 (
            .O(N__6069),
            .I(\U712_CHIP_RAM.N_545 ));
    Odrv4 I__1011 (
            .O(N__6064),
            .I(\U712_CHIP_RAM.N_545 ));
    LocalMux I__1010 (
            .O(N__6061),
            .I(\U712_CHIP_RAM.N_545 ));
    LocalMux I__1009 (
            .O(N__6058),
            .I(\U712_CHIP_RAM.N_545 ));
    LocalMux I__1008 (
            .O(N__6055),
            .I(\U712_CHIP_RAM.N_545 ));
    LocalMux I__1007 (
            .O(N__6052),
            .I(\U712_CHIP_RAM.N_545 ));
    LocalMux I__1006 (
            .O(N__6047),
            .I(\U712_CHIP_RAM.N_545 ));
    InMux I__1005 (
            .O(N__6030),
            .I(N__6023));
    InMux I__1004 (
            .O(N__6029),
            .I(N__6023));
    InMux I__1003 (
            .O(N__6028),
            .I(N__6019));
    LocalMux I__1002 (
            .O(N__6023),
            .I(N__6016));
    InMux I__1001 (
            .O(N__6022),
            .I(N__6013));
    LocalMux I__1000 (
            .O(N__6019),
            .I(\U712_CHIP_RAM.N_572 ));
    Odrv12 I__999 (
            .O(N__6016),
            .I(\U712_CHIP_RAM.N_572 ));
    LocalMux I__998 (
            .O(N__6013),
            .I(\U712_CHIP_RAM.N_572 ));
    CascadeMux I__997 (
            .O(N__6006),
            .I(\U712_CHIP_RAM.N_518_cascade_ ));
    InMux I__996 (
            .O(N__6003),
            .I(N__5999));
    CascadeMux I__995 (
            .O(N__6002),
            .I(N__5996));
    LocalMux I__994 (
            .O(N__5999),
            .I(N__5993));
    InMux I__993 (
            .O(N__5996),
            .I(N__5985));
    Span4Mux_v I__992 (
            .O(N__5993),
            .I(N__5982));
    InMux I__991 (
            .O(N__5992),
            .I(N__5979));
    InMux I__990 (
            .O(N__5991),
            .I(N__5974));
    InMux I__989 (
            .O(N__5990),
            .I(N__5974));
    InMux I__988 (
            .O(N__5989),
            .I(N__5969));
    InMux I__987 (
            .O(N__5988),
            .I(N__5969));
    LocalMux I__986 (
            .O(N__5985),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__985 (
            .O(N__5982),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__984 (
            .O(N__5979),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__983 (
            .O(N__5974),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__982 (
            .O(N__5969),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    InMux I__981 (
            .O(N__5958),
            .I(N__5955));
    LocalMux I__980 (
            .O(N__5955),
            .I(N__5952));
    Odrv4 I__979 (
            .O(N__5952),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0 ));
    InMux I__978 (
            .O(N__5949),
            .I(N__5946));
    LocalMux I__977 (
            .O(N__5946),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ));
    InMux I__976 (
            .O(N__5943),
            .I(N__5940));
    LocalMux I__975 (
            .O(N__5940),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    CascadeMux I__974 (
            .O(N__5937),
            .I(\U712_CHIP_RAM.N_379_cascade_ ));
    InMux I__973 (
            .O(N__5934),
            .I(N__5931));
    LocalMux I__972 (
            .O(N__5931),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    InMux I__971 (
            .O(N__5928),
            .I(N__5925));
    LocalMux I__970 (
            .O(N__5925),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    SRMux I__969 (
            .O(N__5922),
            .I(N__5919));
    LocalMux I__968 (
            .O(N__5919),
            .I(N__5916));
    Odrv12 I__967 (
            .O(N__5916),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    CascadeMux I__966 (
            .O(N__5913),
            .I(\U712_CHIP_RAM.REFRESH_RST_cascade_ ));
    InMux I__965 (
            .O(N__5910),
            .I(N__5907));
    LocalMux I__964 (
            .O(N__5907),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i ));
    IoInMux I__963 (
            .O(N__5904),
            .I(N__5901));
    LocalMux I__962 (
            .O(N__5901),
            .I(N__5898));
    IoSpan4Mux I__961 (
            .O(N__5898),
            .I(N__5895));
    Span4Mux_s2_v I__960 (
            .O(N__5895),
            .I(N__5892));
    Sp12to4 I__959 (
            .O(N__5892),
            .I(N__5888));
    InMux I__958 (
            .O(N__5891),
            .I(N__5885));
    Span12Mux_s8_v I__957 (
            .O(N__5888),
            .I(N__5882));
    LocalMux I__956 (
            .O(N__5885),
            .I(N__5879));
    Span12Mux_v I__955 (
            .O(N__5882),
            .I(N__5876));
    Span4Mux_v I__954 (
            .O(N__5879),
            .I(N__5873));
    Span12Mux_h I__953 (
            .O(N__5876),
            .I(N__5868));
    Sp12to4 I__952 (
            .O(N__5873),
            .I(N__5868));
    Span12Mux_h I__951 (
            .O(N__5868),
            .I(N__5865));
    Odrv12 I__950 (
            .O(N__5865),
            .I(A_c_11));
    InMux I__949 (
            .O(N__5862),
            .I(N__5859));
    LocalMux I__948 (
            .O(N__5859),
            .I(N__5856));
    Span4Mux_v I__947 (
            .O(N__5856),
            .I(N__5853));
    Span4Mux_v I__946 (
            .O(N__5853),
            .I(N__5850));
    Sp12to4 I__945 (
            .O(N__5850),
            .I(N__5847));
    Span12Mux_h I__944 (
            .O(N__5847),
            .I(N__5844));
    Odrv12 I__943 (
            .O(N__5844),
            .I(A_c_4));
    InMux I__942 (
            .O(N__5841),
            .I(N__5838));
    LocalMux I__941 (
            .O(N__5838),
            .I(\U712_CHIP_RAM.N_517 ));
    InMux I__940 (
            .O(N__5835),
            .I(N__5830));
    InMux I__939 (
            .O(N__5834),
            .I(N__5825));
    InMux I__938 (
            .O(N__5833),
            .I(N__5825));
    LocalMux I__937 (
            .O(N__5830),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    LocalMux I__936 (
            .O(N__5825),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    IoInMux I__935 (
            .O(N__5820),
            .I(N__5817));
    LocalMux I__934 (
            .O(N__5817),
            .I(N__5813));
    IoInMux I__933 (
            .O(N__5816),
            .I(N__5810));
    Span4Mux_s0_v I__932 (
            .O(N__5813),
            .I(N__5807));
    LocalMux I__931 (
            .O(N__5810),
            .I(N__5804));
    Sp12to4 I__930 (
            .O(N__5807),
            .I(N__5801));
    IoSpan4Mux I__929 (
            .O(N__5804),
            .I(N__5798));
    Span12Mux_s11_h I__928 (
            .O(N__5801),
            .I(N__5795));
    Sp12to4 I__927 (
            .O(N__5798),
            .I(N__5792));
    Span12Mux_v I__926 (
            .O(N__5795),
            .I(N__5786));
    Span12Mux_v I__925 (
            .O(N__5792),
            .I(N__5786));
    InMux I__924 (
            .O(N__5791),
            .I(N__5783));
    Odrv12 I__923 (
            .O(N__5786),
            .I(ASn_c));
    LocalMux I__922 (
            .O(N__5783),
            .I(ASn_c));
    CascadeMux I__921 (
            .O(N__5778),
            .I(N__5774));
    InMux I__920 (
            .O(N__5777),
            .I(N__5769));
    InMux I__919 (
            .O(N__5774),
            .I(N__5766));
    InMux I__918 (
            .O(N__5773),
            .I(N__5763));
    InMux I__917 (
            .O(N__5772),
            .I(N__5760));
    LocalMux I__916 (
            .O(N__5769),
            .I(N__5757));
    LocalMux I__915 (
            .O(N__5766),
            .I(REG_TACK));
    LocalMux I__914 (
            .O(N__5763),
            .I(REG_TACK));
    LocalMux I__913 (
            .O(N__5760),
            .I(REG_TACK));
    Odrv4 I__912 (
            .O(N__5757),
            .I(REG_TACK));
    InMux I__911 (
            .O(N__5748),
            .I(N__5744));
    InMux I__910 (
            .O(N__5747),
            .I(N__5741));
    LocalMux I__909 (
            .O(N__5744),
            .I(N__5738));
    LocalMux I__908 (
            .O(N__5741),
            .I(N__5735));
    Span4Mux_v I__907 (
            .O(N__5738),
            .I(N__5732));
    Span4Mux_v I__906 (
            .O(N__5735),
            .I(N__5729));
    Sp12to4 I__905 (
            .O(N__5732),
            .I(N__5726));
    Span4Mux_h I__904 (
            .O(N__5729),
            .I(N__5723));
    Span12Mux_h I__903 (
            .O(N__5726),
            .I(N__5718));
    Sp12to4 I__902 (
            .O(N__5723),
            .I(N__5718));
    Odrv12 I__901 (
            .O(N__5718),
            .I(AWEn_c));
    InMux I__900 (
            .O(N__5715),
            .I(N__5711));
    InMux I__899 (
            .O(N__5714),
            .I(N__5708));
    LocalMux I__898 (
            .O(N__5711),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    LocalMux I__897 (
            .O(N__5708),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    IoInMux I__896 (
            .O(N__5703),
            .I(N__5700));
    LocalMux I__895 (
            .O(N__5700),
            .I(N__5697));
    IoSpan4Mux I__894 (
            .O(N__5697),
            .I(N__5694));
    Span4Mux_s3_v I__893 (
            .O(N__5694),
            .I(N__5691));
    Span4Mux_v I__892 (
            .O(N__5691),
            .I(N__5688));
    Sp12to4 I__891 (
            .O(N__5688),
            .I(N__5685));
    Span12Mux_v I__890 (
            .O(N__5685),
            .I(N__5681));
    InMux I__889 (
            .O(N__5684),
            .I(N__5678));
    Odrv12 I__888 (
            .O(N__5681),
            .I(DBDIR_c));
    LocalMux I__887 (
            .O(N__5678),
            .I(DBDIR_c));
    InMux I__886 (
            .O(N__5673),
            .I(N__5670));
    LocalMux I__885 (
            .O(N__5670),
            .I(N__5667));
    Span4Mux_v I__884 (
            .O(N__5667),
            .I(N__5664));
    Odrv4 I__883 (
            .O(N__5664),
            .I(\U712_REG_SM.N_447 ));
    CascadeMux I__882 (
            .O(N__5661),
            .I(\U712_REG_SM.N_447_cascade_ ));
    InMux I__881 (
            .O(N__5658),
            .I(N__5655));
    LocalMux I__880 (
            .O(N__5655),
            .I(\U712_REG_SM.REG_TACK_RNOZ0Z_0 ));
    InMux I__879 (
            .O(N__5652),
            .I(N__5649));
    LocalMux I__878 (
            .O(N__5649),
            .I(\U712_REG_SM.N_478 ));
    IoInMux I__877 (
            .O(N__5646),
            .I(N__5643));
    LocalMux I__876 (
            .O(N__5643),
            .I(N__5640));
    IoSpan4Mux I__875 (
            .O(N__5640),
            .I(N__5637));
    Span4Mux_s2_h I__874 (
            .O(N__5637),
            .I(N__5634));
    Sp12to4 I__873 (
            .O(N__5634),
            .I(N__5631));
    Span12Mux_s11_h I__872 (
            .O(N__5631),
            .I(N__5628));
    Span12Mux_v I__871 (
            .O(N__5628),
            .I(N__5625));
    Odrv12 I__870 (
            .O(N__5625),
            .I(CMA_c_5));
    InMux I__869 (
            .O(N__5622),
            .I(N__5619));
    LocalMux I__868 (
            .O(N__5619),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__867 (
            .O(N__5616),
            .I(N__5613));
    LocalMux I__866 (
            .O(N__5613),
            .I(N__5610));
    Span4Mux_s3_h I__865 (
            .O(N__5610),
            .I(N__5607));
    Sp12to4 I__864 (
            .O(N__5607),
            .I(N__5604));
    Span12Mux_v I__863 (
            .O(N__5604),
            .I(N__5601));
    Span12Mux_h I__862 (
            .O(N__5601),
            .I(N__5598));
    Odrv12 I__861 (
            .O(N__5598),
            .I(CMA_c_7));
    CascadeMux I__860 (
            .O(N__5595),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_ ));
    CEMux I__859 (
            .O(N__5592),
            .I(N__5589));
    LocalMux I__858 (
            .O(N__5589),
            .I(N__5586));
    Span4Mux_h I__857 (
            .O(N__5586),
            .I(N__5583));
    Odrv4 I__856 (
            .O(N__5583),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_1 ));
    InMux I__855 (
            .O(N__5580),
            .I(N__5576));
    InMux I__854 (
            .O(N__5579),
            .I(N__5573));
    LocalMux I__853 (
            .O(N__5576),
            .I(\U712_CHIP_RAM.N_666 ));
    LocalMux I__852 (
            .O(N__5573),
            .I(\U712_CHIP_RAM.N_666 ));
    InMux I__851 (
            .O(N__5568),
            .I(N__5565));
    LocalMux I__850 (
            .O(N__5565),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0 ));
    CascadeMux I__849 (
            .O(N__5562),
            .I(N__5559));
    InMux I__848 (
            .O(N__5559),
            .I(N__5552));
    InMux I__847 (
            .O(N__5558),
            .I(N__5549));
    InMux I__846 (
            .O(N__5557),
            .I(N__5545));
    InMux I__845 (
            .O(N__5556),
            .I(N__5540));
    InMux I__844 (
            .O(N__5555),
            .I(N__5540));
    LocalMux I__843 (
            .O(N__5552),
            .I(N__5535));
    LocalMux I__842 (
            .O(N__5549),
            .I(N__5535));
    InMux I__841 (
            .O(N__5548),
            .I(N__5532));
    LocalMux I__840 (
            .O(N__5545),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__839 (
            .O(N__5540),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__838 (
            .O(N__5535),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__837 (
            .O(N__5532),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__836 (
            .O(N__5523),
            .I(N__5519));
    InMux I__835 (
            .O(N__5522),
            .I(N__5513));
    LocalMux I__834 (
            .O(N__5519),
            .I(N__5510));
    InMux I__833 (
            .O(N__5518),
            .I(N__5507));
    InMux I__832 (
            .O(N__5517),
            .I(N__5504));
    CascadeMux I__831 (
            .O(N__5516),
            .I(N__5500));
    LocalMux I__830 (
            .O(N__5513),
            .I(N__5497));
    Span4Mux_v I__829 (
            .O(N__5510),
            .I(N__5494));
    LocalMux I__828 (
            .O(N__5507),
            .I(N__5489));
    LocalMux I__827 (
            .O(N__5504),
            .I(N__5489));
    InMux I__826 (
            .O(N__5503),
            .I(N__5486));
    InMux I__825 (
            .O(N__5500),
            .I(N__5483));
    Span4Mux_v I__824 (
            .O(N__5497),
            .I(N__5480));
    Odrv4 I__823 (
            .O(N__5494),
            .I(\U712_CHIP_RAM.N_557 ));
    Odrv4 I__822 (
            .O(N__5489),
            .I(\U712_CHIP_RAM.N_557 ));
    LocalMux I__821 (
            .O(N__5486),
            .I(\U712_CHIP_RAM.N_557 ));
    LocalMux I__820 (
            .O(N__5483),
            .I(\U712_CHIP_RAM.N_557 ));
    Odrv4 I__819 (
            .O(N__5480),
            .I(\U712_CHIP_RAM.N_557 ));
    InMux I__818 (
            .O(N__5469),
            .I(N__5466));
    LocalMux I__817 (
            .O(N__5466),
            .I(\U712_CHIP_RAM.N_393 ));
    InMux I__816 (
            .O(N__5463),
            .I(N__5459));
    InMux I__815 (
            .O(N__5462),
            .I(N__5456));
    LocalMux I__814 (
            .O(N__5459),
            .I(N__5453));
    LocalMux I__813 (
            .O(N__5456),
            .I(N__5450));
    Span4Mux_h I__812 (
            .O(N__5453),
            .I(N__5445));
    Span4Mux_h I__811 (
            .O(N__5450),
            .I(N__5445));
    Odrv4 I__810 (
            .O(N__5445),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_0_a2_0 ));
    CascadeMux I__809 (
            .O(N__5442),
            .I(\U712_CHIP_RAM.N_557_cascade_ ));
    CascadeMux I__808 (
            .O(N__5439),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_ ));
    InMux I__807 (
            .O(N__5436),
            .I(N__5433));
    LocalMux I__806 (
            .O(N__5433),
            .I(N__5430));
    Odrv4 I__805 (
            .O(N__5430),
            .I(\U712_CHIP_RAM.N_31 ));
    IoInMux I__804 (
            .O(N__5427),
            .I(N__5424));
    LocalMux I__803 (
            .O(N__5424),
            .I(N__5421));
    Span4Mux_s1_v I__802 (
            .O(N__5421),
            .I(N__5418));
    Sp12to4 I__801 (
            .O(N__5418),
            .I(N__5415));
    Span12Mux_h I__800 (
            .O(N__5415),
            .I(N__5412));
    Span12Mux_v I__799 (
            .O(N__5412),
            .I(N__5408));
    InMux I__798 (
            .O(N__5411),
            .I(N__5405));
    Odrv12 I__797 (
            .O(N__5408),
            .I(LATCH_CLK_c));
    LocalMux I__796 (
            .O(N__5405),
            .I(LATCH_CLK_c));
    CascadeMux I__795 (
            .O(N__5400),
            .I(N__5397));
    InMux I__794 (
            .O(N__5397),
            .I(N__5390));
    InMux I__793 (
            .O(N__5396),
            .I(N__5387));
    InMux I__792 (
            .O(N__5395),
            .I(N__5381));
    InMux I__791 (
            .O(N__5394),
            .I(N__5381));
    InMux I__790 (
            .O(N__5393),
            .I(N__5373));
    LocalMux I__789 (
            .O(N__5390),
            .I(N__5368));
    LocalMux I__788 (
            .O(N__5387),
            .I(N__5368));
    InMux I__787 (
            .O(N__5386),
            .I(N__5365));
    LocalMux I__786 (
            .O(N__5381),
            .I(N__5362));
    InMux I__785 (
            .O(N__5380),
            .I(N__5359));
    InMux I__784 (
            .O(N__5379),
            .I(N__5354));
    InMux I__783 (
            .O(N__5378),
            .I(N__5354));
    InMux I__782 (
            .O(N__5377),
            .I(N__5349));
    InMux I__781 (
            .O(N__5376),
            .I(N__5349));
    LocalMux I__780 (
            .O(N__5373),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__779 (
            .O(N__5368),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__778 (
            .O(N__5365),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__777 (
            .O(N__5362),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__776 (
            .O(N__5359),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__775 (
            .O(N__5354),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__774 (
            .O(N__5349),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__773 (
            .O(N__5334),
            .I(N__5331));
    LocalMux I__772 (
            .O(N__5331),
            .I(N__5327));
    InMux I__771 (
            .O(N__5330),
            .I(N__5324));
    Odrv12 I__770 (
            .O(N__5327),
            .I(\U712_CHIP_RAM.N_566 ));
    LocalMux I__769 (
            .O(N__5324),
            .I(\U712_CHIP_RAM.N_566 ));
    CascadeMux I__768 (
            .O(N__5319),
            .I(N__5314));
    CascadeMux I__767 (
            .O(N__5318),
            .I(N__5311));
    InMux I__766 (
            .O(N__5317),
            .I(N__5307));
    InMux I__765 (
            .O(N__5314),
            .I(N__5302));
    InMux I__764 (
            .O(N__5311),
            .I(N__5302));
    InMux I__763 (
            .O(N__5310),
            .I(N__5299));
    LocalMux I__762 (
            .O(N__5307),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__761 (
            .O(N__5302),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__760 (
            .O(N__5299),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    IoInMux I__759 (
            .O(N__5292),
            .I(N__5288));
    IoInMux I__758 (
            .O(N__5291),
            .I(N__5285));
    LocalMux I__757 (
            .O(N__5288),
            .I(N__5282));
    LocalMux I__756 (
            .O(N__5285),
            .I(N__5279));
    IoSpan4Mux I__755 (
            .O(N__5282),
            .I(N__5276));
    IoSpan4Mux I__754 (
            .O(N__5279),
            .I(N__5273));
    Sp12to4 I__753 (
            .O(N__5276),
            .I(N__5269));
    Span4Mux_s2_h I__752 (
            .O(N__5273),
            .I(N__5266));
    InMux I__751 (
            .O(N__5272),
            .I(N__5263));
    Span12Mux_s7_v I__750 (
            .O(N__5269),
            .I(N__5260));
    Sp12to4 I__749 (
            .O(N__5266),
            .I(N__5257));
    LocalMux I__748 (
            .O(N__5263),
            .I(N__5254));
    Span12Mux_v I__747 (
            .O(N__5260),
            .I(N__5250));
    Span12Mux_h I__746 (
            .O(N__5257),
            .I(N__5247));
    Span4Mux_h I__745 (
            .O(N__5254),
            .I(N__5244));
    InMux I__744 (
            .O(N__5253),
            .I(N__5241));
    Odrv12 I__743 (
            .O(N__5250),
            .I(TACK_OUTn));
    Odrv12 I__742 (
            .O(N__5247),
            .I(TACK_OUTn));
    Odrv4 I__741 (
            .O(N__5244),
            .I(TACK_OUTn));
    LocalMux I__740 (
            .O(N__5241),
            .I(TACK_OUTn));
    CascadeMux I__739 (
            .O(N__5232),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ));
    InMux I__738 (
            .O(N__5229),
            .I(N__5226));
    LocalMux I__737 (
            .O(N__5226),
            .I(N__5223));
    Span12Mux_v I__736 (
            .O(N__5223),
            .I(N__5220));
    Span12Mux_h I__735 (
            .O(N__5220),
            .I(N__5217));
    Odrv12 I__734 (
            .O(N__5217),
            .I(A_c_20));
    CascadeMux I__733 (
            .O(N__5214),
            .I(\U712_CHIP_RAM.N_506_cascade_ ));
    InMux I__732 (
            .O(N__5211),
            .I(N__5207));
    InMux I__731 (
            .O(N__5210),
            .I(N__5204));
    LocalMux I__730 (
            .O(N__5207),
            .I(N__5201));
    LocalMux I__729 (
            .O(N__5204),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    Odrv12 I__728 (
            .O(N__5201),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    InMux I__727 (
            .O(N__5196),
            .I(N__5193));
    LocalMux I__726 (
            .O(N__5193),
            .I(N__5190));
    Span4Mux_v I__725 (
            .O(N__5190),
            .I(N__5187));
    Odrv4 I__724 (
            .O(N__5187),
            .I(\U712_CHIP_RAM.N_375 ));
    InMux I__723 (
            .O(N__5184),
            .I(N__5177));
    InMux I__722 (
            .O(N__5183),
            .I(N__5172));
    InMux I__721 (
            .O(N__5182),
            .I(N__5172));
    InMux I__720 (
            .O(N__5181),
            .I(N__5169));
    InMux I__719 (
            .O(N__5180),
            .I(N__5166));
    LocalMux I__718 (
            .O(N__5177),
            .I(\U712_CHIP_RAM.N_547 ));
    LocalMux I__717 (
            .O(N__5172),
            .I(\U712_CHIP_RAM.N_547 ));
    LocalMux I__716 (
            .O(N__5169),
            .I(\U712_CHIP_RAM.N_547 ));
    LocalMux I__715 (
            .O(N__5166),
            .I(\U712_CHIP_RAM.N_547 ));
    InMux I__714 (
            .O(N__5157),
            .I(N__5154));
    LocalMux I__713 (
            .O(N__5154),
            .I(N__5149));
    CascadeMux I__712 (
            .O(N__5153),
            .I(N__5146));
    InMux I__711 (
            .O(N__5152),
            .I(N__5142));
    Span4Mux_h I__710 (
            .O(N__5149),
            .I(N__5139));
    InMux I__709 (
            .O(N__5146),
            .I(N__5136));
    InMux I__708 (
            .O(N__5145),
            .I(N__5133));
    LocalMux I__707 (
            .O(N__5142),
            .I(N__5130));
    Odrv4 I__706 (
            .O(N__5139),
            .I(\U712_CHIP_RAM.N_522 ));
    LocalMux I__705 (
            .O(N__5136),
            .I(\U712_CHIP_RAM.N_522 ));
    LocalMux I__704 (
            .O(N__5133),
            .I(\U712_CHIP_RAM.N_522 ));
    Odrv4 I__703 (
            .O(N__5130),
            .I(\U712_CHIP_RAM.N_522 ));
    CascadeMux I__702 (
            .O(N__5121),
            .I(\U712_CHIP_RAM.N_523_cascade_ ));
    InMux I__701 (
            .O(N__5118),
            .I(N__5115));
    LocalMux I__700 (
            .O(N__5115),
            .I(\U712_CHIP_RAM.BANK0_9 ));
    IoInMux I__699 (
            .O(N__5112),
            .I(N__5109));
    LocalMux I__698 (
            .O(N__5109),
            .I(N__5106));
    Span12Mux_s5_v I__697 (
            .O(N__5106),
            .I(N__5103));
    Span12Mux_v I__696 (
            .O(N__5103),
            .I(N__5099));
    InMux I__695 (
            .O(N__5102),
            .I(N__5096));
    Odrv12 I__694 (
            .O(N__5099),
            .I(BANK0_c));
    LocalMux I__693 (
            .O(N__5096),
            .I(BANK0_c));
    InMux I__692 (
            .O(N__5091),
            .I(N__5087));
    InMux I__691 (
            .O(N__5090),
            .I(N__5084));
    LocalMux I__690 (
            .O(N__5087),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__689 (
            .O(N__5084),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__688 (
            .O(N__5079),
            .I(N__5075));
    InMux I__687 (
            .O(N__5078),
            .I(N__5072));
    LocalMux I__686 (
            .O(N__5075),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__685 (
            .O(N__5072),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__684 (
            .O(N__5067),
            .I(N__5063));
    InMux I__683 (
            .O(N__5066),
            .I(N__5060));
    LocalMux I__682 (
            .O(N__5063),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__681 (
            .O(N__5060),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__680 (
            .O(N__5055),
            .I(\U712_CHIP_RAM.N_545_cascade_ ));
    InMux I__679 (
            .O(N__5052),
            .I(N__5046));
    CascadeMux I__678 (
            .O(N__5051),
            .I(N__5043));
    InMux I__677 (
            .O(N__5050),
            .I(N__5036));
    InMux I__676 (
            .O(N__5049),
            .I(N__5036));
    LocalMux I__675 (
            .O(N__5046),
            .I(N__5033));
    InMux I__674 (
            .O(N__5043),
            .I(N__5026));
    InMux I__673 (
            .O(N__5042),
            .I(N__5026));
    InMux I__672 (
            .O(N__5041),
            .I(N__5026));
    LocalMux I__671 (
            .O(N__5036),
            .I(\U712_CHIP_RAM.N_549 ));
    Odrv4 I__670 (
            .O(N__5033),
            .I(\U712_CHIP_RAM.N_549 ));
    LocalMux I__669 (
            .O(N__5026),
            .I(\U712_CHIP_RAM.N_549 ));
    InMux I__668 (
            .O(N__5019),
            .I(N__5010));
    InMux I__667 (
            .O(N__5018),
            .I(N__5010));
    InMux I__666 (
            .O(N__5017),
            .I(N__5010));
    LocalMux I__665 (
            .O(N__5010),
            .I(N__5006));
    InMux I__664 (
            .O(N__5009),
            .I(N__5002));
    Span4Mux_h I__663 (
            .O(N__5006),
            .I(N__4999));
    InMux I__662 (
            .O(N__5005),
            .I(N__4996));
    LocalMux I__661 (
            .O(N__5002),
            .I(\U712_CHIP_RAM.N_560 ));
    Odrv4 I__660 (
            .O(N__4999),
            .I(\U712_CHIP_RAM.N_560 ));
    LocalMux I__659 (
            .O(N__4996),
            .I(\U712_CHIP_RAM.N_560 ));
    CascadeMux I__658 (
            .O(N__4989),
            .I(N__4986));
    InMux I__657 (
            .O(N__4986),
            .I(N__4983));
    LocalMux I__656 (
            .O(N__4983),
            .I(\U712_CHIP_RAM.N_501 ));
    InMux I__655 (
            .O(N__4980),
            .I(N__4977));
    LocalMux I__654 (
            .O(N__4977),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1 ));
    InMux I__653 (
            .O(N__4974),
            .I(N__4968));
    InMux I__652 (
            .O(N__4973),
            .I(N__4968));
    LocalMux I__651 (
            .O(N__4968),
            .I(\U712_CHIP_RAM.N_515 ));
    InMux I__650 (
            .O(N__4965),
            .I(N__4962));
    LocalMux I__649 (
            .O(N__4962),
            .I(\U712_CHIP_RAM.N_516 ));
    CascadeMux I__648 (
            .O(N__4959),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ));
    InMux I__647 (
            .O(N__4956),
            .I(N__4952));
    InMux I__646 (
            .O(N__4955),
            .I(N__4949));
    LocalMux I__645 (
            .O(N__4952),
            .I(\U712_CHIP_RAM.N_519 ));
    LocalMux I__644 (
            .O(N__4949),
            .I(\U712_CHIP_RAM.N_519 ));
    InMux I__643 (
            .O(N__4944),
            .I(N__4941));
    LocalMux I__642 (
            .O(N__4941),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0 ));
    IoInMux I__641 (
            .O(N__4938),
            .I(N__4935));
    LocalMux I__640 (
            .O(N__4935),
            .I(N__4932));
    Span4Mux_s2_v I__639 (
            .O(N__4932),
            .I(N__4929));
    Sp12to4 I__638 (
            .O(N__4929),
            .I(N__4925));
    InMux I__637 (
            .O(N__4928),
            .I(N__4922));
    Span12Mux_h I__636 (
            .O(N__4925),
            .I(N__4919));
    LocalMux I__635 (
            .O(N__4922),
            .I(N__4916));
    Odrv12 I__634 (
            .O(N__4919),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__633 (
            .O(N__4916),
            .I(CONSTANT_ONE_NET));
    InMux I__632 (
            .O(N__4911),
            .I(N__4908));
    LocalMux I__631 (
            .O(N__4908),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_0 ));
    CascadeMux I__630 (
            .O(N__4905),
            .I(N__4899));
    InMux I__629 (
            .O(N__4904),
            .I(N__4890));
    InMux I__628 (
            .O(N__4903),
            .I(N__4890));
    InMux I__627 (
            .O(N__4902),
            .I(N__4887));
    InMux I__626 (
            .O(N__4899),
            .I(N__4884));
    InMux I__625 (
            .O(N__4898),
            .I(N__4875));
    InMux I__624 (
            .O(N__4897),
            .I(N__4875));
    InMux I__623 (
            .O(N__4896),
            .I(N__4875));
    InMux I__622 (
            .O(N__4895),
            .I(N__4875));
    LocalMux I__621 (
            .O(N__4890),
            .I(N__4872));
    LocalMux I__620 (
            .O(N__4887),
            .I(\U712_CHIP_RAM.N_78 ));
    LocalMux I__619 (
            .O(N__4884),
            .I(\U712_CHIP_RAM.N_78 ));
    LocalMux I__618 (
            .O(N__4875),
            .I(\U712_CHIP_RAM.N_78 ));
    Odrv4 I__617 (
            .O(N__4872),
            .I(\U712_CHIP_RAM.N_78 ));
    CEMux I__616 (
            .O(N__4863),
            .I(N__4858));
    CEMux I__615 (
            .O(N__4862),
            .I(N__4855));
    CEMux I__614 (
            .O(N__4861),
            .I(N__4852));
    LocalMux I__613 (
            .O(N__4858),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    LocalMux I__612 (
            .O(N__4855),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    LocalMux I__611 (
            .O(N__4852),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    CascadeMux I__610 (
            .O(N__4845),
            .I(\U712_CHIP_RAM.N_559_cascade_ ));
    InMux I__609 (
            .O(N__4842),
            .I(N__4836));
    InMux I__608 (
            .O(N__4841),
            .I(N__4836));
    LocalMux I__607 (
            .O(N__4836),
            .I(\U712_CHIP_RAM.N_665 ));
    CascadeMux I__606 (
            .O(N__4833),
            .I(\U712_CHIP_RAM.N_665_cascade_ ));
    InMux I__605 (
            .O(N__4830),
            .I(N__4827));
    LocalMux I__604 (
            .O(N__4827),
            .I(\U712_CHIP_RAM.N_471 ));
    CascadeMux I__603 (
            .O(N__4824),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ));
    InMux I__602 (
            .O(N__4821),
            .I(N__4817));
    InMux I__601 (
            .O(N__4820),
            .I(N__4814));
    LocalMux I__600 (
            .O(N__4817),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__599 (
            .O(N__4814),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__598 (
            .O(N__4809),
            .I(N__4805));
    InMux I__597 (
            .O(N__4808),
            .I(N__4802));
    LocalMux I__596 (
            .O(N__4805),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__595 (
            .O(N__4802),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__594 (
            .O(N__4797),
            .I(N__4793));
    InMux I__593 (
            .O(N__4796),
            .I(N__4790));
    LocalMux I__592 (
            .O(N__4793),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__591 (
            .O(N__4790),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__590 (
            .O(N__4785),
            .I(N__4782));
    LocalMux I__589 (
            .O(N__4782),
            .I(N__4779));
    Span12Mux_v I__588 (
            .O(N__4779),
            .I(N__4776));
    Span12Mux_h I__587 (
            .O(N__4776),
            .I(N__4773));
    Odrv12 I__586 (
            .O(N__4773),
            .I(A_c_14));
    InMux I__585 (
            .O(N__4770),
            .I(N__4767));
    LocalMux I__584 (
            .O(N__4767),
            .I(N__4764));
    Span4Mux_v I__583 (
            .O(N__4764),
            .I(N__4761));
    Sp12to4 I__582 (
            .O(N__4761),
            .I(N__4758));
    Span12Mux_h I__581 (
            .O(N__4758),
            .I(N__4755));
    Odrv12 I__580 (
            .O(N__4755),
            .I(A_c_7));
    InMux I__579 (
            .O(N__4752),
            .I(N__4748));
    InMux I__578 (
            .O(N__4751),
            .I(N__4745));
    LocalMux I__577 (
            .O(N__4748),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    LocalMux I__576 (
            .O(N__4745),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    InMux I__575 (
            .O(N__4740),
            .I(N__4736));
    InMux I__574 (
            .O(N__4739),
            .I(N__4733));
    LocalMux I__573 (
            .O(N__4736),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    LocalMux I__572 (
            .O(N__4733),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    CascadeMux I__571 (
            .O(N__4728),
            .I(N__4724));
    InMux I__570 (
            .O(N__4727),
            .I(N__4721));
    InMux I__569 (
            .O(N__4724),
            .I(N__4718));
    LocalMux I__568 (
            .O(N__4721),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__567 (
            .O(N__4718),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__566 (
            .O(N__4713),
            .I(N__4709));
    InMux I__565 (
            .O(N__4712),
            .I(N__4706));
    LocalMux I__564 (
            .O(N__4709),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    LocalMux I__563 (
            .O(N__4706),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__562 (
            .O(N__4701),
            .I(N__4698));
    LocalMux I__561 (
            .O(N__4698),
            .I(N__4695));
    Span4Mux_v I__560 (
            .O(N__4695),
            .I(N__4692));
    Sp12to4 I__559 (
            .O(N__4692),
            .I(N__4689));
    Span12Mux_h I__558 (
            .O(N__4689),
            .I(N__4686));
    Odrv12 I__557 (
            .O(N__4686),
            .I(A_c_8));
    InMux I__556 (
            .O(N__4683),
            .I(N__4680));
    LocalMux I__555 (
            .O(N__4680),
            .I(N__4677));
    Span4Mux_v I__554 (
            .O(N__4677),
            .I(N__4674));
    Sp12to4 I__553 (
            .O(N__4674),
            .I(N__4671));
    Span12Mux_h I__552 (
            .O(N__4671),
            .I(N__4668));
    Span12Mux_v I__551 (
            .O(N__4668),
            .I(N__4665));
    Odrv12 I__550 (
            .O(N__4665),
            .I(A_c_15));
    CascadeMux I__549 (
            .O(N__4662),
            .I(\U712_CHIP_RAM.N_669_cascade_ ));
    CascadeMux I__548 (
            .O(N__4659),
            .I(\U712_CHIP_RAM.N_520_cascade_ ));
    CascadeMux I__547 (
            .O(N__4656),
            .I(\U712_CYCLE_TERM.N_539_cascade_ ));
    InMux I__546 (
            .O(N__4653),
            .I(N__4647));
    InMux I__545 (
            .O(N__4652),
            .I(N__4644));
    InMux I__544 (
            .O(N__4651),
            .I(N__4639));
    InMux I__543 (
            .O(N__4650),
            .I(N__4639));
    LocalMux I__542 (
            .O(N__4647),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__541 (
            .O(N__4644),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__540 (
            .O(N__4639),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__539 (
            .O(N__4632),
            .I(N__4624));
    InMux I__538 (
            .O(N__4631),
            .I(N__4624));
    InMux I__537 (
            .O(N__4630),
            .I(N__4621));
    InMux I__536 (
            .O(N__4629),
            .I(N__4618));
    LocalMux I__535 (
            .O(N__4624),
            .I(CPU_TACKm));
    LocalMux I__534 (
            .O(N__4621),
            .I(CPU_TACKm));
    LocalMux I__533 (
            .O(N__4618),
            .I(CPU_TACKm));
    InMux I__532 (
            .O(N__4611),
            .I(N__4608));
    LocalMux I__531 (
            .O(N__4608),
            .I(N__4603));
    InMux I__530 (
            .O(N__4607),
            .I(N__4600));
    InMux I__529 (
            .O(N__4606),
            .I(N__4597));
    Span4Mux_h I__528 (
            .O(N__4603),
            .I(N__4594));
    LocalMux I__527 (
            .O(N__4600),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    LocalMux I__526 (
            .O(N__4597),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    Odrv4 I__525 (
            .O(N__4594),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    InMux I__524 (
            .O(N__4587),
            .I(N__4584));
    LocalMux I__523 (
            .O(N__4584),
            .I(N__4581));
    Span4Mux_v I__522 (
            .O(N__4581),
            .I(N__4578));
    Span4Mux_v I__521 (
            .O(N__4578),
            .I(N__4575));
    Span4Mux_h I__520 (
            .O(N__4575),
            .I(N__4572));
    Sp12to4 I__519 (
            .O(N__4572),
            .I(N__4569));
    Odrv12 I__518 (
            .O(N__4569),
            .I(A_c_6));
    InMux I__517 (
            .O(N__4566),
            .I(N__4563));
    LocalMux I__516 (
            .O(N__4563),
            .I(N__4560));
    Span4Mux_v I__515 (
            .O(N__4560),
            .I(N__4557));
    Sp12to4 I__514 (
            .O(N__4557),
            .I(N__4554));
    Span12Mux_h I__513 (
            .O(N__4554),
            .I(N__4551));
    Odrv12 I__512 (
            .O(N__4551),
            .I(A_c_13));
    InMux I__511 (
            .O(N__4548),
            .I(N__4545));
    LocalMux I__510 (
            .O(N__4545),
            .I(N__4542));
    Span12Mux_v I__509 (
            .O(N__4542),
            .I(N__4539));
    Span12Mux_h I__508 (
            .O(N__4539),
            .I(N__4536));
    Odrv12 I__507 (
            .O(N__4536),
            .I(A_c_18));
    InMux I__506 (
            .O(N__4533),
            .I(N__4530));
    LocalMux I__505 (
            .O(N__4530),
            .I(N__4527));
    Span12Mux_v I__504 (
            .O(N__4527),
            .I(N__4524));
    Span12Mux_h I__503 (
            .O(N__4524),
            .I(N__4521));
    Odrv12 I__502 (
            .O(N__4521),
            .I(A_c_16));
    CascadeMux I__501 (
            .O(N__4518),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_ ));
    InMux I__500 (
            .O(N__4515),
            .I(N__4512));
    LocalMux I__499 (
            .O(N__4512),
            .I(N__4509));
    Span4Mux_h I__498 (
            .O(N__4509),
            .I(N__4506));
    Sp12to4 I__497 (
            .O(N__4506),
            .I(N__4503));
    Span12Mux_v I__496 (
            .O(N__4503),
            .I(N__4500));
    Odrv12 I__495 (
            .O(N__4500),
            .I(A_c_5));
    InMux I__494 (
            .O(N__4497),
            .I(N__4494));
    LocalMux I__493 (
            .O(N__4494),
            .I(N__4491));
    Span12Mux_v I__492 (
            .O(N__4491),
            .I(N__4488));
    Span12Mux_h I__491 (
            .O(N__4488),
            .I(N__4485));
    Odrv12 I__490 (
            .O(N__4485),
            .I(A_c_12));
    InMux I__489 (
            .O(N__4482),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    CascadeMux I__488 (
            .O(N__4479),
            .I(\U712_CHIP_RAM.N_666_cascade_ ));
    CascadeMux I__487 (
            .O(N__4476),
            .I(\U712_CHIP_RAM.N_393_cascade_ ));
    CascadeMux I__486 (
            .O(N__4473),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_ ));
    CEMux I__485 (
            .O(N__4470),
            .I(N__4467));
    LocalMux I__484 (
            .O(N__4467),
            .I(N__4464));
    Span4Mux_h I__483 (
            .O(N__4464),
            .I(N__4461));
    Span4Mux_h I__482 (
            .O(N__4461),
            .I(N__4458));
    Odrv4 I__481 (
            .O(N__4458),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0 ));
    InMux I__480 (
            .O(N__4455),
            .I(N__4452));
    LocalMux I__479 (
            .O(N__4452),
            .I(N__4449));
    Odrv4 I__478 (
            .O(N__4449),
            .I(\U712_CHIP_RAM.CLK_EN_6_0 ));
    CascadeMux I__477 (
            .O(N__4446),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_0_cascade_ ));
    IoInMux I__476 (
            .O(N__4443),
            .I(N__4440));
    LocalMux I__475 (
            .O(N__4440),
            .I(N__4437));
    IoSpan4Mux I__474 (
            .O(N__4437),
            .I(N__4434));
    IoSpan4Mux I__473 (
            .O(N__4434),
            .I(N__4431));
    Sp12to4 I__472 (
            .O(N__4431),
            .I(N__4428));
    Span12Mux_s7_h I__471 (
            .O(N__4428),
            .I(N__4425));
    Span12Mux_h I__470 (
            .O(N__4425),
            .I(N__4421));
    InMux I__469 (
            .O(N__4424),
            .I(N__4418));
    Odrv12 I__468 (
            .O(N__4421),
            .I(CLK_EN_c));
    LocalMux I__467 (
            .O(N__4418),
            .I(CLK_EN_c));
    InMux I__466 (
            .O(N__4413),
            .I(N__4410));
    LocalMux I__465 (
            .O(N__4410),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0 ));
    InMux I__464 (
            .O(N__4407),
            .I(N__4404));
    LocalMux I__463 (
            .O(N__4404),
            .I(\U712_CHIP_RAM.N_504 ));
    CascadeMux I__462 (
            .O(N__4401),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_a2_0_cascade_ ));
    InMux I__461 (
            .O(N__4398),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__460 (
            .O(N__4395),
            .I(N__4392));
    LocalMux I__459 (
            .O(N__4392),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__458 (
            .O(N__4389),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__457 (
            .O(N__4386),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__456 (
            .O(N__4383),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__455 (
            .O(N__4380),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__454 (
            .O(N__4377),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    CascadeMux I__453 (
            .O(N__4374),
            .I(\U712_CHIP_RAM.N_375_cascade_ ));
    CascadeMux I__452 (
            .O(N__4371),
            .I(N__4367));
    InMux I__451 (
            .O(N__4370),
            .I(N__4364));
    InMux I__450 (
            .O(N__4367),
            .I(N__4361));
    LocalMux I__449 (
            .O(N__4364),
            .I(N__4358));
    LocalMux I__448 (
            .O(N__4361),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    Odrv4 I__447 (
            .O(N__4358),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    CascadeMux I__446 (
            .O(N__4353),
            .I(N__4350));
    InMux I__445 (
            .O(N__4350),
            .I(N__4347));
    LocalMux I__444 (
            .O(N__4347),
            .I(\U712_CHIP_RAM.N_498 ));
    CascadeMux I__443 (
            .O(N__4344),
            .I(\U712_CHIP_RAM.N_547_cascade_ ));
    CascadeMux I__442 (
            .O(N__4341),
            .I(\U712_CHIP_RAM.N_501_cascade_ ));
    InMux I__441 (
            .O(N__4338),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__440 (
            .O(N__4335),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__439 (
            .O(N__4332),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__438 (
            .O(N__4329),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__437 (
            .O(N__4326),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__436 (
            .O(N__4323),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__435 (
            .O(N__4320),
            .I(N__4296));
    ClkMux I__434 (
            .O(N__4319),
            .I(N__4296));
    ClkMux I__433 (
            .O(N__4318),
            .I(N__4296));
    ClkMux I__432 (
            .O(N__4317),
            .I(N__4296));
    ClkMux I__431 (
            .O(N__4316),
            .I(N__4296));
    ClkMux I__430 (
            .O(N__4315),
            .I(N__4296));
    ClkMux I__429 (
            .O(N__4314),
            .I(N__4296));
    ClkMux I__428 (
            .O(N__4313),
            .I(N__4296));
    GlobalMux I__427 (
            .O(N__4296),
            .I(N__4293));
    gio2CtrlBuf I__426 (
            .O(N__4293),
            .I(C1_c_g));
    CascadeMux I__425 (
            .O(N__4290),
            .I(\U712_CHIP_RAM.N_371_cascade_ ));
    CascadeMux I__424 (
            .O(N__4287),
            .I(\U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_2_cascade_ ));
    InMux I__423 (
            .O(N__4284),
            .I(N__4281));
    LocalMux I__422 (
            .O(N__4281),
            .I(\U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1 ));
    InMux I__421 (
            .O(N__4278),
            .I(N__4274));
    InMux I__420 (
            .O(N__4277),
            .I(N__4271));
    LocalMux I__419 (
            .O(N__4274),
            .I(N__4268));
    LocalMux I__418 (
            .O(N__4271),
            .I(\U712_CYCLE_TERM.N_565 ));
    Odrv4 I__417 (
            .O(N__4268),
            .I(\U712_CYCLE_TERM.N_565 ));
    InMux I__416 (
            .O(N__4263),
            .I(N__4259));
    InMux I__415 (
            .O(N__4262),
            .I(N__4256));
    LocalMux I__414 (
            .O(N__4259),
            .I(N__4253));
    LocalMux I__413 (
            .O(N__4256),
            .I(\U712_CYCLE_TERM.N_407 ));
    Odrv4 I__412 (
            .O(N__4253),
            .I(\U712_CYCLE_TERM.N_407 ));
    InMux I__411 (
            .O(N__4248),
            .I(N__4245));
    LocalMux I__410 (
            .O(N__4245),
            .I(N__4242));
    Odrv4 I__409 (
            .O(N__4242),
            .I(\U712_CYCLE_TERM.N_534 ));
    InMux I__408 (
            .O(N__4239),
            .I(bfn_9_9_0_));
    InMux I__407 (
            .O(N__4236),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__406 (
            .O(N__4233),
            .I(N__4227));
    InMux I__405 (
            .O(N__4232),
            .I(N__4227));
    LocalMux I__404 (
            .O(N__4227),
            .I(\U712_CHIP_RAM.N_373 ));
    InMux I__403 (
            .O(N__4224),
            .I(N__4221));
    LocalMux I__402 (
            .O(N__4221),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0 ));
    InMux I__401 (
            .O(N__4218),
            .I(N__4215));
    LocalMux I__400 (
            .O(N__4215),
            .I(N__4212));
    Odrv4 I__399 (
            .O(N__4212),
            .I(\U712_CHIP_RAM.N_409 ));
    CascadeMux I__398 (
            .O(N__4209),
            .I(\U712_REG_SM.N_486_cascade_ ));
    InMux I__397 (
            .O(N__4206),
            .I(N__4203));
    LocalMux I__396 (
            .O(N__4203),
            .I(\U712_CHIP_RAM.CLK_EN_6_0_a3_0_a2_1 ));
    IoInMux I__395 (
            .O(N__4200),
            .I(N__4197));
    LocalMux I__394 (
            .O(N__4197),
            .I(N__4194));
    Span12Mux_s9_v I__393 (
            .O(N__4194),
            .I(N__4191));
    Odrv12 I__392 (
            .O(N__4191),
            .I(N_490));
    CEMux I__391 (
            .O(N__4188),
            .I(N__4185));
    LocalMux I__390 (
            .O(N__4185),
            .I(N__4182));
    Span4Mux_v I__389 (
            .O(N__4182),
            .I(N__4179));
    Odrv4 I__388 (
            .O(N__4179),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0 ));
    CascadeMux I__387 (
            .O(N__4176),
            .I(\U712_CHIP_RAM.N_554_cascade_ ));
    CascadeMux I__386 (
            .O(N__4173),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_a2_0_cascade_ ));
    IoInMux I__385 (
            .O(N__4170),
            .I(N__4167));
    LocalMux I__384 (
            .O(N__4167),
            .I(N__4164));
    IoSpan4Mux I__383 (
            .O(N__4164),
            .I(N__4161));
    Span4Mux_s3_v I__382 (
            .O(N__4161),
            .I(N__4158));
    Odrv4 I__381 (
            .O(N__4158),
            .I(CLK80_PLL_i_i));
    CascadeMux I__380 (
            .O(N__4155),
            .I(DBRn_c_i_cascade_));
    IoInMux I__379 (
            .O(N__4152),
            .I(N__4149));
    LocalMux I__378 (
            .O(N__4149),
            .I(N__4146));
    IoSpan4Mux I__377 (
            .O(N__4146),
            .I(N__4143));
    Sp12to4 I__376 (
            .O(N__4143),
            .I(N__4140));
    Odrv12 I__375 (
            .O(N__4140),
            .I(DBRn_c_i_0));
    CascadeMux I__374 (
            .O(N__4137),
            .I(N__4134));
    InMux I__373 (
            .O(N__4134),
            .I(N__4131));
    LocalMux I__372 (
            .O(N__4131),
            .I(DBRn_c_i));
    IoInMux I__371 (
            .O(N__4128),
            .I(N__4125));
    LocalMux I__370 (
            .O(N__4125),
            .I(N__4122));
    IoSpan4Mux I__369 (
            .O(N__4122),
            .I(N__4119));
    Span4Mux_s2_v I__368 (
            .O(N__4119),
            .I(N__4116));
    Sp12to4 I__367 (
            .O(N__4116),
            .I(N__4113));
    Span12Mux_v I__366 (
            .O(N__4113),
            .I(N__4110));
    Span12Mux_h I__365 (
            .O(N__4110),
            .I(N__4107));
    Odrv12 I__364 (
            .O(N__4107),
            .I(U712_CYCLE_TERM_TCIn_0_i));
    CascadeMux I__363 (
            .O(N__4104),
            .I(N__4100));
    InMux I__362 (
            .O(N__4103),
            .I(N__4097));
    InMux I__361 (
            .O(N__4100),
            .I(N__4094));
    LocalMux I__360 (
            .O(N__4097),
            .I(\U712_CYCLE_TERM.RAM_CYCLEZ0 ));
    LocalMux I__359 (
            .O(N__4094),
            .I(\U712_CYCLE_TERM.RAM_CYCLEZ0 ));
    IoInMux I__358 (
            .O(N__4089),
            .I(N__4086));
    LocalMux I__357 (
            .O(N__4086),
            .I(N__4083));
    IoSpan4Mux I__356 (
            .O(N__4083),
            .I(N__4080));
    Span4Mux_s2_v I__355 (
            .O(N__4080),
            .I(N__4077));
    Sp12to4 I__354 (
            .O(N__4077),
            .I(N__4074));
    Span12Mux_v I__353 (
            .O(N__4074),
            .I(N__4071));
    Odrv12 I__352 (
            .O(N__4071),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__4314));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__4317));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .I(N__4318));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__4313));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .I(N__4315));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .I(N__4316));
    INV \INVU712_CHIP_RAM.DMA_A20C  (
            .O(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .I(N__4319));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__6962),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7959),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4152),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__7011),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_2_1_3.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_2_1_3.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_2_1_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_2_1_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9042),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_5_12_3.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_5_12_3.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_5_12_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_5_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7499),
            .lcout(DBRn_c_i),
            .ltout(DBRn_c_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_12_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4155),
            .in3(N__10293),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_A20_LC_6_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A20_LC_6_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A20_LC_6_12_0 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A20_LC_6_12_0  (
            .in0(N__10416),
            .in1(N__10629),
            .in2(N__4137),
            .in3(N__5210),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .ce(),
            .sr(N__10254));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_7_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_7_10_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_7_10_6  (
            .in0(N__10292),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4224),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.RAM_CYCLE_RNILITE_LC_7_11_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.RAM_CYCLE_RNILITE_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.RAM_CYCLE_RNILITE_LC_7_11_4 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U712_CYCLE_TERM.RAM_CYCLE_RNILITE_LC_7_11_4  (
            .in0(N__5272),
            .in1(N__4103),
            .in2(_gnd_net_),
            .in3(N__7396),
            .lcout(U712_CYCLE_TERM_TCIn_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.RAM_CYCLE_LC_7_12_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.RAM_CYCLE_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.RAM_CYCLE_LC_7_12_0 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \U712_CYCLE_TERM.RAM_CYCLE_LC_7_12_0  (
            .in0(N__8516),
            .in1(N__4248),
            .in2(N__4104),
            .in3(N__7442),
            .lcout(\U712_CYCLE_TERM.RAM_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9031),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_7_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_7_12_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_2_LC_7_12_1  (
            .in0(N__9932),
            .in1(N__11216),
            .in2(_gnd_net_),
            .in3(N__6774),
            .lcout(\U712_CHIP_RAM.CLK_EN_6_0_a3_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__8097),
            .in2(_gnd_net_),
            .in3(N__7898),
            .lcout(),
            .ltout(\U712_REG_SM.N_486_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_7_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_7_13_1 .LUT_INIT=16'b1110110011100100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_7_13_1  (
            .in0(N__8518),
            .in1(N__10117),
            .in2(N__4209),
            .in3(N__5673),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9035),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_13_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_13_4  (
            .in0(N__4206),
            .in1(N__5334),
            .in2(N__6186),
            .in3(N__6101),
            .lcout(\U712_CHIP_RAM.CLK_EN_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_i_i_a2_LC_8_6_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_i_i_a2_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_i_i_a2_LC_8_6_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_i_i_a2_LC_8_6_2  (
            .in0(N__10130),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9946),
            .lcout(N_490),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_8_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_8_10_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_8_10_0  (
            .in0(N__6903),
            .in1(N__6294),
            .in2(_gnd_net_),
            .in3(N__6003),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9019),
            .ce(N__4188),
            .sr(N__10255));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_8_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_8_11_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_8_11_0  (
            .in0(N__6766),
            .in1(N__6579),
            .in2(_gnd_net_),
            .in3(N__8628),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_554_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOJRU2_1_LC_8_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOJRU2_1_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOJRU2_1_LC_8_11_1 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOJRU2_1_LC_8_11_1  (
            .in0(N__4232),
            .in1(N__6657),
            .in2(N__4176),
            .in3(N__5380),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_1_LC_8_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_1_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_1_LC_8_11_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_1_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4173),
            .in3(N__5180),
            .lcout(\U712_CHIP_RAM.N_522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_8_11_3 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_8_11_3  (
            .in0(N__11213),
            .in1(N__6765),
            .in2(_gnd_net_),
            .in3(N__6578),
            .lcout(\U712_CHIP_RAM.N_373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_8_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_8_11_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_8_11_4  (
            .in0(N__6767),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8431),
            .lcout(\U712_CHIP_RAM.N_560 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_8_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_8_11_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_8_11_5  (
            .in0(N__8430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5557),
            .lcout(\U712_CHIP_RAM.N_572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_8_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_8_11_6 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_8_11_6  (
            .in0(N__4218),
            .in1(N__11214),
            .in2(N__4371),
            .in3(N__8432),
            .lcout(WRITE_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9023),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_11_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_11_7  (
            .in0(N__4233),
            .in1(N__5522),
            .in2(N__4353),
            .in3(N__6658),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_12_0 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_12_0  (
            .in0(N__4395),
            .in1(N__8482),
            .in2(N__4905),
            .in3(N__4370),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9027),
            .ce(N__4863),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_0_LC_8_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_0_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_0_LC_8_12_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_0_LC_8_12_1  (
            .in0(N__11215),
            .in1(N__6768),
            .in2(_gnd_net_),
            .in3(N__6594),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNIDG0M2_4_LC_8_12_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNIDG0M2_4_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNIDG0M2_4_LC_8_12_3 .LUT_INIT=16'b1010111110101110;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNIDG0M2_4_LC_8_12_3  (
            .in0(N__4611),
            .in1(N__4278),
            .in2(N__6323),
            .in3(N__4263),
            .lcout(\U712_CYCLE_TERM.un13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_13_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__6901),
            .in2(_gnd_net_),
            .in3(N__6243),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9032),
            .ce(N__4470),
            .sr(N__10243));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_13_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__8620),
            .in2(_gnd_net_),
            .in3(N__5393),
            .lcout(\U712_CHIP_RAM.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_13_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_13_6  (
            .in0(N__10068),
            .in1(N__5747),
            .in2(_gnd_net_),
            .in3(N__6900),
            .lcout(\U712_CHIP_RAM.N_409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_8_14_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_8_14_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_8_14_0  (
            .in0(N__4284),
            .in1(N__11231),
            .in2(_gnd_net_),
            .in3(N__6807),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_8_14_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_8_14_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_8_14_1  (
            .in0(N__6177),
            .in1(N__6102),
            .in2(N__4287),
            .in3(N__5396),
            .lcout(\U712_CHIP_RAM.N_504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_0_a2_1_0_LC_8_14_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_0_a2_1_0_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_0_a2_1_0_LC_8_14_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_0_a2_1_0_LC_8_14_2  (
            .in0(N__4629),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5777),
            .lcout(\U712_CYCLE_TERM.N_565 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_5_LC_8_14_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_5_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_5_LC_8_14_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_5_LC_8_14_3  (
            .in0(N__9895),
            .in1(N__6690),
            .in2(_gnd_net_),
            .in3(N__6595),
            .lcout(\U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNI05SV_3_LC_8_14_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNI05SV_3_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNI05SV_3_LC_8_14_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNI05SV_3_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__6340),
            .in2(_gnd_net_),
            .in3(N__5310),
            .lcout(\U712_CYCLE_TERM.N_407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_14_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_14_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_8_14_7  (
            .in0(N__4606),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8517),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9036),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_15_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_15_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_15_0 .LUT_INIT=16'b0101000001010100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_8_15_0  (
            .in0(N__4607),
            .in1(N__4277),
            .in2(N__6324),
            .in3(N__4262),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9038),
            .ce(),
            .sr(N__10231));
    defparam \U712_CYCLE_TERM.RAM_CYCLE_RNO_0_LC_8_15_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.RAM_CYCLE_RNO_0_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.RAM_CYCLE_RNO_0_LC_8_15_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CYCLE_TERM.RAM_CYCLE_RNO_0_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__4652),
            .in2(_gnd_net_),
            .in3(N__4630),
            .lcout(\U712_CYCLE_TERM.N_534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_9_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_9_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__4713),
            .in2(_gnd_net_),
            .in3(N__4239),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__4320),
            .ce(),
            .sr(N__5922));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_9_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_9_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__4740),
            .in2(_gnd_net_),
            .in3(N__4236),
            .lcout(\U712_CHIP_RAM.REFRESH5lto1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__4320),
            .ce(),
            .sr(N__5922));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_9_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__4752),
            .in2(_gnd_net_),
            .in3(N__4338),
            .lcout(\U712_CHIP_RAM.REFRESH5lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__4320),
            .ce(),
            .sr(N__5922));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_9_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_9_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__6377),
            .in2(_gnd_net_),
            .in3(N__4335),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__4320),
            .ce(),
            .sr(N__5922));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_9_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__4727),
            .in2(_gnd_net_),
            .in3(N__4332),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__4320),
            .ce(),
            .sr(N__5922));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_9_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_9_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__4797),
            .in2(_gnd_net_),
            .in3(N__4329),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__4320),
            .ce(),
            .sr(N__5922));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_9_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_9_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__4809),
            .in2(_gnd_net_),
            .in3(N__4326),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__4320),
            .ce(),
            .sr(N__5922));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_9_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__4821),
            .in2(_gnd_net_),
            .in3(N__4323),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4320),
            .ce(),
            .sr(N__5922));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_10_0 .LUT_INIT=16'b0000001001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_10_0  (
            .in0(N__6806),
            .in1(N__5394),
            .in2(N__6692),
            .in3(N__6566),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_371_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_4_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_4_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_4_LC_9_10_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_4_LC_9_10_1  (
            .in0(N__6164),
            .in1(N__6022),
            .in2(N__4290),
            .in3(N__6094),
            .lcout(\U712_CHIP_RAM.N_519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_10_2 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_10_2  (
            .in0(N__8520),
            .in1(_gnd_net_),
            .in2(N__5153),
            .in3(N__4830),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_10_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_10_3  (
            .in0(N__5009),
            .in1(N__5517),
            .in2(N__6587),
            .in3(N__6687),
            .lcout(\U712_CHIP_RAM.N_516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_1_LC_9_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_1_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_1_LC_9_10_4 .LUT_INIT=16'b0010000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_1_LC_9_10_4  (
            .in0(N__8519),
            .in1(N__5395),
            .in2(N__6693),
            .in3(N__6567),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIR9VE1_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIR9VE1_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIR9VE1_LC_9_10_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIR9VE1_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__6897),
            .in2(_gnd_net_),
            .in3(N__6293),
            .lcout(\U712_CHIP_RAM.N_375 ),
            .ltout(\U712_CHIP_RAM.N_375_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIPCS25_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIPCS25_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIPCS25_LC_9_10_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIPCS25_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4374),
            .in3(N__6238),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_11_0 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_11_0  (
            .in0(N__5556),
            .in1(N__8427),
            .in2(N__6808),
            .in3(N__4842),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9020),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_9_11_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_9_11_1  (
            .in0(N__6896),
            .in1(N__6286),
            .in2(_gnd_net_),
            .in3(N__6227),
            .lcout(\U712_CHIP_RAM.N_498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_9_11_2 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_9_11_2  (
            .in0(N__5990),
            .in1(N__6028),
            .in2(N__6178),
            .in3(N__6201),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_9_11_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_9_11_3  (
            .in0(N__6144),
            .in1(N__5555),
            .in2(_gnd_net_),
            .in3(N__6075),
            .lcout(\U712_CHIP_RAM.N_547 ),
            .ltout(\U712_CHIP_RAM.N_547_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_4_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_4_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_4_LC_9_11_4 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_4_LC_9_11_4  (
            .in0(N__5005),
            .in1(N__4841),
            .in2(N__4344),
            .in3(N__5049),
            .lcout(\U712_CHIP_RAM.N_501 ),
            .ltout(\U712_CHIP_RAM.N_501_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG9KPG_2_LC_9_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG9KPG_2_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG9KPG_2_LC_9_11_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIG9KPG_2_LC_9_11_5  (
            .in0(N__8428),
            .in1(N__5145),
            .in2(N__4341),
            .in3(N__5991),
            .lcout(\U712_CHIP_RAM.N_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVTLS1_7_LC_9_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVTLS1_7_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVTLS1_7_LC_9_11_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVTLS1_7_LC_9_11_6  (
            .in0(N__6076),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8429),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE24B8_2_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE24B8_2_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE24B8_2_LC_9_11_7 .LUT_INIT=16'b1100000011100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIE24B8_2_LC_9_11_7  (
            .in0(N__5050),
            .in1(N__4955),
            .in2(N__4401),
            .in3(N__6785),
            .lcout(\U712_CHIP_RAM.N_515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_9_12_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_9_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__6571),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_12_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_12_1  (
            .in0(N__4895),
            .in1(N__5386),
            .in2(_gnd_net_),
            .in3(N__4398),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__9024),
            .ce(N__4861),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_12_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__6784),
            .in2(_gnd_net_),
            .in3(N__4389),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_12_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_12_3  (
            .in0(N__4896),
            .in1(N__6678),
            .in2(_gnd_net_),
            .in3(N__4386),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__9024),
            .ce(N__4861),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_12_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_12_4  (
            .in0(N__4903),
            .in1(N__6163),
            .in2(_gnd_net_),
            .in3(N__4383),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__9024),
            .ce(N__4861),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_12_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_12_5  (
            .in0(N__4897),
            .in1(N__5067),
            .in2(_gnd_net_),
            .in3(N__4380),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__9024),
            .ce(N__4861),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_12_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_12_6  (
            .in0(N__4904),
            .in1(N__5079),
            .in2(_gnd_net_),
            .in3(N__4377),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__9024),
            .ce(N__4861),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_12_7  (
            .in0(N__4898),
            .in1(N__5091),
            .in2(_gnd_net_),
            .in3(N__4482),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9024),
            .ce(N__4861),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_9_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_9_13_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_9_13_1  (
            .in0(N__6146),
            .in1(N__5330),
            .in2(N__5562),
            .in3(N__6080),
            .lcout(\U712_CHIP_RAM.N_666 ),
            .ltout(\U712_CHIP_RAM.N_666_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIJH788_LC_9_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIJH788_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIJH788_LC_9_13_2 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNIJH788_LC_9_13_2  (
            .in0(N__6810),
            .in1(N__8618),
            .in2(N__4479),
            .in3(N__5714),
            .lcout(\U712_CHIP_RAM.N_393 ),
            .ltout(\U712_CHIP_RAM.N_393_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFS4TD_2_LC_9_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFS4TD_2_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFS4TD_2_LC_9_13_3 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIFS4TD_2_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__6811),
            .in2(N__4476),
            .in3(N__5152),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_13_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4473),
            .in3(N__10290),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_13_5 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_13_5  (
            .in0(N__8619),
            .in1(N__6812),
            .in2(_gnd_net_),
            .in3(N__5580),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_13_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_13_6 .LUT_INIT=16'b0101111101010000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_9_13_6  (
            .in0(N__4455),
            .in1(_gnd_net_),
            .in2(N__4446),
            .in3(N__4424),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9028),
            .ce(),
            .sr(N__10236));
    defparam \U712_CHIP_RAM.DBENn_LC_9_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_9_13_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_9_13_7 .LUT_INIT=16'b0010111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_9_13_7  (
            .in0(N__8679),
            .in1(N__4413),
            .in2(N__6002),
            .in3(N__9516),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9028),
            .ce(),
            .sr(N__10236));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_9_14_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_9_14_1 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_LC_9_14_1  (
            .in0(N__4407),
            .in1(N__11235),
            .in2(N__5400),
            .in3(N__9964),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9033),
            .ce(N__5592),
            .sr(N__10232));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_15_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_15_0 .LUT_INIT=16'b0000000100001111;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_15_0  (
            .in0(N__4632),
            .in1(N__5773),
            .in2(N__5318),
            .in3(N__4651),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_539_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_15_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_15_1 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_9_15_1  (
            .in0(N__8047),
            .in1(N__4653),
            .in2(N__4656),
            .in3(N__8521),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9037),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_15_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_15_3 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_15_3  (
            .in0(N__4650),
            .in1(N__5772),
            .in2(_gnd_net_),
            .in3(N__4631),
            .lcout(\U712_CYCLE_TERM.TACK_EN_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_15_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_15_6 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_9_15_6  (
            .in0(N__8522),
            .in1(_gnd_net_),
            .in2(N__5319),
            .in3(N__8048),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9037),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_0  (
            .in0(N__4587),
            .in1(N__4566),
            .in2(_gnd_net_),
            .in3(N__9739),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_7_2  (
            .in0(N__4548),
            .in1(N__4533),
            .in2(_gnd_net_),
            .in3(N__9740),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_7_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_7_3  (
            .in0(N__9741),
            .in1(N__9965),
            .in2(N__4518),
            .in3(N__7920),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_10_8_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_8_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_8_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_8_3  (
            .in0(N__4515),
            .in1(N__4497),
            .in2(_gnd_net_),
            .in3(N__9742),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_8_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_8_4  (
            .in0(N__9743),
            .in1(N__9950),
            .in2(N__4824),
            .in3(N__7935),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_9_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_9_1  (
            .in0(N__4820),
            .in1(N__4808),
            .in2(_gnd_net_),
            .in3(N__4796),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_9_3  (
            .in0(N__4785),
            .in1(N__4770),
            .in2(_gnd_net_),
            .in3(N__9698),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_9_4 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_9_4  (
            .in0(N__4751),
            .in1(N__4739),
            .in2(N__4728),
            .in3(N__4712),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_9_5  (
            .in0(N__4701),
            .in1(N__4683),
            .in2(_gnd_net_),
            .in3(N__9697),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_10_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_10_0  (
            .in0(N__5523),
            .in1(N__6688),
            .in2(_gnd_net_),
            .in3(N__5019),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_669_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_10_1 .LUT_INIT=16'b1000100010001011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_10_1  (
            .in0(N__7216),
            .in1(N__5834),
            .in2(N__4662),
            .in3(N__4974),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9012),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_2  (
            .in0(N__5183),
            .in1(N__6689),
            .in2(N__6597),
            .in3(N__5018),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_520_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_3 .LUT_INIT=16'b1100110100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_3  (
            .in0(N__4944),
            .in1(N__5833),
            .in2(N__4659),
            .in3(N__9738),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9012),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_10_4 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_10_4  (
            .in0(N__11242),
            .in1(N__5017),
            .in2(N__6596),
            .in3(N__5518),
            .lcout(\U712_CHIP_RAM.N_517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_10_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_10_10_5 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_10_10_5  (
            .in0(N__6200),
            .in1(N__5182),
            .in2(N__4989),
            .in3(N__4980),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_10_6 .LUT_INIT=16'b1111000100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_10_6  (
            .in0(N__4973),
            .in1(N__4965),
            .in2(N__4959),
            .in3(N__7120),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9012),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_10_7 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_10_7  (
            .in0(N__6435),
            .in1(N__4956),
            .in2(N__6902),
            .in3(N__6239),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_11_1 .LUT_INIT=16'b0011001101011010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_11_1  (
            .in0(N__4928),
            .in1(N__4911),
            .in2(N__6577),
            .in3(N__4902),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9015),
            .ce(N__4862),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_1_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_1_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_1_LC_10_11_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_1_LC_10_11_2  (
            .in0(N__5376),
            .in1(N__6651),
            .in2(_gnd_net_),
            .in3(N__6546),
            .lcout(\U712_CHIP_RAM.N_549 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_0_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_0_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_0_LC_10_11_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_0_LC_10_11_3  (
            .in0(N__6547),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6659),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_559_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_4_LC_10_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_4_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_4_LC_10_11_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_4_LC_10_11_4  (
            .in0(N__5377),
            .in1(N__6147),
            .in2(N__4845),
            .in3(N__6081),
            .lcout(\U712_CHIP_RAM.N_665 ),
            .ltout(\U712_CHIP_RAM.N_665_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_11_5 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_11_5  (
            .in0(N__6813),
            .in1(N__5181),
            .in2(N__4833),
            .in3(N__5052),
            .lcout(\U712_CHIP_RAM.N_471 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_10_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_10_12_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_10_12_0  (
            .in0(N__6277),
            .in1(N__6898),
            .in2(_gnd_net_),
            .in3(N__5988),
            .lcout(),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_10_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_10_12_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_2_LC_10_12_1  (
            .in0(N__10624),
            .in1(_gnd_net_),
            .in2(N__5232),
            .in3(N__5229),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_506_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_10_12_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_1_LC_10_12_2  (
            .in0(N__6881),
            .in1(N__5989),
            .in2(N__5214),
            .in3(N__5211),
            .lcout(\U712_CHIP_RAM.BANK0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_2_LC_10_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_2_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_2_LC_10_12_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_2_LC_10_12_3  (
            .in0(N__6790),
            .in1(N__6082),
            .in2(_gnd_net_),
            .in3(N__5042),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_10_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_10_12_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_0_LC_10_12_4  (
            .in0(N__5196),
            .in1(N__6791),
            .in2(N__5051),
            .in3(N__5184),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_523_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.BANK0_LC_10_12_5 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \U712_CHIP_RAM.BANK0_LC_10_12_5  (
            .in0(N__5102),
            .in1(N__5157),
            .in2(N__5121),
            .in3(N__5118),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9021),
            .ce(),
            .sr(N__10237));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_10_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_10_12_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_10_12_6  (
            .in0(N__5090),
            .in1(N__5078),
            .in2(_gnd_net_),
            .in3(N__5066),
            .lcout(\U712_CHIP_RAM.N_545 ),
            .ltout(\U712_CHIP_RAM.N_545_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_10_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_10_12_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_10_12_7  (
            .in0(N__5548),
            .in1(N__6789),
            .in2(N__5055),
            .in3(N__5041),
            .lcout(\U712_CHIP_RAM.N_562 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_10_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_10_13_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_10_13_0  (
            .in0(N__5462),
            .in1(N__5503),
            .in2(N__6680),
            .in3(N__5568),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_10_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_10_13_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_10_13_1  (
            .in0(N__10289),
            .in1(_gnd_net_),
            .in2(N__5595),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_10_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_10_13_2 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_10_13_2  (
            .in0(N__6653),
            .in1(N__5579),
            .in2(N__5516),
            .in3(N__6809),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_13_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_13_3  (
            .in0(N__5379),
            .in1(N__6145),
            .in2(N__6093),
            .in3(N__5558),
            .lcout(\U712_CHIP_RAM.N_557 ),
            .ltout(\U712_CHIP_RAM.N_557_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_13_4 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_13_4  (
            .in0(N__5469),
            .in1(N__5463),
            .in2(N__5442),
            .in3(N__6679),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_10_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_10_13_5 .LUT_INIT=16'b0000100010101000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_10_13_5  (
            .in0(N__8505),
            .in1(N__5411),
            .in2(N__5439),
            .in3(N__5436),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9025),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_1_LC_10_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_1_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_1_LC_10_13_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_1_LC_10_13_6  (
            .in0(N__6652),
            .in1(N__5378),
            .in2(_gnd_net_),
            .in3(N__6586),
            .lcout(\U712_CHIP_RAM.N_566 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_13_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__6861),
            .in2(_gnd_net_),
            .in3(N__6226),
            .lcout(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_14_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_14_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_14_0 .LUT_INIT=16'b1110110011101110;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_10_14_0  (
            .in0(N__5253),
            .in1(N__6350),
            .in2(N__8049),
            .in3(N__5317),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9029),
            .ce(),
            .sr(N__10228));
    defparam \U712_REG_SM.ASn_LC_10_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_LC_10_14_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_LC_10_14_1 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \U712_REG_SM.ASn_LC_10_14_1  (
            .in0(N__7017),
            .in1(N__8194),
            .in2(N__7728),
            .in3(N__5791),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9029),
            .ce(),
            .sr(N__10228));
    defparam \U712_REG_SM.REG_TACK_LC_10_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_10_14_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_10_14_2  (
            .in0(N__7880),
            .in1(N__5652),
            .in2(N__5778),
            .in3(N__5658),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9029),
            .ce(),
            .sr(N__10228));
    defparam \U712_CHIP_RAM.DBDIR_LC_10_14_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_10_14_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_10_14_3 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_10_14_3  (
            .in0(N__5748),
            .in1(N__5684),
            .in2(_gnd_net_),
            .in3(N__5715),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9029),
            .ce(),
            .sr(N__10228));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_15_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_15_2 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_15_2  (
            .in0(N__8124),
            .in1(N__7688),
            .in2(_gnd_net_),
            .in3(N__8178),
            .lcout(\U712_REG_SM.N_447 ),
            .ltout(\U712_REG_SM.N_447_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_15_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_10_15_3  (
            .in0(N__10082),
            .in1(_gnd_net_),
            .in2(N__5661),
            .in3(N__7778),
            .lcout(\U712_REG_SM.REG_TACK_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_15_6 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_10_15_6  (
            .in0(N__7779),
            .in1(N__7689),
            .in2(_gnd_net_),
            .in3(N__8179),
            .lcout(\U712_REG_SM.N_478 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_7_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_11_7_2  (
            .in0(N__5928),
            .in1(N__5934),
            .in2(_gnd_net_),
            .in3(N__5943),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9001),
            .ce(N__8891),
            .sr(N__10256));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_7_6 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_11_7_6  (
            .in0(N__9095),
            .in1(N__10641),
            .in2(N__9192),
            .in3(N__5622),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9001),
            .ce(N__8891),
            .sr(N__10256));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_11_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_11_8_0 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_11_8_0  (
            .in0(N__10291),
            .in1(N__5910),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_8_2 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_8_2  (
            .in0(N__9953),
            .in1(N__5949),
            .in2(N__9612),
            .in3(N__9759),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_8_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__7113),
            .in2(_gnd_net_),
            .in3(N__7065),
            .lcout(\U712_CHIP_RAM.N_379 ),
            .ltout(\U712_CHIP_RAM.N_379_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_8_4 .LUT_INIT=16'b0100000000001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_8_4  (
            .in0(N__9951),
            .in1(N__8858),
            .in2(N__5937),
            .in3(N__9758),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_8_7 .LUT_INIT=16'b1100111110001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_8_7  (
            .in0(N__8859),
            .in1(N__9094),
            .in2(N__9779),
            .in3(N__9952),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_9_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_9_0  (
            .in0(N__9694),
            .in1(N__7052),
            .in2(N__7212),
            .in3(N__7099),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(\U712_CHIP_RAM.REFRESH_RST_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_9_1 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_9_1  (
            .in0(N__9695),
            .in1(N__7202),
            .in2(N__5913),
            .in3(N__7100),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_9_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_9_7  (
            .in0(N__9696),
            .in1(N__5891),
            .in2(_gnd_net_),
            .in3(N__5862),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_10_0 .LUT_INIT=16'b1100000011010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_10_0  (
            .in0(N__5841),
            .in1(N__5835),
            .in2(N__7070),
            .in3(N__5958),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9009),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_10_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_10_1  (
            .in0(N__8515),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6261),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_10_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_10_5  (
            .in0(N__6422),
            .in1(N__6399),
            .in2(_gnd_net_),
            .in3(N__9717),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_11_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_10_7 .LUT_INIT=16'b0011000010110000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_11_10_7  (
            .in0(N__6381),
            .in1(N__6363),
            .in2(N__8523),
            .in3(N__6357),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9009),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_11_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__8426),
            .in2(_gnd_net_),
            .in3(N__6351),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9013),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_11_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_11_11_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_11_11_3  (
            .in0(N__6259),
            .in1(N__6457),
            .in2(_gnd_net_),
            .in3(N__7797),
            .lcout(\U712_CHIP_RAM.N_567 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIHSHE1_LC_11_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIHSHE1_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIHSHE1_LC_11_11_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIHSHE1_LC_11_11_4  (
            .in0(N__8425),
            .in1(N__6862),
            .in2(_gnd_net_),
            .in3(N__6260),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_11_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_11_11_5 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_11_11_5  (
            .in0(N__7808),
            .in1(N__6458),
            .in2(N__6246),
            .in3(N__6228),
            .lcout(\U712_CHIP_RAM.N_502 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_11_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_11_11_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_11_11_6  (
            .in0(N__6029),
            .in1(N__6498),
            .in2(N__6185),
            .in3(N__6092),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_518_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_11_7 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(N__6030),
            .in2(N__6006),
            .in3(N__5992),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_12_0 .LUT_INIT=16'b1011100011111000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_12_0  (
            .in0(N__8541),
            .in1(N__8504),
            .in2(N__6899),
            .in3(N__8640),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9016),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_11_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_11_12_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_11_12_2  (
            .in0(N__6792),
            .in1(N__6691),
            .in2(_gnd_net_),
            .in3(N__6565),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_11_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_11_12_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__9938),
            .in2(_gnd_net_),
            .in3(N__6459),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_492_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_12_4 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_12_4  (
            .in0(N__6492),
            .in1(N__7640),
            .in2(N__6462),
            .in3(N__8503),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9016),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_11_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_11_13_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_11_13_2  (
            .in0(N__7839),
            .in1(N__7770),
            .in2(_gnd_net_),
            .in3(N__8132),
            .lcout(),
            .ltout(\U712_REG_SM.STATE_COUNT_srsts_i_0_0_a2_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_13_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_13_3 .LUT_INIT=16'b0000000011110001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_11_13_3  (
            .in0(N__7771),
            .in1(N__6441),
            .in2(N__6444),
            .in3(N__7881),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9022),
            .ce(),
            .sr(N__10229));
    defparam \U712_REG_SM.C3_SYNC_RNI347S_1_LC_11_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI347S_1_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI347S_1_LC_11_13_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI347S_1_LC_11_13_4  (
            .in0(N__7701),
            .in1(N__8195),
            .in2(_gnd_net_),
            .in3(N__7807),
            .lcout(\U712_REG_SM.N_661 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_11_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_11_14_1 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_11_14_1  (
            .in0(N__10072),
            .in1(N__8089),
            .in2(_gnd_net_),
            .in3(N__8127),
            .lcout(\U712_REG_SM.DS_EN_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_14_2 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_14_2  (
            .in0(N__8125),
            .in1(N__7695),
            .in2(_gnd_net_),
            .in3(N__8188),
            .lcout(\U712_REG_SM.N_374 ),
            .ltout(\U712_REG_SM.N_374_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_14_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_14_3 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_11_14_3  (
            .in0(N__8506),
            .in1(N__7772),
            .in2(N__7020),
            .in3(N__8128),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9026),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_11_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_11_14_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__8088),
            .in2(_gnd_net_),
            .in3(N__8224),
            .lcout(\U712_REG_SM.N_389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_RNO_0_LC_11_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_RNO_0_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_RNO_0_LC_11_14_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_REG_SM.ASn_RNO_0_LC_11_14_7  (
            .in0(N__8187),
            .in1(N__8225),
            .in2(_gnd_net_),
            .in3(N__8126),
            .lcout(\U712_REG_SM.N_417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_15_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6927),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9030),
            .ce(),
            .sr(N__10226));
    defparam \U712_REG_SM.C3_SYNC_0_LC_11_15_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_11_15_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_11_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6992),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9030),
            .ce(),
            .sr(N__10226));
    defparam \U712_REG_SM.DS_EN_LC_11_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_11_15_5 .LUT_INIT=16'b1111101100000001;
    LogicCell40 \U712_REG_SM.DS_EN_LC_11_15_5  (
            .in0(N__7647),
            .in1(N__6975),
            .in2(N__8058),
            .in3(N__11054),
            .lcout(DS_ENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9030),
            .ce(),
            .sr(N__10226));
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_15_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6969),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9030),
            .ce(),
            .sr(N__10226));
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_16_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_16_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_16_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_11_16_2  (
            .in0(N__6963),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9034),
            .ce(),
            .sr(N__10225));
    defparam \U712_CHIP_RAM.RASn_LC_12_2_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_12_2_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_12_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_12_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7128),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8997),
            .ce(),
            .sr(N__10270));
    defparam \U712_CHIP_RAM.WEn_LC_12_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_12_6_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_12_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7071),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8998),
            .ce(),
            .sr(N__10253));
    defparam \U712_CHIP_RAM.CRCSn_LC_12_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_12_6_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_12_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7221),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8998),
            .ce(),
            .sr(N__10253));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_7_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_12_7_0  (
            .in0(N__7029),
            .in1(N__10374),
            .in2(N__9975),
            .in3(N__7314),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8999),
            .ce(N__8912),
            .sr(N__10247));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_7_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_12_7_2  (
            .in0(N__7028),
            .in1(N__7272),
            .in2(N__9974),
            .in3(N__7947),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8999),
            .ce(N__8912),
            .sr(N__10247));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_3 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_7_3  (
            .in0(N__9121),
            .in1(N__7545),
            .in2(N__9789),
            .in3(N__7515),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8999),
            .ce(N__8912),
            .sr(N__10247));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_7_5 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_12_7_5  (
            .in0(N__9782),
            .in1(_gnd_net_),
            .in2(N__9131),
            .in3(N__7220),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8999),
            .ce(N__8912),
            .sr(N__10247));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_7_7 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_12_7_7  (
            .in0(N__7941),
            .in1(N__9125),
            .in2(N__9193),
            .in3(N__7134),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8999),
            .ce(N__8912),
            .sr(N__10247));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_1 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_1  (
            .in0(N__7140),
            .in1(N__9781),
            .in2(N__9967),
            .in3(N__8550),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_8_3 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_8_3  (
            .in0(N__7121),
            .in1(N__9780),
            .in2(_gnd_net_),
            .in3(N__7066),
            .lcout(\U712_CHIP_RAM.CMA_5_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_12_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_12_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__7470),
            .in2(_gnd_net_),
            .in3(N__7831),
            .lcout(),
            .ltout(\U712_REG_SM.N_477_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_12_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_12_10_2 .LUT_INIT=16'b1010000010100010;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_12_10_2  (
            .in0(N__8497),
            .in1(N__7641),
            .in2(N__7611),
            .in3(N__7608),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9004),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_10_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_10_3  (
            .in0(N__7577),
            .in1(N__9936),
            .in2(_gnd_net_),
            .in3(N__8772),
            .lcout(\U712_CHIP_RAM.N_422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_10_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_10_5  (
            .in0(N__7536),
            .in1(N__9937),
            .in2(_gnd_net_),
            .in3(N__7926),
            .lcout(\U712_CHIP_RAM.N_445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_0_LC_12_11_1.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_12_11_1.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_12_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_12_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7506),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9005),
            .ce(),
            .sr(N__10230));
    defparam DBR_SYNC_1_LC_12_11_6.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_12_11_6.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_12_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_12_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7476),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9005),
            .ce(),
            .sr(N__10230));
    defparam \U712_REG_SM.START_RST_LC_12_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.START_RST_LC_12_12_4 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_REG_SM.START_RST_LC_12_12_4  (
            .in0(N__7469),
            .in1(N__7742),
            .in2(_gnd_net_),
            .in3(N__8232),
            .lcout(\U712_REG_SM.START_RSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9011),
            .ce(),
            .sr(N__10227));
    defparam \U712_CYCLE_TERM.TACK_EN_LC_12_12_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_12_12_6 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_LC_12_12_6  (
            .in0(N__7372),
            .in1(N__7455),
            .in2(_gnd_net_),
            .in3(N__7443),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9011),
            .ce(),
            .sr(N__10227));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_12_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_12_13_0 .LUT_INIT=16'b0011001100110000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__8093),
            .in2(N__7724),
            .in3(N__8197),
            .lcout(),
            .ltout(\U712_REG_SM.N_475_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_12_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_12_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_12_13_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_12_13_1  (
            .in0(N__7899),
            .in1(N__7879),
            .in2(N__7863),
            .in3(N__8494),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9014),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_57_i_LC_12_13_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_57_i_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_57_i_LC_12_13_3 .LUT_INIT=16'b0101010101000101;
    LogicCell40 \U712_BYTE_ENABLE.N_57_i_LC_12_13_3  (
            .in0(N__8565),
            .in1(N__11174),
            .in2(N__8662),
            .in3(N__8689),
            .lcout(N_57_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_12_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_12_13_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_12_13_4  (
            .in0(N__7838),
            .in1(N__8196),
            .in2(N__7723),
            .in3(N__7818),
            .lcout(\U712_REG_SM.START_RST_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_12_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_12_13_5 .LUT_INIT=16'b0001101110111011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_12_13_5  (
            .in0(N__8094),
            .in1(N__7769),
            .in2(N__7812),
            .in3(N__7716),
            .lcout(),
            .ltout(\U712_REG_SM.N_449_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_13_6 .LUT_INIT=16'b0000101000000010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_12_13_6  (
            .in0(N__8495),
            .in1(N__7712),
            .in2(N__7782),
            .in3(N__8198),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9014),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_12_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_12_14_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__7700),
            .in2(_gnd_net_),
            .in3(N__8193),
            .lcout(),
            .ltout(\U712_REG_SM.N_396_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_12_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_12_14_2 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_12_14_2  (
            .in0(N__8231),
            .in1(N__7743),
            .in2(N__7731),
            .in3(N__8496),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9018),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_12_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_12_15_4 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_2_LC_12_15_4  (
            .in0(N__8095),
            .in1(N__8226),
            .in2(N__8199),
            .in3(N__7696),
            .lcout(\U712_REG_SM.un1_STATE_COUNT_4_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_12_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_12_15_5 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_1_LC_12_15_5  (
            .in0(N__8227),
            .in1(N__8192),
            .in2(N__8133),
            .in3(N__8096),
            .lcout(\U712_REG_SM.N_479 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pll_RNI8MQ3_LC_12_16_1.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_12_16_1.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_12_16_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 pll_RNI8MQ3_LC_12_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8043),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_16_5.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_16_5.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_16_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8481),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_7_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_7_3  (
            .in0(N__10736),
            .in1(_gnd_net_),
            .in2(N__10623),
            .in3(N__10434),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10365),
            .ce(N__10331),
            .sr(N__10257));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_7_7  (
            .in0(N__10603),
            .in1(N__8280),
            .in2(_gnd_net_),
            .in3(N__8820),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10365),
            .ce(N__10331),
            .sr(N__10257));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_5  (
            .in0(N__9435),
            .in1(N__10602),
            .in2(_gnd_net_),
            .in3(N__9387),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__10330),
            .sr(N__10248));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_4  (
            .in0(N__8816),
            .in1(N__10598),
            .in2(_gnd_net_),
            .in3(N__8279),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10329),
            .sr(N__10245));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_6  (
            .in0(N__10728),
            .in1(N__10599),
            .in2(_gnd_net_),
            .in3(N__10429),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10329),
            .sr(N__10245));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_10_0 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_10_0  (
            .in0(N__9745),
            .in1(N__7908),
            .in2(N__9959),
            .in3(N__8556),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_13_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_13_10_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__9744),
            .in2(_gnd_net_),
            .in3(N__9918),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_11_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_11_3  (
            .in0(N__9588),
            .in1(N__10608),
            .in2(_gnd_net_),
            .in3(N__8809),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10326),
            .sr(N__10238));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_11_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_11_5  (
            .in0(N__9382),
            .in1(N__10609),
            .in2(_gnd_net_),
            .in3(N__8272),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10326),
            .sr(N__10238));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_13_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_13_12_1 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_13_12_1  (
            .in0(N__8492),
            .in1(N__10029),
            .in2(_gnd_net_),
            .in3(N__11170),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9017),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_12_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__8331),
            .in2(_gnd_net_),
            .in3(N__8531),
            .lcout(\U712_CHIP_RAM.un3_DMA_CYCLE_START ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_13_12_4  (
            .in0(N__8532),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8493),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9017),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_6_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_6_3  (
            .in0(N__9945),
            .in1(N__8325),
            .in2(N__9787),
            .in3(N__9627),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_14_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_14_7_2 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_14_7_2  (
            .in0(N__9112),
            .in1(N__8238),
            .in2(N__9194),
            .in3(N__8313),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9002),
            .ce(N__8908),
            .sr(N__10260));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_0  (
            .in0(N__9386),
            .in1(N__10600),
            .in2(_gnd_net_),
            .in3(N__8271),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10364),
            .ce(N__10332),
            .sr(N__10258));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_8_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_8_1  (
            .in0(N__10601),
            .in1(N__9495),
            .in2(_gnd_net_),
            .in3(N__9431),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10364),
            .ce(N__10332),
            .sr(N__10258));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_9_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_14_9_7  (
            .in0(N__9132),
            .in1(N__9597),
            .in2(N__9173),
            .in3(N__8847),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9010),
            .ce(N__8907),
            .sr(N__10249));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_11_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_11_1  (
            .in0(N__9587),
            .in1(N__10545),
            .in2(_gnd_net_),
            .in3(N__8795),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10363),
            .ce(N__10327),
            .sr(N__10244));
    defparam \U712_BYTE_ENABLE.N_295_i_LC_14_12_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_295_i_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_295_i_LC_14_12_2 .LUT_INIT=16'b0101000101010101;
    LogicCell40 \U712_BYTE_ENABLE.N_295_i_LC_14_12_2  (
            .in0(N__8574),
            .in1(N__8706),
            .in2(N__10028),
            .in3(N__8655),
            .lcout(N_295_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_299_i_LC_14_12_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_299_i_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_299_i_LC_14_12_6 .LUT_INIT=16'b0011001100100011;
    LogicCell40 \U712_BYTE_ENABLE.N_299_i_LC_14_12_6  (
            .in0(N__10024),
            .in1(N__9309),
            .in2(N__8664),
            .in3(N__8708),
            .lcout(N_299_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_297_i_LC_14_12_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_297_i_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_297_i_LC_14_12_7 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \U712_BYTE_ENABLE.N_297_i_LC_14_12_7  (
            .in0(N__8707),
            .in1(N__9315),
            .in2(N__8663),
            .in3(N__11169),
            .lcout(N_297_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_13_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_13_2 .LUT_INIT=16'b0000101000101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_13_2  (
            .in0(N__9963),
            .in1(N__10950),
            .in2(N__9300),
            .in3(N__10873),
            .lcout(\U712_BYTE_ENABLE.N_528 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_o2_LC_14_13_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_o2_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_o2_LC_14_13_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_LDSn_i_o2_LC_14_13_3  (
            .in0(N__10874),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10781),
            .lcout(\U712_BYTE_ENABLE.N_377 ),
            .ltout(\U712_BYTE_ENABLE.N_377_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_14_13_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_14_13_4 .LUT_INIT=16'b1000000010101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_14_13_4  (
            .in0(N__9961),
            .in1(N__10948),
            .in2(N__8568),
            .in3(N__9295),
            .lcout(\U712_BYTE_ENABLE.N_508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_14_13_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_14_13_6 .LUT_INIT=16'b0010000010101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_14_13_6  (
            .in0(N__9962),
            .in1(N__10949),
            .in2(N__9324),
            .in3(N__9296),
            .lcout(\U712_BYTE_ENABLE.N_530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_14_14_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_14_14_0 .LUT_INIT=16'b0101110100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_14_14_0  (
            .in0(N__9294),
            .in1(N__10947),
            .in2(N__10882),
            .in3(N__9966),
            .lcout(\U712_BYTE_ENABLE.N_532 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_i_x2_LC_14_17_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_i_x2_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_i_x2_LC_14_17_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_i_x2_LC_14_17_4  (
            .in0(N__11023),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10780),
            .lcout(\U712_BYTE_ENABLE.N_364_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_14_20_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_14_20_5 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_14_20_5  (
            .in0(N__10020),
            .in1(N__11178),
            .in2(_gnd_net_),
            .in3(N__11255),
            .lcout(DMA_LATCH_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_403_i_LC_14_20_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_403_i_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_403_i_LC_14_20_7 .LUT_INIT=16'b0000111011100000;
    LogicCell40 \U712_BYTE_ENABLE.N_403_i_LC_14_20_7  (
            .in0(N__10935),
            .in1(N__10883),
            .in2(N__11014),
            .in3(N__10779),
            .lcout(N_403_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CASn_LC_15_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_15_4_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_15_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_15_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9788),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9000),
            .ce(),
            .sr(N__10272));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_15_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_15_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_15_6_0 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_15_6_0  (
            .in0(N__9333),
            .in1(N__9127),
            .in2(N__9195),
            .in3(N__9633),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9003),
            .ce(N__8913),
            .sr(N__10269));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_15_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_15_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_15_6_6 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_15_6_6  (
            .in0(N__9191),
            .in1(N__9126),
            .in2(N__9447),
            .in3(N__9069),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9003),
            .ce(N__8913),
            .sr(N__10269));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_7_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_7_3  (
            .in0(N__9960),
            .in1(N__9798),
            .in2(N__9786),
            .in3(N__9618),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_8_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_8_2  (
            .in0(N__10611),
            .in1(N__10737),
            .in2(_gnd_net_),
            .in3(N__10685),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__10335),
            .sr(N__10261));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_8_5  (
            .in0(N__10612),
            .in1(N__9494),
            .in2(_gnd_net_),
            .in3(N__9430),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__10335),
            .sr(N__10261));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_9_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_9_5  (
            .in0(N__10684),
            .in1(N__10610),
            .in2(_gnd_net_),
            .in3(N__9486),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__10333),
            .sr(N__10259));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_11_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_11_1  (
            .in0(N__9543),
            .in1(N__10572),
            .in2(_gnd_net_),
            .in3(N__9586),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10360),
            .ce(N__10328),
            .sr(N__10246));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_13_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_15_13_3  (
            .in0(N__9582),
            .in1(N__10607),
            .in2(_gnd_net_),
            .in3(N__9539),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10334),
            .sr(N__10239));
    defparam \U712_BYTE_ENABLE.N_402_i_LC_15_20_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_402_i_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_402_i_LC_15_20_3 .LUT_INIT=16'b0000110111010000;
    LogicCell40 \U712_BYTE_ENABLE.N_402_i_LC_15_20_3  (
            .in0(N__10936),
            .in1(N__10884),
            .in2(N__11024),
            .in3(N__10802),
            .lcout(N_402_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_2  (
            .in0(N__9493),
            .in1(_gnd_net_),
            .in2(N__10628),
            .in3(N__10680),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10361),
            .ce(N__10336),
            .sr(N__10268));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_8_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_8_4  (
            .in0(N__10619),
            .in1(N__9429),
            .in2(_gnd_net_),
            .in3(N__9369),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10361),
            .ce(N__10336),
            .sr(N__10268));
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_16_19_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_16_19_7 .LUT_INIT=16'b0010100011111111;
    LogicCell40 \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_16_19_7  (
            .in0(N__10864),
            .in1(N__10986),
            .in2(N__10815),
            .in3(N__11069),
            .lcout(N_291),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_400_i_LC_16_20_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_400_i_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_400_i_LC_16_20_0 .LUT_INIT=16'b0000101110100000;
    LogicCell40 \U712_BYTE_ENABLE.N_400_i_LC_16_20_0  (
            .in0(N__10933),
            .in1(N__10865),
            .in2(N__10811),
            .in3(N__11018),
            .lcout(N_400_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_20_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_20_5 .LUT_INIT=16'b0001000011111111;
    LogicCell40 \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_20_5  (
            .in0(N__10869),
            .in1(N__10807),
            .in2(N__11025),
            .in3(N__11073),
            .lcout(N_293),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_401_i_LC_16_20_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_401_i_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_401_i_LC_16_20_7 .LUT_INIT=16'b0001000100101010;
    LogicCell40 \U712_BYTE_ENABLE.N_401_i_LC_16_20_7  (
            .in0(N__11019),
            .in1(N__10934),
            .in2(N__10881),
            .in3(N__10806),
            .lcout(N_401_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_7_1  (
            .in0(N__10550),
            .in1(N__10729),
            .in2(_gnd_net_),
            .in3(N__10686),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10362),
            .ce(N__10337),
            .sr(N__10271));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_19_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_19_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_19_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_19_7_7  (
            .in0(N__10549),
            .in1(N__10449),
            .in2(_gnd_net_),
            .in3(N__10433),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10359),
            .ce(N__10338),
            .sr(N__10273));
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_20_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_20_2 .LUT_INIT=16'b0010000000100000;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_20_2  (
            .in0(N__11156),
            .in1(N__10140),
            .in2(N__10019),
            .in3(_gnd_net_),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_24_20_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_24_20_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_24_20_5 .LUT_INIT=16'b0100011100001111;
    LogicCell40 \U712_BUFFERS.DRDDIR_0_m2_LC_24_20_5  (
            .in0(N__10086),
            .in1(N__10004),
            .in2(N__11262),
            .in3(N__11155),
            .lcout(N_450),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

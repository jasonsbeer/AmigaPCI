// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 19 2024 10:10:35

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U111_TOP" view "INTERFACE"

module U111_TOP (
    D_LL_AMIGA,
    D_LM_AMIGA,
    D_UU_AMIGA,
    D_UM_AMIGA,
    D_UU_040,
    D_LL_040,
    D_LM_040,
    D_UM_040,
    A_AMIGA,
    A_040,
    SIZ,
    TSn,
    RESETn,
    CLKRAMA,
    PORTSIZE,
    CLK40B,
    TBI_CPUn,
    TAn,
    CPUBGn,
    BUFENn,
    RnW,
    CLK80_CPU,
    BUFDIR,
    TCI_CPUn,
    TS_CPUn,
    CLKRAMB,
    CLK40A,
    DMAn,
    CLK40C,
    CLK40_IN,
    TACKn,
    BGn);

    inout [7:0] D_LL_AMIGA;
    inout [7:0] D_LM_AMIGA;
    inout [7:0] D_UU_AMIGA;
    inout [7:0] D_UM_AMIGA;
    inout [7:0] D_UU_040;
    inout [7:0] D_LL_040;
    inout [7:0] D_LM_040;
    inout [7:0] D_UM_040;
    output [1:0] A_AMIGA;
    input [1:0] A_040;
    input [1:0] SIZ;
    output TSn;
    input RESETn;
    output CLKRAMA;
    input PORTSIZE;
    output CLK40B;
    output TBI_CPUn;
    output TAn;
    output CPUBGn;
    output BUFENn;
    input RnW;
    output CLK80_CPU;
    output BUFDIR;
    output TCI_CPUn;
    input TS_CPUn;
    output CLKRAMB;
    output CLK40A;
    output DMAn;
    output CLK40C;
    input CLK40_IN;
    input TACKn;
    input BGn;

    wire N__8230;
    wire N__8214;
    wire N__8213;
    wire N__8212;
    wire N__8205;
    wire N__8204;
    wire N__8203;
    wire N__8196;
    wire N__8195;
    wire N__8194;
    wire N__8187;
    wire N__8186;
    wire N__8185;
    wire N__8178;
    wire N__8177;
    wire N__8176;
    wire N__8169;
    wire N__8168;
    wire N__8167;
    wire N__8160;
    wire N__8159;
    wire N__8158;
    wire N__8151;
    wire N__8150;
    wire N__8149;
    wire N__8142;
    wire N__8141;
    wire N__8140;
    wire N__8133;
    wire N__8132;
    wire N__8131;
    wire N__8124;
    wire N__8123;
    wire N__8122;
    wire N__8115;
    wire N__8114;
    wire N__8113;
    wire N__8106;
    wire N__8105;
    wire N__8104;
    wire N__8097;
    wire N__8096;
    wire N__8095;
    wire N__8088;
    wire N__8087;
    wire N__8086;
    wire N__8079;
    wire N__8078;
    wire N__8077;
    wire N__8070;
    wire N__8069;
    wire N__8068;
    wire N__8061;
    wire N__8060;
    wire N__8059;
    wire N__8052;
    wire N__8051;
    wire N__8050;
    wire N__8043;
    wire N__8042;
    wire N__8041;
    wire N__8034;
    wire N__8033;
    wire N__8032;
    wire N__8025;
    wire N__8024;
    wire N__8023;
    wire N__8016;
    wire N__8015;
    wire N__8014;
    wire N__8007;
    wire N__8006;
    wire N__8005;
    wire N__7998;
    wire N__7997;
    wire N__7996;
    wire N__7989;
    wire N__7988;
    wire N__7987;
    wire N__7980;
    wire N__7979;
    wire N__7978;
    wire N__7971;
    wire N__7970;
    wire N__7969;
    wire N__7962;
    wire N__7961;
    wire N__7960;
    wire N__7953;
    wire N__7952;
    wire N__7951;
    wire N__7944;
    wire N__7943;
    wire N__7942;
    wire N__7935;
    wire N__7934;
    wire N__7933;
    wire N__7926;
    wire N__7925;
    wire N__7924;
    wire N__7917;
    wire N__7916;
    wire N__7915;
    wire N__7908;
    wire N__7907;
    wire N__7906;
    wire N__7899;
    wire N__7898;
    wire N__7897;
    wire N__7890;
    wire N__7889;
    wire N__7888;
    wire N__7881;
    wire N__7880;
    wire N__7879;
    wire N__7872;
    wire N__7871;
    wire N__7870;
    wire N__7863;
    wire N__7862;
    wire N__7861;
    wire N__7854;
    wire N__7853;
    wire N__7852;
    wire N__7845;
    wire N__7844;
    wire N__7843;
    wire N__7836;
    wire N__7835;
    wire N__7834;
    wire N__7827;
    wire N__7826;
    wire N__7825;
    wire N__7818;
    wire N__7817;
    wire N__7816;
    wire N__7809;
    wire N__7808;
    wire N__7807;
    wire N__7800;
    wire N__7799;
    wire N__7798;
    wire N__7791;
    wire N__7790;
    wire N__7789;
    wire N__7782;
    wire N__7781;
    wire N__7780;
    wire N__7773;
    wire N__7772;
    wire N__7771;
    wire N__7764;
    wire N__7763;
    wire N__7762;
    wire N__7755;
    wire N__7754;
    wire N__7753;
    wire N__7746;
    wire N__7745;
    wire N__7744;
    wire N__7737;
    wire N__7736;
    wire N__7735;
    wire N__7728;
    wire N__7727;
    wire N__7726;
    wire N__7719;
    wire N__7718;
    wire N__7717;
    wire N__7710;
    wire N__7709;
    wire N__7708;
    wire N__7701;
    wire N__7700;
    wire N__7699;
    wire N__7692;
    wire N__7691;
    wire N__7690;
    wire N__7683;
    wire N__7682;
    wire N__7681;
    wire N__7674;
    wire N__7673;
    wire N__7672;
    wire N__7665;
    wire N__7664;
    wire N__7663;
    wire N__7656;
    wire N__7655;
    wire N__7654;
    wire N__7647;
    wire N__7646;
    wire N__7645;
    wire N__7638;
    wire N__7637;
    wire N__7636;
    wire N__7629;
    wire N__7628;
    wire N__7627;
    wire N__7620;
    wire N__7619;
    wire N__7618;
    wire N__7611;
    wire N__7610;
    wire N__7609;
    wire N__7602;
    wire N__7601;
    wire N__7600;
    wire N__7593;
    wire N__7592;
    wire N__7591;
    wire N__7584;
    wire N__7583;
    wire N__7582;
    wire N__7575;
    wire N__7574;
    wire N__7573;
    wire N__7566;
    wire N__7565;
    wire N__7564;
    wire N__7557;
    wire N__7556;
    wire N__7555;
    wire N__7548;
    wire N__7547;
    wire N__7546;
    wire N__7539;
    wire N__7538;
    wire N__7537;
    wire N__7530;
    wire N__7529;
    wire N__7528;
    wire N__7521;
    wire N__7520;
    wire N__7519;
    wire N__7512;
    wire N__7511;
    wire N__7510;
    wire N__7503;
    wire N__7502;
    wire N__7501;
    wire N__7494;
    wire N__7493;
    wire N__7492;
    wire N__7485;
    wire N__7484;
    wire N__7483;
    wire N__7476;
    wire N__7475;
    wire N__7474;
    wire N__7467;
    wire N__7466;
    wire N__7465;
    wire N__7458;
    wire N__7457;
    wire N__7456;
    wire N__7449;
    wire N__7448;
    wire N__7447;
    wire N__7440;
    wire N__7439;
    wire N__7438;
    wire N__7431;
    wire N__7430;
    wire N__7429;
    wire N__7422;
    wire N__7421;
    wire N__7420;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7393;
    wire N__7390;
    wire N__7389;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7374;
    wire N__7371;
    wire N__7368;
    wire N__7363;
    wire N__7360;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7345;
    wire N__7340;
    wire N__7339;
    wire N__7338;
    wire N__7335;
    wire N__7334;
    wire N__7333;
    wire N__7332;
    wire N__7331;
    wire N__7326;
    wire N__7325;
    wire N__7324;
    wire N__7323;
    wire N__7322;
    wire N__7321;
    wire N__7318;
    wire N__7317;
    wire N__7316;
    wire N__7315;
    wire N__7308;
    wire N__7305;
    wire N__7304;
    wire N__7301;
    wire N__7296;
    wire N__7293;
    wire N__7288;
    wire N__7287;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7275;
    wire N__7270;
    wire N__7267;
    wire N__7258;
    wire N__7253;
    wire N__7252;
    wire N__7251;
    wire N__7248;
    wire N__7243;
    wire N__7238;
    wire N__7233;
    wire N__7230;
    wire N__7227;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7192;
    wire N__7191;
    wire N__7190;
    wire N__7189;
    wire N__7188;
    wire N__7185;
    wire N__7182;
    wire N__7179;
    wire N__7176;
    wire N__7173;
    wire N__7170;
    wire N__7165;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7145;
    wire N__7144;
    wire N__7143;
    wire N__7140;
    wire N__7139;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7125;
    wire N__7122;
    wire N__7119;
    wire N__7116;
    wire N__7111;
    wire N__7108;
    wire N__7105;
    wire N__7100;
    wire N__7093;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7081;
    wire N__7080;
    wire N__7077;
    wire N__7074;
    wire N__7071;
    wire N__7068;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7047;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7035;
    wire N__7032;
    wire N__7027;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6997;
    wire N__6996;
    wire N__6993;
    wire N__6990;
    wire N__6987;
    wire N__6984;
    wire N__6981;
    wire N__6978;
    wire N__6975;
    wire N__6970;
    wire N__6967;
    wire N__6964;
    wire N__6961;
    wire N__6958;
    wire N__6953;
    wire N__6950;
    wire N__6947;
    wire N__6944;
    wire N__6941;
    wire N__6938;
    wire N__6935;
    wire N__6932;
    wire N__6929;
    wire N__6926;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6911;
    wire N__6910;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6900;
    wire N__6895;
    wire N__6892;
    wire N__6889;
    wire N__6886;
    wire N__6883;
    wire N__6880;
    wire N__6877;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6839;
    wire N__6838;
    wire N__6835;
    wire N__6832;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6819;
    wire N__6814;
    wire N__6811;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6769;
    wire N__6766;
    wire N__6763;
    wire N__6762;
    wire N__6759;
    wire N__6756;
    wire N__6753;
    wire N__6750;
    wire N__6745;
    wire N__6742;
    wire N__6739;
    wire N__6736;
    wire N__6733;
    wire N__6730;
    wire N__6727;
    wire N__6722;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6710;
    wire N__6707;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6682;
    wire N__6681;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6663;
    wire N__6658;
    wire N__6655;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6617;
    wire N__6614;
    wire N__6611;
    wire N__6608;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6596;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6586;
    wire N__6583;
    wire N__6582;
    wire N__6579;
    wire N__6576;
    wire N__6573;
    wire N__6570;
    wire N__6567;
    wire N__6564;
    wire N__6561;
    wire N__6558;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6544;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6507;
    wire N__6502;
    wire N__6499;
    wire N__6494;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6467;
    wire N__6464;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6456;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6416;
    wire N__6413;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6385;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6375;
    wire N__6372;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6328;
    wire N__6327;
    wire N__6326;
    wire N__6323;
    wire N__6322;
    wire N__6321;
    wire N__6318;
    wire N__6317;
    wire N__6316;
    wire N__6311;
    wire N__6308;
    wire N__6303;
    wire N__6302;
    wire N__6299;
    wire N__6296;
    wire N__6293;
    wire N__6292;
    wire N__6291;
    wire N__6290;
    wire N__6289;
    wire N__6288;
    wire N__6285;
    wire N__6284;
    wire N__6279;
    wire N__6276;
    wire N__6271;
    wire N__6270;
    wire N__6269;
    wire N__6268;
    wire N__6267;
    wire N__6266;
    wire N__6265;
    wire N__6262;
    wire N__6257;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6247;
    wire N__6246;
    wire N__6245;
    wire N__6244;
    wire N__6241;
    wire N__6238;
    wire N__6237;
    wire N__6234;
    wire N__6231;
    wire N__6230;
    wire N__6229;
    wire N__6226;
    wire N__6221;
    wire N__6218;
    wire N__6213;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6188;
    wire N__6185;
    wire N__6184;
    wire N__6179;
    wire N__6176;
    wire N__6171;
    wire N__6168;
    wire N__6165;
    wire N__6164;
    wire N__6163;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6144;
    wire N__6139;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6123;
    wire N__6118;
    wire N__6115;
    wire N__6110;
    wire N__6109;
    wire N__6106;
    wire N__6101;
    wire N__6098;
    wire N__6089;
    wire N__6086;
    wire N__6077;
    wire N__6074;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6050;
    wire N__6047;
    wire N__6044;
    wire N__6041;
    wire N__6040;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__5998;
    wire N__5993;
    wire N__5992;
    wire N__5989;
    wire N__5986;
    wire N__5985;
    wire N__5984;
    wire N__5983;
    wire N__5978;
    wire N__5971;
    wire N__5970;
    wire N__5969;
    wire N__5968;
    wire N__5967;
    wire N__5966;
    wire N__5961;
    wire N__5958;
    wire N__5957;
    wire N__5956;
    wire N__5955;
    wire N__5950;
    wire N__5949;
    wire N__5946;
    wire N__5945;
    wire N__5942;
    wire N__5941;
    wire N__5940;
    wire N__5935;
    wire N__5930;
    wire N__5927;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5919;
    wire N__5914;
    wire N__5913;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5887;
    wire N__5884;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5874;
    wire N__5871;
    wire N__5868;
    wire N__5865;
    wire N__5864;
    wire N__5861;
    wire N__5860;
    wire N__5859;
    wire N__5854;
    wire N__5853;
    wire N__5852;
    wire N__5851;
    wire N__5846;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5834;
    wire N__5833;
    wire N__5826;
    wire N__5823;
    wire N__5820;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5806;
    wire N__5803;
    wire N__5798;
    wire N__5797;
    wire N__5796;
    wire N__5795;
    wire N__5790;
    wire N__5787;
    wire N__5784;
    wire N__5779;
    wire N__5770;
    wire N__5765;
    wire N__5762;
    wire N__5757;
    wire N__5754;
    wire N__5751;
    wire N__5746;
    wire N__5743;
    wire N__5732;
    wire N__5723;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5705;
    wire N__5702;
    wire N__5701;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5686;
    wire N__5683;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5633;
    wire N__5632;
    wire N__5631;
    wire N__5630;
    wire N__5629;
    wire N__5628;
    wire N__5627;
    wire N__5626;
    wire N__5625;
    wire N__5624;
    wire N__5623;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5583;
    wire N__5580;
    wire N__5577;
    wire N__5574;
    wire N__5571;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5545;
    wire N__5544;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5532;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5522;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5503;
    wire N__5502;
    wire N__5501;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5489;
    wire N__5486;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5459;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5447;
    wire N__5446;
    wire N__5445;
    wire N__5444;
    wire N__5441;
    wire N__5434;
    wire N__5431;
    wire N__5426;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5401;
    wire N__5400;
    wire N__5399;
    wire N__5398;
    wire N__5397;
    wire N__5396;
    wire N__5395;
    wire N__5394;
    wire N__5391;
    wire N__5386;
    wire N__5381;
    wire N__5372;
    wire N__5363;
    wire N__5362;
    wire N__5361;
    wire N__5358;
    wire N__5357;
    wire N__5356;
    wire N__5355;
    wire N__5354;
    wire N__5351;
    wire N__5350;
    wire N__5347;
    wire N__5346;
    wire N__5343;
    wire N__5338;
    wire N__5333;
    wire N__5324;
    wire N__5315;
    wire N__5314;
    wire N__5313;
    wire N__5312;
    wire N__5311;
    wire N__5310;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5296;
    wire N__5291;
    wire N__5288;
    wire N__5287;
    wire N__5278;
    wire N__5275;
    wire N__5270;
    wire N__5267;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5238;
    wire N__5237;
    wire N__5236;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5224;
    wire N__5223;
    wire N__5222;
    wire N__5221;
    wire N__5220;
    wire N__5217;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5194;
    wire N__5193;
    wire N__5190;
    wire N__5189;
    wire N__5188;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5166;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5158;
    wire N__5157;
    wire N__5156;
    wire N__5155;
    wire N__5154;
    wire N__5153;
    wire N__5146;
    wire N__5145;
    wire N__5142;
    wire N__5139;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5115;
    wire N__5114;
    wire N__5113;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5105;
    wire N__5100;
    wire N__5099;
    wire N__5098;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5066;
    wire N__5063;
    wire N__5062;
    wire N__5061;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5040;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5023;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5010;
    wire N__5007;
    wire N__4996;
    wire N__4993;
    wire N__4990;
    wire N__4987;
    wire N__4982;
    wire N__4977;
    wire N__4972;
    wire N__4969;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4945;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4930;
    wire N__4927;
    wire N__4924;
    wire N__4921;
    wire N__4918;
    wire N__4915;
    wire N__4912;
    wire N__4909;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4868;
    wire N__4867;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4822;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4795;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4732;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4666;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4573;
    wire N__4570;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4558;
    wire N__4555;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4543;
    wire N__4540;
    wire N__4537;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4483;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4465;
    wire N__4462;
    wire N__4459;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4423;
    wire N__4420;
    wire N__4417;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4393;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4375;
    wire N__4372;
    wire N__4369;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4212;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4145;
    wire N__4144;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4129;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4117;
    wire N__4114;
    wire N__4111;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4066;
    wire N__4063;
    wire N__4060;
    wire N__4057;
    wire N__4054;
    wire N__4051;
    wire N__4048;
    wire N__4045;
    wire N__4042;
    wire N__4039;
    wire N__4036;
    wire N__4033;
    wire N__4030;
    wire N__4027;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__4000;
    wire N__3997;
    wire N__3994;
    wire N__3991;
    wire N__3988;
    wire N__3985;
    wire N__3982;
    wire N__3979;
    wire N__3976;
    wire N__3973;
    wire N__3970;
    wire N__3967;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3953;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3941;
    wire N__3938;
    wire N__3935;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3914;
    wire N__3911;
    wire N__3908;
    wire N__3905;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3887;
    wire N__3884;
    wire N__3881;
    wire N__3878;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3845;
    wire N__3842;
    wire N__3839;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3817;
    wire N__3814;
    wire N__3811;
    wire N__3808;
    wire N__3805;
    wire N__3802;
    wire N__3799;
    wire N__3796;
    wire N__3793;
    wire N__3788;
    wire N__3785;
    wire N__3782;
    wire N__3779;
    wire N__3776;
    wire N__3773;
    wire N__3770;
    wire N__3767;
    wire N__3764;
    wire N__3761;
    wire N__3758;
    wire N__3755;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3730;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3680;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3668;
    wire N__3665;
    wire N__3662;
    wire N__3661;
    wire N__3658;
    wire N__3655;
    wire N__3652;
    wire N__3649;
    wire N__3646;
    wire N__3643;
    wire N__3640;
    wire N__3637;
    wire N__3634;
    wire N__3631;
    wire N__3628;
    wire N__3625;
    wire N__3622;
    wire N__3617;
    wire N__3614;
    wire N__3611;
    wire N__3608;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire N__3596;
    wire N__3593;
    wire N__3590;
    wire N__3587;
    wire N__3584;
    wire N__3581;
    wire N__3578;
    wire N__3575;
    wire N__3572;
    wire N__3569;
    wire N__3566;
    wire N__3563;
    wire N__3560;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3548;
    wire N__3545;
    wire N__3542;
    wire N__3539;
    wire N__3536;
    wire N__3533;
    wire N__3530;
    wire N__3527;
    wire N__3524;
    wire N__3521;
    wire N__3518;
    wire N__3515;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire N__3497;
    wire N__3494;
    wire N__3491;
    wire N__3488;
    wire N__3485;
    wire N__3482;
    wire N__3479;
    wire N__3476;
    wire N__3473;
    wire N__3470;
    wire N__3467;
    wire N__3464;
    wire N__3461;
    wire N__3458;
    wire N__3455;
    wire N__3452;
    wire N__3449;
    wire N__3446;
    wire N__3443;
    wire N__3440;
    wire N__3437;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3425;
    wire N__3422;
    wire N__3419;
    wire N__3416;
    wire N__3413;
    wire N__3412;
    wire N__3409;
    wire N__3406;
    wire N__3403;
    wire N__3400;
    wire N__3397;
    wire N__3394;
    wire N__3391;
    wire N__3388;
    wire N__3385;
    wire N__3382;
    wire N__3377;
    wire N__3374;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3362;
    wire N__3359;
    wire N__3356;
    wire N__3353;
    wire N__3350;
    wire N__3347;
    wire N__3344;
    wire N__3341;
    wire N__3338;
    wire N__3335;
    wire N__3332;
    wire N__3329;
    wire N__3326;
    wire N__3323;
    wire N__3320;
    wire N__3317;
    wire N__3314;
    wire N__3311;
    wire N__3308;
    wire N__3305;
    wire N__3302;
    wire N__3299;
    wire N__3296;
    wire N__3293;
    wire N__3290;
    wire N__3287;
    wire N__3284;
    wire N__3281;
    wire N__3278;
    wire N__3275;
    wire N__3272;
    wire N__3269;
    wire N__3266;
    wire N__3263;
    wire N__3260;
    wire N__3257;
    wire N__3254;
    wire N__3251;
    wire N__3248;
    wire N__3245;
    wire N__3242;
    wire N__3239;
    wire N__3236;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3190;
    wire N__3187;
    wire N__3184;
    wire N__3179;
    wire N__3176;
    wire N__3173;
    wire N__3170;
    wire N__3167;
    wire N__3164;
    wire N__3163;
    wire N__3160;
    wire N__3157;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3121;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3104;
    wire N__3101;
    wire N__3098;
    wire N__3095;
    wire N__3092;
    wire N__3089;
    wire N__3086;
    wire N__3083;
    wire N__3080;
    wire N__3077;
    wire N__3076;
    wire N__3073;
    wire N__3070;
    wire N__3067;
    wire N__3064;
    wire N__3061;
    wire N__3058;
    wire N__3055;
    wire N__3052;
    wire N__3049;
    wire N__3046;
    wire N__3043;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3031;
    wire N__3026;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3011;
    wire N__3008;
    wire N__3005;
    wire N__3002;
    wire N__2999;
    wire N__2996;
    wire N__2993;
    wire N__2990;
    wire N__2987;
    wire N__2984;
    wire N__2981;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2966;
    wire N__2963;
    wire N__2960;
    wire N__2957;
    wire N__2956;
    wire N__2953;
    wire N__2950;
    wire N__2947;
    wire N__2944;
    wire N__2941;
    wire N__2938;
    wire N__2935;
    wire N__2932;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2920;
    wire N__2917;
    wire N__2914;
    wire N__2909;
    wire N__2906;
    wire N__2903;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2888;
    wire N__2885;
    wire N__2882;
    wire N__2879;
    wire N__2876;
    wire N__2873;
    wire N__2870;
    wire N__2867;
    wire N__2864;
    wire N__2861;
    wire N__2858;
    wire N__2857;
    wire N__2854;
    wire N__2851;
    wire N__2848;
    wire N__2845;
    wire N__2842;
    wire N__2839;
    wire N__2836;
    wire N__2833;
    wire N__2830;
    wire N__2827;
    wire N__2822;
    wire N__2819;
    wire N__2816;
    wire N__2813;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2795;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2780;
    wire N__2777;
    wire N__2776;
    wire N__2773;
    wire N__2770;
    wire N__2767;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2755;
    wire N__2752;
    wire N__2749;
    wire N__2746;
    wire N__2743;
    wire N__2740;
    wire N__2737;
    wire N__2732;
    wire N__2729;
    wire N__2726;
    wire N__2723;
    wire N__2720;
    wire N__2717;
    wire N__2714;
    wire N__2711;
    wire N__2708;
    wire N__2705;
    wire N__2702;
    wire N__2699;
    wire N__2696;
    wire N__2693;
    wire N__2690;
    wire N__2689;
    wire N__2686;
    wire N__2683;
    wire N__2682;
    wire N__2681;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2669;
    wire N__2668;
    wire N__2661;
    wire N__2658;
    wire N__2655;
    wire N__2648;
    wire N__2647;
    wire N__2646;
    wire N__2645;
    wire N__2644;
    wire N__2643;
    wire N__2642;
    wire N__2639;
    wire N__2636;
    wire N__2635;
    wire N__2634;
    wire N__2633;
    wire N__2632;
    wire N__2631;
    wire N__2630;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2620;
    wire N__2617;
    wire N__2614;
    wire N__2609;
    wire N__2606;
    wire N__2603;
    wire N__2600;
    wire N__2597;
    wire N__2596;
    wire N__2595;
    wire N__2594;
    wire N__2593;
    wire N__2590;
    wire N__2587;
    wire N__2584;
    wire N__2575;
    wire N__2574;
    wire N__2573;
    wire N__2570;
    wire N__2569;
    wire N__2568;
    wire N__2567;
    wire N__2556;
    wire N__2553;
    wire N__2550;
    wire N__2547;
    wire N__2544;
    wire N__2535;
    wire N__2532;
    wire N__2529;
    wire N__2526;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2516;
    wire N__2515;
    wire N__2508;
    wire N__2497;
    wire N__2494;
    wire N__2491;
    wire N__2490;
    wire N__2489;
    wire N__2484;
    wire N__2481;
    wire N__2478;
    wire N__2473;
    wire N__2468;
    wire N__2465;
    wire N__2462;
    wire N__2459;
    wire N__2456;
    wire N__2453;
    wire N__2450;
    wire N__2447;
    wire N__2442;
    wire N__2439;
    wire N__2434;
    wire N__2429;
    wire N__2426;
    wire N__2417;
    wire N__2414;
    wire N__2411;
    wire N__2408;
    wire N__2405;
    wire N__2402;
    wire N__2399;
    wire N__2396;
    wire N__2393;
    wire N__2390;
    wire N__2387;
    wire N__2384;
    wire N__2381;
    wire N__2378;
    wire N__2375;
    wire N__2372;
    wire N__2369;
    wire N__2366;
    wire N__2363;
    wire N__2360;
    wire N__2357;
    wire N__2354;
    wire N__2351;
    wire N__2348;
    wire N__2345;
    wire N__2342;
    wire N__2339;
    wire N__2336;
    wire N__2333;
    wire N__2330;
    wire N__2327;
    wire N__2324;
    wire N__2321;
    wire N__2318;
    wire N__2315;
    wire N__2312;
    wire N__2309;
    wire N__2306;
    wire N__2303;
    wire N__2300;
    wire N__2297;
    wire N__2294;
    wire N__2291;
    wire N__2288;
    wire N__2285;
    wire N__2282;
    wire N__2279;
    wire N__2276;
    wire N__2275;
    wire N__2272;
    wire N__2269;
    wire N__2266;
    wire N__2263;
    wire N__2260;
    wire N__2257;
    wire N__2254;
    wire N__2251;
    wire N__2248;
    wire N__2245;
    wire N__2242;
    wire N__2239;
    wire N__2236;
    wire N__2233;
    wire N__2228;
    wire N__2225;
    wire N__2222;
    wire N__2219;
    wire N__2216;
    wire N__2213;
    wire VCCG0;
    wire GNDG0;
    wire A_040_c_0;
    wire A_AMIGA_c_0;
    wire A_040_c_1;
    wire A_AMIGA_c_1_cascade_;
    wire D_LL_AMIGA_in_3;
    wire un1_D_LL_AMIGA_3;
    wire D_LL_AMIGA_in_4;
    wire un1_D_LL_AMIGA_4;
    wire D_UM_040_in_0;
    wire D_LL_040_in_0;
    wire un1_D_UM_040_0;
    wire D_UM_040_in_2;
    wire D_LL_040_in_2;
    wire un1_D_UM_040_2;
    wire D_LL_040_in_1;
    wire D_UM_040_in_1;
    wire un1_D_UM_040_1;
    wire D_LL_040_in_7;
    wire D_UM_040_in_7;
    wire un1_D_UM_040_7;
    wire D_UU_040_in_1;
    wire D_LM_040_in_1;
    wire un1_D_UU_040_1;
    wire D_LM_AMIGA_in_3;
    wire un1_D_LM_AMIGA_3;
    wire D_LM_040_in_7;
    wire D_UU_040_in_7;
    wire un1_D_UU_040_7;
    wire D_LM_040_in_3;
    wire D_UU_040_in_3;
    wire un1_D_UU_040_3;
    wire RnW_c_i_0;
    wire D_LL_AMIGA_in_6;
    wire un1_D_LL_AMIGA_6;
    wire D_LM_AMIGA_in_5;
    wire un1_D_LM_AMIGA_5;
    wire D_LM_AMIGA_in_7;
    wire un1_D_LM_AMIGA_7;
    wire TSn_c;
    wire \INVU111_CYCLE_SM.TSnC_net ;
    wire D_LL_AMIGA_in_0;
    wire un1_D_LL_AMIGA_0;
    wire D_UU_040_in_4;
    wire D_LM_040_in_4;
    wire un1_D_UU_040_4;
    wire D_LL_AMIGA_in_1;
    wire un1_D_LL_AMIGA_1;
    wire D_LL_AMIGA_in_2;
    wire un1_D_LL_AMIGA_2;
    wire D_LM_AMIGA_in_0;
    wire un1_D_LM_AMIGA_0;
    wire D_UU_040_in_2;
    wire D_LM_040_in_2;
    wire un1_D_UU_040_2;
    wire D_UU_040_in_0;
    wire D_LM_040_in_0;
    wire un1_D_UU_040_0;
    wire D_LL_040_in_4;
    wire D_UM_040_in_4;
    wire un1_D_UM_040_4;
    wire D_LM_AMIGA_in_2;
    wire un1_D_LM_AMIGA_2;
    wire D_LM_AMIGA_in_6;
    wire un1_D_LM_AMIGA_6;
    wire D_UM_040_in_3;
    wire D_LL_040_in_3;
    wire un1_D_UM_040_3;
    wire D_UU_040_in_5;
    wire D_LM_040_in_5;
    wire un1_D_UU_040_5;
    wire D_UM_040_in_5;
    wire D_LL_040_in_5;
    wire un1_D_UM_040_5;
    wire D_LL_AMIGA_in_5;
    wire un1_D_LL_AMIGA_5;
    wire D_LL_AMIGA_in_7;
    wire un1_D_LL_AMIGA_7;
    wire un1_D_UM_AMIGA_2;
    wire \INVU111_CYCLE_SM.TA_ENC_net ;
    wire \U111_CYCLE_SM.RESETn_c_i ;
    wire D_UM_AMIGA_in_2;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_2C_net ;
    wire \U111_CYCLE_SM.un3_LW_CYCLE_START_cascade_ ;
    wire TS_CPUn_c;
    wire \U111_CYCLE_SM.N_69_0_cascade_ ;
    wire \U111_CYCLE_SM.TS_EN_5 ;
    wire \U111_CYCLE_SM.TS_ENZ0 ;
    wire \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net ;
    wire \INVU111_CYCLE_SM.UU_LATCHED_nesr_6C_net ;
    wire PORTSIZE_c;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire CONSTANT_ONE_NET;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ;
    wire D_UU_AMIGA_in_3;
    wire un1_D_UU_AMIGA_3;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ;
    wire D_UU_AMIGA_in_6;
    wire un1_D_UU_AMIGA_6;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ;
    wire D_UU_AMIGA_in_2;
    wire un1_D_UU_AMIGA_2;
    wire GB_BUFFER_CLK40_THRU_CO;
    wire D_LM_AMIGA_in_1;
    wire un1_D_LM_AMIGA_1;
    wire D_UM_040_in_6;
    wire D_LL_040_in_6;
    wire un1_D_UM_040_6;
    wire \U111_CYCLE_SM.TA_ENZ0 ;
    wire U111_CYCLE_SM_TAn_0_i;
    wire D_LM_AMIGA_in_4;
    wire un1_D_LM_AMIGA_4;
    wire \INVU111_CYCLE_SM.LW_CYCLEC_net ;
    wire \U111_CYCLE_SM.LW_CYCLE_0 ;
    wire \U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0 ;
    wire CLK40;
    wire \U111_CYCLE_SM.N_91_cascade_ ;
    wire \U111_CYCLE_SM.LW_CYCLE_STARTZ0 ;
    wire \U111_CYCLE_SM.A_OUT_0_cascade_ ;
    wire \U111_CYCLE_SM.A_OUTZ0 ;
    wire \INVU111_CYCLE_SM.CYCLE_STATE_0C_net ;
    wire TACKn_c;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ;
    wire RESETn_c;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_ ;
    wire RnW_c;
    wire \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa ;
    wire \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net ;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ;
    wire D_UU_AMIGA_in_0;
    wire un1_D_UU_AMIGA_0;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ;
    wire D_UM_AMIGA_in_5;
    wire un1_D_UM_AMIGA_5;
    wire \U111_CYCLE_SM.un1_LW_TRANS_1_0 ;
    wire D_UU_040_in_6;
    wire D_LM_040_in_6;
    wire A_AMIGA_c_1;
    wire un1_D_UU_040_6;
    wire D_UU_AMIGA_in_4;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ;
    wire un1_D_UU_AMIGA_4;
    wire CLK80;
    wire GB_BUFFER_CLK80_THRU_CO;
    wire un1_D_UM_AMIGA_0;
    wire un1_D_UM_AMIGA_6;
    wire D_UM_AMIGA_in_6;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ;
    wire D_UM_AMIGA_in_0;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net ;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_1C_net ;
    wire \INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net ;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ;
    wire \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0 ;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ;
    wire D_UM_AMIGA_in_3;
    wire un1_D_UM_AMIGA_3;
    wire D_UM_AMIGA_in_1;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ;
    wire un1_D_UM_AMIGA_1;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ;
    wire D_UU_AMIGA_in_1;
    wire un1_D_UU_AMIGA_1;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ;
    wire D_UM_AMIGA_in_4;
    wire un1_D_UM_AMIGA_4;
    wire D_UM_AMIGA_in_7;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ;
    wire un1_D_UM_AMIGA_7;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ;
    wire D_UU_AMIGA_in_7;
    wire un1_D_UU_AMIGA_7;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ;
    wire D_UU_AMIGA_in_5;
    wire \U111_CYCLE_SM.LW_CYCLEZ0 ;
    wire un1_D_UU_AMIGA_5;
    wire _gnd_net_;

    defparam pll_pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll_pll.TEST_MODE=1'b0;
    defparam pll_pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll_pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll_pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll_pll.FILTER_RANGE=3'b011;
    defparam pll_pll.FEEDBACK_PATH="SIMPLE";
    defparam pll_pll.FDA_RELATIVE=4'b0000;
    defparam pll_pll.FDA_FEEDBACK=4'b0000;
    defparam pll_pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll_pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll_pll.DIVR=4'b0000;
    defparam pll_pll.DIVQ=3'b011;
    defparam pll_pll.DIVF=7'b0001111;
    defparam pll_pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40_2F pll_pll (
            .SCLK(),
            .PLLOUTGLOBALA(CLK80),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALB(CLK40),
            .SDI(),
            .PLLOUTCOREA(),
            .BYPASS(),
            .RESETB(N__4458),
            .PLLOUTCOREB(),
            .LOCK(),
            .SDO(),
            .EXTFEEDBACK(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__8230));
    IO_PAD pll_iopad (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__8230),
            .PACKAGEPIN(CLK40_IN));
    defparam D_UM_040_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_3_iopad (
            .OE(N__8214),
            .DIN(N__8213),
            .DOUT(N__8212),
            .PACKAGEPIN(D_UM_040[3]));
    defparam D_UM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_3_preio (
            .PADOEN(N__8214),
            .PADOUT(N__8213),
            .PADIN(N__8212),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5114),
            .DIN0(D_UM_040_in_3),
            .DOUT0(N__7022),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_1_iopad (
            .OE(N__8205),
            .DIN(N__8204),
            .DOUT(N__8203),
            .PACKAGEPIN(D_LL_AMIGA[1]));
    defparam D_LL_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_1_preio (
            .PADOEN(N__8205),
            .PADOUT(N__8204),
            .PADIN(N__8203),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2682),
            .DIN0(D_LL_AMIGA_in_1),
            .DOUT0(N__3163),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_5_iopad (
            .OE(N__8196),
            .DIN(N__8195),
            .DOUT(N__8194),
            .PACKAGEPIN(D_UU_AMIGA[5]));
    defparam D_UU_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_5_preio (
            .PADOEN(N__8196),
            .PADOUT(N__8195),
            .PADIN(N__8194),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2630),
            .DIN0(D_UU_AMIGA_in_5),
            .DOUT0(N__3707),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_ibuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_ibuf_iopad (
            .OE(N__8187),
            .DIN(N__8186),
            .DOUT(N__8185),
            .PACKAGEPIN(TACKn));
    defparam TACKn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TACKn_ibuf_preio (
            .PADOEN(N__8187),
            .PADOUT(N__8186),
            .PADIN(N__8185),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TACKn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_6_iopad (
            .OE(N__8178),
            .DIN(N__8177),
            .DOUT(N__8176),
            .PACKAGEPIN(D_UU_040[6]));
    defparam D_UU_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_6_preio (
            .PADOEN(N__8178),
            .PADOUT(N__8177),
            .PADIN(N__8176),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5158),
            .DIN0(D_UU_040_in_6),
            .DOUT0(N__4904),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam CPUBGn_obuf_iopad.PULLUP=1'b1;
    IO_PAD CPUBGn_obuf_iopad (
            .OE(N__8169),
            .DIN(N__8168),
            .DOUT(N__8167),
            .PACKAGEPIN(CPUBGn));
    defparam CPUBGn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUBGn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CPUBGn_obuf_preio (
            .PADOEN(N__8169),
            .PADOUT(N__8168),
            .PADIN(N__8167),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_7_iopad (
            .OE(N__8160),
            .DIN(N__8159),
            .DOUT(N__8158),
            .PACKAGEPIN(D_LL_040[7]));
    defparam D_LL_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_7_preio (
            .PADOEN(N__8160),
            .PADOUT(N__8159),
            .PADIN(N__8158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5220),
            .DIN0(D_LL_040_in_7),
            .DOUT0(N__4283),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_4_iopad (
            .OE(N__8151),
            .DIN(N__8150),
            .DOUT(N__8149),
            .PACKAGEPIN(D_LL_AMIGA[4]));
    defparam D_LL_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_4_preio (
            .PADOEN(N__8151),
            .PADOUT(N__8150),
            .PADIN(N__8149),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2681),
            .DIN0(D_LL_AMIGA_in_4),
            .DOUT0(N__4004),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_3_iopad (
            .OE(N__8142),
            .DIN(N__8141),
            .DOUT(N__8140),
            .PACKAGEPIN(D_UM_AMIGA[3]));
    defparam D_UM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_3_preio (
            .PADOEN(N__8142),
            .PADOUT(N__8141),
            .PADIN(N__8140),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2574),
            .DIN0(D_UM_AMIGA_in_3),
            .DOUT0(N__3788),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_3_iopad (
            .OE(N__8133),
            .DIN(N__8132),
            .DOUT(N__8131),
            .PACKAGEPIN(D_UU_040[3]));
    defparam D_UU_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_3_preio (
            .PADOEN(N__8133),
            .PADOUT(N__8132),
            .PADIN(N__8131),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5153),
            .DIN0(D_UU_040_in_3),
            .DOUT0(N__4361),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_1_iopad (
            .OE(N__8124),
            .DIN(N__8123),
            .DOUT(N__8122),
            .PACKAGEPIN(A_040[1]));
    defparam A_040_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_1_preio (
            .PADOEN(N__8124),
            .PADOUT(N__8123),
            .PADIN(N__8122),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_3_iopad (
            .OE(N__8115),
            .DIN(N__8114),
            .DOUT(N__8113),
            .PACKAGEPIN(D_LM_AMIGA[3]));
    defparam D_LM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_3_preio (
            .PADOEN(N__8115),
            .PADOUT(N__8114),
            .PADIN(N__8113),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2647),
            .DIN0(D_LM_AMIGA_in_3),
            .DOUT0(N__2780),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_0_iopad (
            .OE(N__8106),
            .DIN(N__8105),
            .DOUT(N__8104),
            .PACKAGEPIN(D_LM_040[0]));
    defparam D_LM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_0_preio (
            .PADOEN(N__8106),
            .PADOUT(N__8105),
            .PADIN(N__8104),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5221),
            .DIN0(D_LM_040_in_0),
            .DOUT0(N__3260),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_6_iopad (
            .OE(N__8097),
            .DIN(N__8096),
            .DOUT(N__8095),
            .PACKAGEPIN(D_UM_AMIGA[6]));
    defparam D_UM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_6_preio (
            .PADOEN(N__8097),
            .PADOUT(N__8096),
            .PADIN(N__8095),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2629),
            .DIN0(D_UM_AMIGA_in_6),
            .DOUT0(N__4685),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_4_iopad (
            .OE(N__8088),
            .DIN(N__8087),
            .DOUT(N__8086),
            .PACKAGEPIN(D_LM_AMIGA[4]));
    defparam D_LM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_4_preio (
            .PADOEN(N__8088),
            .PADOUT(N__8087),
            .PADIN(N__8086),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2632),
            .DIN0(D_LM_AMIGA_in_4),
            .DOUT0(N__3419),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_1_iopad (
            .OE(N__8079),
            .DIN(N__8078),
            .DOUT(N__8077),
            .PACKAGEPIN(A_AMIGA[1]));
    defparam A_AMIGA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_1_preio (
            .PADOEN(N__8079),
            .PADOUT(N__8078),
            .PADIN(N__8077),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5833),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_7_iopad (
            .OE(N__8070),
            .DIN(N__8069),
            .DOUT(N__8068),
            .PACKAGEPIN(D_LM_040[7]));
    defparam D_LM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_7_preio (
            .PADOEN(N__8070),
            .PADOUT(N__8069),
            .PADIN(N__8068),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5039),
            .DIN0(D_LM_040_in_7),
            .DOUT0(N__3500),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_4_iopad (
            .OE(N__8061),
            .DIN(N__8060),
            .DOUT(N__8059),
            .PACKAGEPIN(D_UM_040[4]));
    defparam D_UM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_4_preio (
            .PADOEN(N__8061),
            .PADOUT(N__8060),
            .PADIN(N__8059),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5154),
            .DIN0(D_UM_040_in_4),
            .DOUT0(N__6794),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_obuf_iopad (
            .OE(N__8052),
            .DIN(N__8051),
            .DOUT(N__8050),
            .PACKAGEPIN(CLK40B));
    defparam CLK40B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_obuf_preio (
            .PADOEN(N__8052),
            .PADOUT(N__8051),
            .PADIN(N__8050),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4823),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_0_iopad (
            .OE(N__8043),
            .DIN(N__8042),
            .DOUT(N__8041),
            .PACKAGEPIN(D_UU_AMIGA[0]));
    defparam D_UU_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_0_preio (
            .PADOEN(N__8043),
            .PADOUT(N__8042),
            .PADIN(N__8041),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2644),
            .DIN0(D_UU_AMIGA_in_0),
            .DOUT0(N__4022),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_0_iopad (
            .OE(N__8034),
            .DIN(N__8033),
            .DOUT(N__8032),
            .PACKAGEPIN(A_040[0]));
    defparam A_040_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_0_preio (
            .PADOEN(N__8034),
            .PADOUT(N__8033),
            .PADIN(N__8032),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_0_iopad (
            .OE(N__8025),
            .DIN(N__8024),
            .DOUT(N__8023),
            .PACKAGEPIN(D_LM_AMIGA[0]));
    defparam D_LM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_0_preio (
            .PADOEN(N__8025),
            .PADOUT(N__8024),
            .PADIN(N__8023),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2569),
            .DIN0(D_LM_AMIGA_in_0),
            .DOUT0(N__4070),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_1_iopad (
            .OE(N__8016),
            .DIN(N__8015),
            .DOUT(N__8014),
            .PACKAGEPIN(D_UM_040[1]));
    defparam D_UM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_1_preio (
            .PADOEN(N__8016),
            .PADOUT(N__8015),
            .PADIN(N__8014),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5112),
            .DIN0(D_UM_040_in_1),
            .DOUT0(N__6944),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBI_CPUn_obuf_iopad (
            .OE(N__8007),
            .DIN(N__8006),
            .DOUT(N__8005),
            .PACKAGEPIN(TBI_CPUn));
    defparam TBI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TBI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TBI_CPUn_obuf_preio (
            .PADOEN(N__8007),
            .PADOUT(N__8006),
            .PADIN(N__8005),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40A_obuf_iopad (
            .OE(N__7998),
            .DIN(N__7997),
            .DOUT(N__7996),
            .PACKAGEPIN(CLK40A));
    defparam CLK40A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40A_obuf_preio (
            .PADOEN(N__7998),
            .PADOUT(N__7997),
            .PADIN(N__7996),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4822),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_3_iopad (
            .OE(N__7989),
            .DIN(N__7988),
            .DOUT(N__7987),
            .PACKAGEPIN(D_LM_040[3]));
    defparam D_LM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_3_preio (
            .PADOEN(N__7989),
            .PADOUT(N__7988),
            .PADIN(N__7987),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5145),
            .DIN0(D_LM_040_in_3),
            .DOUT0(N__2885),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_4_iopad (
            .OE(N__7980),
            .DIN(N__7979),
            .DOUT(N__7978),
            .PACKAGEPIN(D_LL_040[4]));
    defparam D_LL_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_4_preio (
            .PADOEN(N__7980),
            .PADOUT(N__7979),
            .PADIN(N__7978),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5238),
            .DIN0(D_LL_040_in_4),
            .DOUT0(N__2318),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_7_iopad (
            .OE(N__7971),
            .DIN(N__7970),
            .DOUT(N__7969),
            .PACKAGEPIN(D_LL_AMIGA[7]));
    defparam D_LL_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_7_preio (
            .PADOEN(N__7971),
            .PADOUT(N__7970),
            .PADIN(N__7969),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2568),
            .DIN0(D_LL_AMIGA_in_7),
            .DOUT0(N__3077),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_7_iopad (
            .OE(N__7962),
            .DIN(N__7961),
            .DOUT(N__7960),
            .PACKAGEPIN(D_UU_AMIGA[7]));
    defparam D_UU_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_7_preio (
            .PADOEN(N__7962),
            .PADOUT(N__7961),
            .PADIN(N__7960),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2642),
            .DIN0(D_UU_AMIGA_in_7),
            .DOUT0(N__2798),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFDIR_obuf_iopad (
            .OE(N__7953),
            .DIN(N__7952),
            .DOUT(N__7951),
            .PACKAGEPIN(BUFDIR));
    defparam BUFDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFDIR_obuf_preio (
            .PADOEN(N__7953),
            .PADOUT(N__7952),
            .PADIN(N__7951),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5236),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_5_iopad (
            .OE(N__7944),
            .DIN(N__7943),
            .DOUT(N__7942),
            .PACKAGEPIN(D_LM_AMIGA[5]));
    defparam D_LM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_5_preio (
            .PADOEN(N__7944),
            .PADOUT(N__7943),
            .PADIN(N__7942),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2595),
            .DIN0(D_LM_AMIGA_in_5),
            .DOUT0(N__3743),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_4_iopad (
            .OE(N__7935),
            .DIN(N__7934),
            .DOUT(N__7933),
            .PACKAGEPIN(D_UU_040[4]));
    defparam D_UU_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_4_preio (
            .PADOEN(N__7935),
            .PADOUT(N__7934),
            .PADIN(N__7933),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5189),
            .DIN0(D_UU_040_in_4),
            .DOUT0(N__5660),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SIZ_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__7926),
            .DIN(N__7925),
            .DOUT(N__7924),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__7926),
            .PADOUT(N__7925),
            .PADIN(N__7924),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_6_iopad (
            .OE(N__7917),
            .DIN(N__7916),
            .DOUT(N__7915),
            .PACKAGEPIN(D_LM_040[6]));
    defparam D_LM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_6_preio (
            .PADOEN(N__7917),
            .PADOUT(N__7916),
            .PADIN(N__7915),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5022),
            .DIN0(D_LM_040_in_6),
            .DOUT0(N__3872),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_5_iopad (
            .OE(N__7908),
            .DIN(N__7907),
            .DOUT(N__7906),
            .PACKAGEPIN(D_UM_040[5]));
    defparam D_UM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_5_preio (
            .PADOEN(N__7908),
            .PADOUT(N__7907),
            .PADIN(N__7906),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5155),
            .DIN0(D_UM_040_in_5),
            .DOUT0(N__6347),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TS_CPUn_ibuf_iopad (
            .OE(N__7899),
            .DIN(N__7898),
            .DOUT(N__7897),
            .PACKAGEPIN(TS_CPUn));
    defparam TS_CPUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TS_CPUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TS_CPUn_ibuf_preio (
            .PADOEN(N__7899),
            .PADOUT(N__7898),
            .PADIN(N__7897),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TS_CPUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_1_iopad (
            .OE(N__7890),
            .DIN(N__7889),
            .DOUT(N__7888),
            .PACKAGEPIN(D_LL_040[1]));
    defparam D_LL_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_1_preio (
            .PADOEN(N__7890),
            .PADOUT(N__7889),
            .PADIN(N__7888),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5237),
            .DIN0(D_LL_040_in_1),
            .DOUT0(N__3341),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_3_iopad (
            .OE(N__7881),
            .DIN(N__7880),
            .DOUT(N__7879),
            .PACKAGEPIN(D_LL_AMIGA[3]));
    defparam D_LL_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_3_preio (
            .PADOEN(N__7881),
            .PADOUT(N__7880),
            .PADIN(N__7879),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2689),
            .DIN0(D_LL_AMIGA_in_3),
            .DOUT0(N__3830),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_5_iopad (
            .OE(N__7872),
            .DIN(N__7871),
            .DOUT(N__7870),
            .PACKAGEPIN(D_UM_AMIGA[5]));
    defparam D_UM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_5_preio (
            .PADOEN(N__7872),
            .PADOUT(N__7871),
            .PADIN(N__7870),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2645),
            .DIN0(D_UM_AMIGA_in_5),
            .DOUT0(N__3614),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_1_iopad (
            .OE(N__7863),
            .DIN(N__7862),
            .DOUT(N__7861),
            .PACKAGEPIN(D_UU_040[1]));
    defparam D_UU_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_1_preio (
            .PADOEN(N__7863),
            .PADOUT(N__7862),
            .PADIN(N__7861),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5115),
            .DIN0(D_UU_040_in_1),
            .DOUT0(N__6872),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_3_iopad (
            .OE(N__7854),
            .DIN(N__7853),
            .DOUT(N__7852),
            .PACKAGEPIN(D_UU_AMIGA[3]));
    defparam D_UU_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_3_preio (
            .PADOEN(N__7854),
            .PADOUT(N__7853),
            .PADIN(N__7852),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2631),
            .DIN0(D_UU_AMIGA_in_3),
            .DOUT0(N__2708),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_1_iopad (
            .OE(N__7845),
            .DIN(N__7844),
            .DOUT(N__7843),
            .PACKAGEPIN(D_LM_AMIGA[1]));
    defparam D_LM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_1_preio (
            .PADOEN(N__7845),
            .PADOUT(N__7844),
            .PADIN(N__7843),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2515),
            .DIN0(D_LM_AMIGA_in_1),
            .DOUT0(N__2956),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_2_iopad (
            .OE(N__7836),
            .DIN(N__7835),
            .DOUT(N__7834),
            .PACKAGEPIN(D_LM_040[2]));
    defparam D_LM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_2_preio (
            .PADOEN(N__7836),
            .PADOUT(N__7835),
            .PADIN(N__7834),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5194),
            .DIN0(D_LM_040_in_2),
            .DOUT0(N__3905),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_5_iopad (
            .OE(N__7827),
            .DIN(N__7826),
            .DOUT(N__7825),
            .PACKAGEPIN(D_LL_040[5]));
    defparam D_LL_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_5_preio (
            .PADOEN(N__7827),
            .PADOUT(N__7826),
            .PADIN(N__7825),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5222),
            .DIN0(D_LL_040_in_5),
            .DOUT0(N__4319),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_6_iopad (
            .OE(N__7818),
            .DIN(N__7817),
            .DOUT(N__7816),
            .PACKAGEPIN(D_LL_AMIGA[6]));
    defparam D_LL_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_6_preio (
            .PADOEN(N__7818),
            .PADOUT(N__7817),
            .PADIN(N__7816),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2668),
            .DIN0(D_LL_AMIGA_in_6),
            .DOUT0(N__4736),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_6_iopad (
            .OE(N__7809),
            .DIN(N__7808),
            .DOUT(N__7807),
            .PACKAGEPIN(D_UU_AMIGA[6]));
    defparam D_UU_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_6_preio (
            .PADOEN(N__7809),
            .PADOUT(N__7808),
            .PADIN(N__7807),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2646),
            .DIN0(D_UU_AMIGA_in_6),
            .DOUT0(N__5723),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_1_iopad (
            .OE(N__7800),
            .DIN(N__7799),
            .DOUT(N__7798),
            .PACKAGEPIN(D_UM_AMIGA[1]));
    defparam D_UM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_1_preio (
            .PADOEN(N__7800),
            .PADOUT(N__7799),
            .PADIN(N__7798),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2596),
            .DIN0(D_UM_AMIGA_in_1),
            .DOUT0(N__3092),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_5_iopad (
            .OE(N__7791),
            .DIN(N__7790),
            .DOUT(N__7789),
            .PACKAGEPIN(D_UU_040[5]));
    defparam D_UU_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_5_preio (
            .PADOEN(N__7791),
            .PADOUT(N__7790),
            .PADIN(N__7789),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5156),
            .DIN0(D_UU_040_in_5),
            .DOUT0(N__7214),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMA_obuf_iopad (
            .OE(N__7782),
            .DIN(N__7781),
            .DOUT(N__7780),
            .PACKAGEPIN(CLKRAMA));
    defparam CLKRAMA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMA_obuf_preio (
            .PADOEN(N__7782),
            .PADOUT(N__7781),
            .PADIN(N__7780),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5597),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_2_iopad (
            .OE(N__7773),
            .DIN(N__7772),
            .DOUT(N__7771),
            .PACKAGEPIN(D_UM_040[2]));
    defparam D_UM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_2_preio (
            .PADOEN(N__7773),
            .PADOUT(N__7772),
            .PADIN(N__7771),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5060),
            .DIN0(D_UM_040_in_2),
            .DOUT0(N__4262),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_2_iopad (
            .OE(N__7764),
            .DIN(N__7763),
            .DOUT(N__7762),
            .PACKAGEPIN(D_LL_040[2]));
    defparam D_LL_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_2_preio (
            .PADOEN(N__7764),
            .PADOUT(N__7763),
            .PADIN(N__7762),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5224),
            .DIN0(D_LL_040_in_2),
            .DOUT0(N__3299),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TCI_CPUn_obuf_iopad.PULLUP=1'b1;
    IO_PAD TCI_CPUn_obuf_iopad (
            .OE(N__7755),
            .DIN(N__7754),
            .DOUT(N__7753),
            .PACKAGEPIN(TCI_CPUn));
    defparam TCI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TCI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TCI_CPUn_obuf_preio (
            .PADOEN(N__7755),
            .PADOUT(N__7754),
            .PADIN(N__7753),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4466),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMB_obuf_iopad (
            .OE(N__7746),
            .DIN(N__7745),
            .DOUT(N__7744),
            .PACKAGEPIN(CLKRAMB));
    defparam CLKRAMB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMB_obuf_preio (
            .PADOEN(N__7746),
            .PADOUT(N__7745),
            .PADIN(N__7744),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5583),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_2_iopad (
            .OE(N__7737),
            .DIN(N__7736),
            .DOUT(N__7735),
            .PACKAGEPIN(D_LL_AMIGA[2]));
    defparam D_LL_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_2_preio (
            .PADOEN(N__7737),
            .PADOUT(N__7736),
            .PADIN(N__7735),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2690),
            .DIN0(D_LL_AMIGA_in_2),
            .DOUT0(N__3226),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_4_iopad (
            .OE(N__7728),
            .DIN(N__7727),
            .DOUT(N__7726),
            .PACKAGEPIN(D_UM_AMIGA[4]));
    defparam D_UM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_4_preio (
            .PADOEN(N__7728),
            .PADOUT(N__7727),
            .PADIN(N__7726),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2594),
            .DIN0(D_UM_AMIGA_in_4),
            .DOUT0(N__3938),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_2_iopad (
            .OE(N__7719),
            .DIN(N__7718),
            .DOUT(N__7717),
            .PACKAGEPIN(D_UU_AMIGA[2]));
    defparam D_UU_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_2_preio (
            .PADOEN(N__7719),
            .PADOUT(N__7718),
            .PADIN(N__7717),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2643),
            .DIN0(D_UU_AMIGA_in_2),
            .DOUT0(N__4106),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__7710),
            .DIN(N__7709),
            .DOUT(N__7708),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__7710),
            .PADOUT(N__7709),
            .PADIN(N__7708),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_6_iopad (
            .OE(N__7701),
            .DIN(N__7700),
            .DOUT(N__7699),
            .PACKAGEPIN(D_LM_AMIGA[6]));
    defparam D_LM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_6_preio (
            .PADOEN(N__7701),
            .PADOUT(N__7700),
            .PADIN(N__7699),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2490),
            .DIN0(D_LM_AMIGA_in_6),
            .DOUT0(N__6041),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam RnW_ibuf_iopad.PULLUP=1'b1;
    IO_PAD RnW_ibuf_iopad (
            .OE(N__7692),
            .DIN(N__7691),
            .DOUT(N__7690),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__7692),
            .PADOUT(N__7691),
            .PADIN(N__7690),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_5_iopad (
            .OE(N__7683),
            .DIN(N__7682),
            .DOUT(N__7681),
            .PACKAGEPIN(D_LM_040[5]));
    defparam D_LM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_5_preio (
            .PADOEN(N__7683),
            .PADOUT(N__7682),
            .PADIN(N__7681),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5062),
            .DIN0(D_LM_040_in_5),
            .DOUT0(N__3539),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_6_iopad (
            .OE(N__7674),
            .DIN(N__7673),
            .DOUT(N__7672),
            .PACKAGEPIN(D_UM_040[6]));
    defparam D_UM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_6_preio (
            .PADOEN(N__7674),
            .PADOUT(N__7673),
            .PADIN(N__7672),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5023),
            .DIN0(D_UM_040_in_6),
            .DOUT0(N__6608),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TAn_obuf_iopad.PULLUP=1'b1;
    IO_PAD TAn_obuf_iopad (
            .OE(N__7665),
            .DIN(N__7664),
            .DOUT(N__7663),
            .PACKAGEPIN(TAn));
    defparam TAn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TAn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TAn_obuf_preio (
            .PADOEN(N__7665),
            .PADOUT(N__7664),
            .PADIN(N__7663),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4652),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMAn_obuf_iopad (
            .OE(N__7656),
            .DIN(N__7655),
            .DOUT(N__7654),
            .PACKAGEPIN(DMAn));
    defparam DMAn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMAn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMAn_obuf_preio (
            .PADOEN(N__7656),
            .PADOUT(N__7655),
            .PADIN(N__7654),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4465),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_6_iopad (
            .OE(N__7647),
            .DIN(N__7646),
            .DOUT(N__7645),
            .PACKAGEPIN(D_LL_040[6]));
    defparam D_LL_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_6_preio (
            .PADOEN(N__7647),
            .PADOUT(N__7646),
            .PADIN(N__7645),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5223),
            .DIN0(D_LL_040_in_6),
            .DOUT0(N__3578),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_5_iopad (
            .OE(N__7638),
            .DIN(N__7637),
            .DOUT(N__7636),
            .PACKAGEPIN(D_LL_AMIGA[5]));
    defparam D_LL_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_5_preio (
            .PADOEN(N__7638),
            .PADOUT(N__7637),
            .PADIN(N__7636),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2669),
            .DIN0(D_LL_AMIGA_in_5),
            .DOUT0(N__3662),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_0_iopad (
            .OE(N__7629),
            .DIN(N__7628),
            .DOUT(N__7627),
            .PACKAGEPIN(D_UM_AMIGA[0]));
    defparam D_UM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_0_preio (
            .PADOEN(N__7629),
            .PADOUT(N__7628),
            .PADIN(N__7627),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2635),
            .DIN0(D_UM_AMIGA_in_0),
            .DOUT0(N__2228),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_2_iopad (
            .OE(N__7620),
            .DIN(N__7619),
            .DOUT(N__7618),
            .PACKAGEPIN(D_UU_040[2]));
    defparam D_UU_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_2_preio (
            .PADOEN(N__7620),
            .PADOUT(N__7619),
            .PADIN(N__7618),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5188),
            .DIN0(D_UU_040_in_2),
            .DOUT0(N__4838),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_2_iopad (
            .OE(N__7611),
            .DIN(N__7610),
            .DOUT(N__7609),
            .PACKAGEPIN(D_LM_AMIGA[2]));
    defparam D_LM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_2_preio (
            .PADOEN(N__7611),
            .PADOUT(N__7610),
            .PADIN(N__7609),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2634),
            .DIN0(D_LM_AMIGA_in_2),
            .DOUT0(N__4144),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK80_CPU_obuf_iopad (
            .OE(N__7602),
            .DIN(N__7601),
            .DOUT(N__7600),
            .PACKAGEPIN(CLK80_CPU));
    defparam CLK80_CPU_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK80_CPU_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK80_CPU_obuf_preio (
            .PADOEN(N__7602),
            .PADOUT(N__7601),
            .PADIN(N__7600),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5593),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_3_iopad (
            .OE(N__7593),
            .DIN(N__7592),
            .DOUT(N__7591),
            .PACKAGEPIN(D_LL_040[3]));
    defparam D_LL_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_3_preio (
            .PADOEN(N__7593),
            .PADOUT(N__7592),
            .PADIN(N__7591),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5245),
            .DIN0(D_LL_040_in_3),
            .DOUT0(N__2357),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_1_iopad (
            .OE(N__7584),
            .DIN(N__7583),
            .DOUT(N__7582),
            .PACKAGEPIN(D_LM_040[1]));
    defparam D_LM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_1_preio (
            .PADOEN(N__7584),
            .PADOUT(N__7583),
            .PADIN(N__7582),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5193),
            .DIN0(D_LM_040_in_1),
            .DOUT0(N__4775),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TSn_obuf_iopad.PULLUP=1'b1;
    IO_PAD TSn_obuf_iopad (
            .OE(N__7575),
            .DIN(N__7574),
            .DOUT(N__7573),
            .PACKAGEPIN(TSn));
    defparam TSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TSn_obuf_preio (
            .PADOEN(N__7575),
            .PADOUT(N__7574),
            .PADIN(N__7573),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3485),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_7_iopad (
            .OE(N__7566),
            .DIN(N__7565),
            .DOUT(N__7564),
            .PACKAGEPIN(D_UM_AMIGA[7]));
    defparam D_UM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_7_preio (
            .PADOEN(N__7566),
            .PADOUT(N__7565),
            .PADIN(N__7564),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2593),
            .DIN0(D_UM_AMIGA_in_7),
            .DOUT0(N__2999),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_7_iopad (
            .OE(N__7557),
            .DIN(N__7556),
            .DOUT(N__7555),
            .PACKAGEPIN(D_LM_AMIGA[7]));
    defparam D_LM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_7_preio (
            .PADOEN(N__7557),
            .PADOUT(N__7556),
            .PADIN(N__7555),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2489),
            .DIN0(D_LM_AMIGA_in_7),
            .DOUT0(N__2864),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PORTSIZE_ibuf_iopad.PULLUP=1'b1;
    IO_PAD PORTSIZE_ibuf_iopad (
            .OE(N__7548),
            .DIN(N__7547),
            .DOUT(N__7546),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PORTSIZE_ibuf_preio (
            .PADOEN(N__7548),
            .PADOUT(N__7547),
            .PADIN(N__7546),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PORTSIZE_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_0_iopad (
            .OE(N__7539),
            .DIN(N__7538),
            .DOUT(N__7537),
            .PACKAGEPIN(A_AMIGA[0]));
    defparam A_AMIGA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_0_preio (
            .PADOEN(N__7539),
            .PADOUT(N__7538),
            .PADIN(N__7537),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2402),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_4_iopad (
            .OE(N__7530),
            .DIN(N__7529),
            .DOUT(N__7528),
            .PACKAGEPIN(D_LM_040[4]));
    defparam D_LM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_4_preio (
            .PADOEN(N__7530),
            .PADOUT(N__7529),
            .PADIN(N__7528),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5105),
            .DIN0(D_LM_040_in_4),
            .DOUT0(N__4613),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_7_iopad (
            .OE(N__7521),
            .DIN(N__7520),
            .DOUT(N__7519),
            .PACKAGEPIN(D_UM_040[7]));
    defparam D_UM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_7_preio (
            .PADOEN(N__7521),
            .PADOUT(N__7520),
            .PADIN(N__7519),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5113),
            .DIN0(D_UM_040_in_7),
            .DOUT0(N__6713),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__7512),
            .DIN(N__7511),
            .DOUT(N__7510),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__7512),
            .PADOUT(N__7511),
            .PADIN(N__7510),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_1_iopad (
            .OE(N__7503),
            .DIN(N__7502),
            .DOUT(N__7501),
            .PACKAGEPIN(D_UU_AMIGA[1]));
    defparam D_UU_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_1_preio (
            .PADOEN(N__7503),
            .PADOUT(N__7502),
            .PADIN(N__7501),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2573),
            .DIN0(D_UU_AMIGA_in_1),
            .DOUT0(N__2909),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__7494),
            .DIN(N__7493),
            .DOUT(N__7492),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__7494),
            .PADOUT(N__7493),
            .PADIN(N__7492),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4821),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_0_iopad (
            .OE(N__7485),
            .DIN(N__7484),
            .DOUT(N__7483),
            .PACKAGEPIN(D_UM_040[0]));
    defparam D_UM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_0_preio (
            .PADOEN(N__7485),
            .PADOUT(N__7484),
            .PADIN(N__7483),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5061),
            .DIN0(D_UM_040_in_0),
            .DOUT0(N__6629),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_0_iopad (
            .OE(N__7476),
            .DIN(N__7475),
            .DOUT(N__7474),
            .PACKAGEPIN(D_LL_AMIGA[0]));
    defparam D_LL_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_0_preio (
            .PADOEN(N__7476),
            .PADOUT(N__7475),
            .PADIN(N__7474),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2567),
            .DIN0(D_LL_AMIGA_in_0),
            .DOUT0(N__2275),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_4_iopad (
            .OE(N__7467),
            .DIN(N__7466),
            .DOUT(N__7465),
            .PACKAGEPIN(D_UU_AMIGA[4]));
    defparam D_UU_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_4_preio (
            .PADOEN(N__7467),
            .PADOUT(N__7466),
            .PADIN(N__7465),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2525),
            .DIN0(D_UU_AMIGA_in_4),
            .DOUT0(N__3377),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_7_iopad (
            .OE(N__7458),
            .DIN(N__7457),
            .DOUT(N__7456),
            .PACKAGEPIN(D_UU_040[7]));
    defparam D_UU_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_7_preio (
            .PADOEN(N__7458),
            .PADOUT(N__7457),
            .PADIN(N__7456),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5157),
            .DIN0(D_UU_040_in_7),
            .DOUT0(N__6644),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SIZ_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__7449),
            .DIN(N__7448),
            .DOUT(N__7447),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__7449),
            .PADOUT(N__7448),
            .PADIN(N__7447),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_0_iopad (
            .OE(N__7440),
            .DIN(N__7439),
            .DOUT(N__7438),
            .PACKAGEPIN(D_LL_040[0]));
    defparam D_LL_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_0_preio (
            .PADOEN(N__7440),
            .PADOUT(N__7439),
            .PADIN(N__7438),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5246),
            .DIN0(D_LL_040_in_0),
            .DOUT0(N__3458),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_2_iopad (
            .OE(N__7431),
            .DIN(N__7430),
            .DOUT(N__7429),
            .PACKAGEPIN(D_UM_AMIGA[2]));
    defparam D_UM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_2_preio (
            .PADOEN(N__7431),
            .PADOUT(N__7430),
            .PADIN(N__7429),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2633),
            .DIN0(D_UM_AMIGA_in_2),
            .DOUT0(N__3179),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_0_iopad (
            .OE(N__7422),
            .DIN(N__7421),
            .DOUT(N__7420),
            .PACKAGEPIN(D_UU_040[0]));
    defparam D_UU_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_0_preio (
            .PADOEN(N__7422),
            .PADOUT(N__7421),
            .PADIN(N__7420),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5099),
            .DIN0(D_UU_040_in_0),
            .DOUT0(N__6416),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1925 (
            .O(N__7403),
            .I(N__7400));
    LocalMux I__1924 (
            .O(N__7400),
            .I(N__7397));
    Odrv12 I__1923 (
            .O(N__7397),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ));
    InMux I__1922 (
            .O(N__7394),
            .I(N__7390));
    CascadeMux I__1921 (
            .O(N__7393),
            .I(N__7386));
    LocalMux I__1920 (
            .O(N__7390),
            .I(N__7383));
    InMux I__1919 (
            .O(N__7389),
            .I(N__7380));
    InMux I__1918 (
            .O(N__7386),
            .I(N__7377));
    Span4Mux_h I__1917 (
            .O(N__7383),
            .I(N__7374));
    LocalMux I__1916 (
            .O(N__7380),
            .I(N__7371));
    LocalMux I__1915 (
            .O(N__7377),
            .I(N__7368));
    Span4Mux_v I__1914 (
            .O(N__7374),
            .I(N__7363));
    Span4Mux_h I__1913 (
            .O(N__7371),
            .I(N__7363));
    Span4Mux_v I__1912 (
            .O(N__7368),
            .I(N__7360));
    Span4Mux_h I__1911 (
            .O(N__7363),
            .I(N__7355));
    Span4Mux_v I__1910 (
            .O(N__7360),
            .I(N__7355));
    Span4Mux_v I__1909 (
            .O(N__7355),
            .I(N__7352));
    Sp12to4 I__1908 (
            .O(N__7352),
            .I(N__7349));
    Odrv12 I__1907 (
            .O(N__7349),
            .I(D_UU_AMIGA_in_5));
    InMux I__1906 (
            .O(N__7346),
            .I(N__7340));
    InMux I__1905 (
            .O(N__7345),
            .I(N__7340));
    LocalMux I__1904 (
            .O(N__7340),
            .I(N__7335));
    InMux I__1903 (
            .O(N__7339),
            .I(N__7326));
    InMux I__1902 (
            .O(N__7338),
            .I(N__7326));
    Span4Mux_v I__1901 (
            .O(N__7335),
            .I(N__7318));
    InMux I__1900 (
            .O(N__7334),
            .I(N__7308));
    InMux I__1899 (
            .O(N__7333),
            .I(N__7308));
    InMux I__1898 (
            .O(N__7332),
            .I(N__7308));
    InMux I__1897 (
            .O(N__7331),
            .I(N__7305));
    LocalMux I__1896 (
            .O(N__7326),
            .I(N__7301));
    InMux I__1895 (
            .O(N__7325),
            .I(N__7296));
    InMux I__1894 (
            .O(N__7324),
            .I(N__7296));
    InMux I__1893 (
            .O(N__7323),
            .I(N__7293));
    InMux I__1892 (
            .O(N__7322),
            .I(N__7288));
    InMux I__1891 (
            .O(N__7321),
            .I(N__7288));
    Sp12to4 I__1890 (
            .O(N__7318),
            .I(N__7283));
    InMux I__1889 (
            .O(N__7317),
            .I(N__7280));
    InMux I__1888 (
            .O(N__7316),
            .I(N__7275));
    InMux I__1887 (
            .O(N__7315),
            .I(N__7275));
    LocalMux I__1886 (
            .O(N__7308),
            .I(N__7270));
    LocalMux I__1885 (
            .O(N__7305),
            .I(N__7270));
    InMux I__1884 (
            .O(N__7304),
            .I(N__7267));
    Span4Mux_v I__1883 (
            .O(N__7301),
            .I(N__7258));
    LocalMux I__1882 (
            .O(N__7296),
            .I(N__7258));
    LocalMux I__1881 (
            .O(N__7293),
            .I(N__7258));
    LocalMux I__1880 (
            .O(N__7288),
            .I(N__7258));
    InMux I__1879 (
            .O(N__7287),
            .I(N__7253));
    InMux I__1878 (
            .O(N__7286),
            .I(N__7253));
    Span12Mux_h I__1877 (
            .O(N__7283),
            .I(N__7248));
    LocalMux I__1876 (
            .O(N__7280),
            .I(N__7243));
    LocalMux I__1875 (
            .O(N__7275),
            .I(N__7243));
    Span4Mux_v I__1874 (
            .O(N__7270),
            .I(N__7238));
    LocalMux I__1873 (
            .O(N__7267),
            .I(N__7238));
    Span4Mux_v I__1872 (
            .O(N__7258),
            .I(N__7233));
    LocalMux I__1871 (
            .O(N__7253),
            .I(N__7233));
    InMux I__1870 (
            .O(N__7252),
            .I(N__7230));
    InMux I__1869 (
            .O(N__7251),
            .I(N__7227));
    Odrv12 I__1868 (
            .O(N__7248),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    Odrv12 I__1867 (
            .O(N__7243),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    Odrv4 I__1866 (
            .O(N__7238),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    Odrv4 I__1865 (
            .O(N__7233),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    LocalMux I__1864 (
            .O(N__7230),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    LocalMux I__1863 (
            .O(N__7227),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    IoInMux I__1862 (
            .O(N__7214),
            .I(N__7211));
    LocalMux I__1861 (
            .O(N__7211),
            .I(N__7208));
    Span4Mux_s2_v I__1860 (
            .O(N__7208),
            .I(N__7205));
    Span4Mux_v I__1859 (
            .O(N__7205),
            .I(N__7202));
    Sp12to4 I__1858 (
            .O(N__7202),
            .I(N__7199));
    Span12Mux_s10_h I__1857 (
            .O(N__7199),
            .I(N__7196));
    Odrv12 I__1856 (
            .O(N__7196),
            .I(un1_D_UU_AMIGA_5));
    CEMux I__1855 (
            .O(N__7193),
            .I(N__7185));
    CEMux I__1854 (
            .O(N__7192),
            .I(N__7182));
    CEMux I__1853 (
            .O(N__7191),
            .I(N__7179));
    CEMux I__1852 (
            .O(N__7190),
            .I(N__7176));
    CEMux I__1851 (
            .O(N__7189),
            .I(N__7173));
    CEMux I__1850 (
            .O(N__7188),
            .I(N__7170));
    LocalMux I__1849 (
            .O(N__7185),
            .I(N__7165));
    LocalMux I__1848 (
            .O(N__7182),
            .I(N__7165));
    LocalMux I__1847 (
            .O(N__7179),
            .I(N__7160));
    LocalMux I__1846 (
            .O(N__7176),
            .I(N__7160));
    LocalMux I__1845 (
            .O(N__7173),
            .I(N__7157));
    LocalMux I__1844 (
            .O(N__7170),
            .I(N__7154));
    Odrv4 I__1843 (
            .O(N__7165),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    Odrv4 I__1842 (
            .O(N__7160),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    Odrv4 I__1841 (
            .O(N__7157),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    Odrv4 I__1840 (
            .O(N__7154),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    SRMux I__1839 (
            .O(N__7145),
            .I(N__7140));
    SRMux I__1838 (
            .O(N__7144),
            .I(N__7135));
    SRMux I__1837 (
            .O(N__7143),
            .I(N__7132));
    LocalMux I__1836 (
            .O(N__7140),
            .I(N__7129));
    SRMux I__1835 (
            .O(N__7139),
            .I(N__7126));
    SRMux I__1834 (
            .O(N__7138),
            .I(N__7122));
    LocalMux I__1833 (
            .O(N__7135),
            .I(N__7119));
    LocalMux I__1832 (
            .O(N__7132),
            .I(N__7116));
    Span4Mux_h I__1831 (
            .O(N__7129),
            .I(N__7111));
    LocalMux I__1830 (
            .O(N__7126),
            .I(N__7111));
    SRMux I__1829 (
            .O(N__7125),
            .I(N__7108));
    LocalMux I__1828 (
            .O(N__7122),
            .I(N__7105));
    Span4Mux_h I__1827 (
            .O(N__7119),
            .I(N__7100));
    Span4Mux_h I__1826 (
            .O(N__7116),
            .I(N__7100));
    Span4Mux_h I__1825 (
            .O(N__7111),
            .I(N__7093));
    LocalMux I__1824 (
            .O(N__7108),
            .I(N__7093));
    Span4Mux_h I__1823 (
            .O(N__7105),
            .I(N__7093));
    Odrv4 I__1822 (
            .O(N__7100),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0 ));
    Odrv4 I__1821 (
            .O(N__7093),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0 ));
    InMux I__1820 (
            .O(N__7088),
            .I(N__7085));
    LocalMux I__1819 (
            .O(N__7085),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ));
    InMux I__1818 (
            .O(N__7082),
            .I(N__7077));
    InMux I__1817 (
            .O(N__7081),
            .I(N__7074));
    InMux I__1816 (
            .O(N__7080),
            .I(N__7071));
    LocalMux I__1815 (
            .O(N__7077),
            .I(N__7068));
    LocalMux I__1814 (
            .O(N__7074),
            .I(N__7065));
    LocalMux I__1813 (
            .O(N__7071),
            .I(N__7062));
    Span4Mux_h I__1812 (
            .O(N__7068),
            .I(N__7059));
    Span4Mux_v I__1811 (
            .O(N__7065),
            .I(N__7056));
    Span4Mux_h I__1810 (
            .O(N__7062),
            .I(N__7053));
    Sp12to4 I__1809 (
            .O(N__7059),
            .I(N__7050));
    Span4Mux_v I__1808 (
            .O(N__7056),
            .I(N__7047));
    Span4Mux_v I__1807 (
            .O(N__7053),
            .I(N__7044));
    Span12Mux_v I__1806 (
            .O(N__7050),
            .I(N__7041));
    Sp12to4 I__1805 (
            .O(N__7047),
            .I(N__7038));
    Span4Mux_h I__1804 (
            .O(N__7044),
            .I(N__7035));
    Span12Mux_v I__1803 (
            .O(N__7041),
            .I(N__7032));
    Span12Mux_h I__1802 (
            .O(N__7038),
            .I(N__7027));
    Sp12to4 I__1801 (
            .O(N__7035),
            .I(N__7027));
    Odrv12 I__1800 (
            .O(N__7032),
            .I(D_UM_AMIGA_in_3));
    Odrv12 I__1799 (
            .O(N__7027),
            .I(D_UM_AMIGA_in_3));
    IoInMux I__1798 (
            .O(N__7022),
            .I(N__7019));
    LocalMux I__1797 (
            .O(N__7019),
            .I(N__7016));
    Span4Mux_s3_h I__1796 (
            .O(N__7016),
            .I(N__7013));
    Span4Mux_h I__1795 (
            .O(N__7013),
            .I(N__7010));
    Span4Mux_h I__1794 (
            .O(N__7010),
            .I(N__7007));
    Span4Mux_h I__1793 (
            .O(N__7007),
            .I(N__7004));
    Span4Mux_v I__1792 (
            .O(N__7004),
            .I(N__7001));
    Odrv4 I__1791 (
            .O(N__7001),
            .I(un1_D_UM_AMIGA_3));
    InMux I__1790 (
            .O(N__6998),
            .I(N__6993));
    InMux I__1789 (
            .O(N__6997),
            .I(N__6990));
    InMux I__1788 (
            .O(N__6996),
            .I(N__6987));
    LocalMux I__1787 (
            .O(N__6993),
            .I(N__6984));
    LocalMux I__1786 (
            .O(N__6990),
            .I(N__6981));
    LocalMux I__1785 (
            .O(N__6987),
            .I(N__6978));
    Sp12to4 I__1784 (
            .O(N__6984),
            .I(N__6975));
    Span4Mux_v I__1783 (
            .O(N__6981),
            .I(N__6970));
    Span4Mux_v I__1782 (
            .O(N__6978),
            .I(N__6970));
    Span12Mux_v I__1781 (
            .O(N__6975),
            .I(N__6967));
    Sp12to4 I__1780 (
            .O(N__6970),
            .I(N__6964));
    Span12Mux_h I__1779 (
            .O(N__6967),
            .I(N__6961));
    Span12Mux_h I__1778 (
            .O(N__6964),
            .I(N__6958));
    Odrv12 I__1777 (
            .O(N__6961),
            .I(D_UM_AMIGA_in_1));
    Odrv12 I__1776 (
            .O(N__6958),
            .I(D_UM_AMIGA_in_1));
    InMux I__1775 (
            .O(N__6953),
            .I(N__6950));
    LocalMux I__1774 (
            .O(N__6950),
            .I(N__6947));
    Odrv4 I__1773 (
            .O(N__6947),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ));
    IoInMux I__1772 (
            .O(N__6944),
            .I(N__6941));
    LocalMux I__1771 (
            .O(N__6941),
            .I(N__6938));
    Span4Mux_s3_h I__1770 (
            .O(N__6938),
            .I(N__6935));
    Sp12to4 I__1769 (
            .O(N__6935),
            .I(N__6932));
    Span12Mux_s10_v I__1768 (
            .O(N__6932),
            .I(N__6929));
    Span12Mux_h I__1767 (
            .O(N__6929),
            .I(N__6926));
    Odrv12 I__1766 (
            .O(N__6926),
            .I(un1_D_UM_AMIGA_1));
    InMux I__1765 (
            .O(N__6923),
            .I(N__6920));
    LocalMux I__1764 (
            .O(N__6920),
            .I(N__6917));
    Odrv4 I__1763 (
            .O(N__6917),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ));
    InMux I__1762 (
            .O(N__6914),
            .I(N__6911));
    LocalMux I__1761 (
            .O(N__6911),
            .I(N__6906));
    InMux I__1760 (
            .O(N__6910),
            .I(N__6903));
    InMux I__1759 (
            .O(N__6909),
            .I(N__6900));
    Span4Mux_v I__1758 (
            .O(N__6906),
            .I(N__6895));
    LocalMux I__1757 (
            .O(N__6903),
            .I(N__6895));
    LocalMux I__1756 (
            .O(N__6900),
            .I(N__6892));
    Span4Mux_v I__1755 (
            .O(N__6895),
            .I(N__6889));
    Span12Mux_v I__1754 (
            .O(N__6892),
            .I(N__6886));
    Sp12to4 I__1753 (
            .O(N__6889),
            .I(N__6883));
    Span12Mux_h I__1752 (
            .O(N__6886),
            .I(N__6880));
    Span12Mux_h I__1751 (
            .O(N__6883),
            .I(N__6877));
    Odrv12 I__1750 (
            .O(N__6880),
            .I(D_UU_AMIGA_in_1));
    Odrv12 I__1749 (
            .O(N__6877),
            .I(D_UU_AMIGA_in_1));
    IoInMux I__1748 (
            .O(N__6872),
            .I(N__6869));
    LocalMux I__1747 (
            .O(N__6869),
            .I(N__6866));
    IoSpan4Mux I__1746 (
            .O(N__6866),
            .I(N__6863));
    IoSpan4Mux I__1745 (
            .O(N__6863),
            .I(N__6860));
    Span4Mux_s2_h I__1744 (
            .O(N__6860),
            .I(N__6857));
    Sp12to4 I__1743 (
            .O(N__6857),
            .I(N__6854));
    Odrv12 I__1742 (
            .O(N__6854),
            .I(un1_D_UU_AMIGA_1));
    InMux I__1741 (
            .O(N__6851),
            .I(N__6848));
    LocalMux I__1740 (
            .O(N__6848),
            .I(N__6845));
    Odrv4 I__1739 (
            .O(N__6845),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ));
    InMux I__1738 (
            .O(N__6842),
            .I(N__6839));
    LocalMux I__1737 (
            .O(N__6839),
            .I(N__6835));
    InMux I__1736 (
            .O(N__6838),
            .I(N__6832));
    Span4Mux_v I__1735 (
            .O(N__6835),
            .I(N__6828));
    LocalMux I__1734 (
            .O(N__6832),
            .I(N__6825));
    InMux I__1733 (
            .O(N__6831),
            .I(N__6822));
    Span4Mux_v I__1732 (
            .O(N__6828),
            .I(N__6819));
    Span4Mux_v I__1731 (
            .O(N__6825),
            .I(N__6814));
    LocalMux I__1730 (
            .O(N__6822),
            .I(N__6814));
    Sp12to4 I__1729 (
            .O(N__6819),
            .I(N__6811));
    Span4Mux_v I__1728 (
            .O(N__6814),
            .I(N__6808));
    Span12Mux_s5_h I__1727 (
            .O(N__6811),
            .I(N__6805));
    Sp12to4 I__1726 (
            .O(N__6808),
            .I(N__6802));
    Span12Mux_v I__1725 (
            .O(N__6805),
            .I(N__6797));
    Span12Mux_h I__1724 (
            .O(N__6802),
            .I(N__6797));
    Odrv12 I__1723 (
            .O(N__6797),
            .I(D_UM_AMIGA_in_4));
    IoInMux I__1722 (
            .O(N__6794),
            .I(N__6791));
    LocalMux I__1721 (
            .O(N__6791),
            .I(N__6788));
    IoSpan4Mux I__1720 (
            .O(N__6788),
            .I(N__6785));
    IoSpan4Mux I__1719 (
            .O(N__6785),
            .I(N__6782));
    Span4Mux_s3_v I__1718 (
            .O(N__6782),
            .I(N__6779));
    Span4Mux_h I__1717 (
            .O(N__6779),
            .I(N__6776));
    Span4Mux_v I__1716 (
            .O(N__6776),
            .I(N__6773));
    Odrv4 I__1715 (
            .O(N__6773),
            .I(un1_D_UM_AMIGA_4));
    InMux I__1714 (
            .O(N__6770),
            .I(N__6766));
    InMux I__1713 (
            .O(N__6769),
            .I(N__6763));
    LocalMux I__1712 (
            .O(N__6766),
            .I(N__6759));
    LocalMux I__1711 (
            .O(N__6763),
            .I(N__6756));
    InMux I__1710 (
            .O(N__6762),
            .I(N__6753));
    Span4Mux_h I__1709 (
            .O(N__6759),
            .I(N__6750));
    Span4Mux_v I__1708 (
            .O(N__6756),
            .I(N__6745));
    LocalMux I__1707 (
            .O(N__6753),
            .I(N__6745));
    Span4Mux_v I__1706 (
            .O(N__6750),
            .I(N__6742));
    Span4Mux_v I__1705 (
            .O(N__6745),
            .I(N__6739));
    Sp12to4 I__1704 (
            .O(N__6742),
            .I(N__6736));
    Sp12to4 I__1703 (
            .O(N__6739),
            .I(N__6733));
    Span12Mux_v I__1702 (
            .O(N__6736),
            .I(N__6730));
    Span12Mux_h I__1701 (
            .O(N__6733),
            .I(N__6727));
    Odrv12 I__1700 (
            .O(N__6730),
            .I(D_UM_AMIGA_in_7));
    Odrv12 I__1699 (
            .O(N__6727),
            .I(D_UM_AMIGA_in_7));
    InMux I__1698 (
            .O(N__6722),
            .I(N__6719));
    LocalMux I__1697 (
            .O(N__6719),
            .I(N__6716));
    Odrv12 I__1696 (
            .O(N__6716),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ));
    IoInMux I__1695 (
            .O(N__6713),
            .I(N__6710));
    LocalMux I__1694 (
            .O(N__6710),
            .I(N__6707));
    IoSpan4Mux I__1693 (
            .O(N__6707),
            .I(N__6704));
    Span4Mux_s1_h I__1692 (
            .O(N__6704),
            .I(N__6701));
    Sp12to4 I__1691 (
            .O(N__6701),
            .I(N__6698));
    Span12Mux_h I__1690 (
            .O(N__6698),
            .I(N__6695));
    Odrv12 I__1689 (
            .O(N__6695),
            .I(un1_D_UM_AMIGA_7));
    InMux I__1688 (
            .O(N__6692),
            .I(N__6689));
    LocalMux I__1687 (
            .O(N__6689),
            .I(N__6686));
    Odrv12 I__1686 (
            .O(N__6686),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ));
    InMux I__1685 (
            .O(N__6683),
            .I(N__6678));
    InMux I__1684 (
            .O(N__6682),
            .I(N__6675));
    InMux I__1683 (
            .O(N__6681),
            .I(N__6672));
    LocalMux I__1682 (
            .O(N__6678),
            .I(N__6669));
    LocalMux I__1681 (
            .O(N__6675),
            .I(N__6666));
    LocalMux I__1680 (
            .O(N__6672),
            .I(N__6663));
    Span4Mux_v I__1679 (
            .O(N__6669),
            .I(N__6658));
    Span4Mux_v I__1678 (
            .O(N__6666),
            .I(N__6658));
    Span4Mux_v I__1677 (
            .O(N__6663),
            .I(N__6655));
    Sp12to4 I__1676 (
            .O(N__6658),
            .I(N__6650));
    Sp12to4 I__1675 (
            .O(N__6655),
            .I(N__6650));
    Span12Mux_h I__1674 (
            .O(N__6650),
            .I(N__6647));
    Odrv12 I__1673 (
            .O(N__6647),
            .I(D_UU_AMIGA_in_7));
    IoInMux I__1672 (
            .O(N__6644),
            .I(N__6641));
    LocalMux I__1671 (
            .O(N__6641),
            .I(N__6638));
    Span12Mux_s10_v I__1670 (
            .O(N__6638),
            .I(N__6635));
    Span12Mux_h I__1669 (
            .O(N__6635),
            .I(N__6632));
    Odrv12 I__1668 (
            .O(N__6632),
            .I(un1_D_UU_AMIGA_7));
    IoInMux I__1667 (
            .O(N__6629),
            .I(N__6626));
    LocalMux I__1666 (
            .O(N__6626),
            .I(N__6623));
    Span4Mux_s2_h I__1665 (
            .O(N__6623),
            .I(N__6620));
    Span4Mux_h I__1664 (
            .O(N__6620),
            .I(N__6617));
    Span4Mux_h I__1663 (
            .O(N__6617),
            .I(N__6614));
    Span4Mux_h I__1662 (
            .O(N__6614),
            .I(N__6611));
    Odrv4 I__1661 (
            .O(N__6611),
            .I(un1_D_UM_AMIGA_0));
    IoInMux I__1660 (
            .O(N__6608),
            .I(N__6605));
    LocalMux I__1659 (
            .O(N__6605),
            .I(N__6602));
    Span4Mux_s2_h I__1658 (
            .O(N__6602),
            .I(N__6599));
    Span4Mux_h I__1657 (
            .O(N__6599),
            .I(N__6596));
    Sp12to4 I__1656 (
            .O(N__6596),
            .I(N__6593));
    Span12Mux_v I__1655 (
            .O(N__6593),
            .I(N__6590));
    Odrv12 I__1654 (
            .O(N__6590),
            .I(un1_D_UM_AMIGA_6));
    InMux I__1653 (
            .O(N__6587),
            .I(N__6583));
    InMux I__1652 (
            .O(N__6586),
            .I(N__6579));
    LocalMux I__1651 (
            .O(N__6583),
            .I(N__6576));
    InMux I__1650 (
            .O(N__6582),
            .I(N__6573));
    LocalMux I__1649 (
            .O(N__6579),
            .I(N__6570));
    Span4Mux_h I__1648 (
            .O(N__6576),
            .I(N__6567));
    LocalMux I__1647 (
            .O(N__6573),
            .I(N__6564));
    Sp12to4 I__1646 (
            .O(N__6570),
            .I(N__6561));
    Sp12to4 I__1645 (
            .O(N__6567),
            .I(N__6558));
    Span12Mux_h I__1644 (
            .O(N__6564),
            .I(N__6553));
    Span12Mux_v I__1643 (
            .O(N__6561),
            .I(N__6553));
    Span12Mux_v I__1642 (
            .O(N__6558),
            .I(N__6550));
    Span12Mux_v I__1641 (
            .O(N__6553),
            .I(N__6547));
    Span12Mux_h I__1640 (
            .O(N__6550),
            .I(N__6544));
    Odrv12 I__1639 (
            .O(N__6547),
            .I(D_UM_AMIGA_in_6));
    Odrv12 I__1638 (
            .O(N__6544),
            .I(D_UM_AMIGA_in_6));
    InMux I__1637 (
            .O(N__6539),
            .I(N__6536));
    LocalMux I__1636 (
            .O(N__6536),
            .I(N__6533));
    Odrv4 I__1635 (
            .O(N__6533),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ));
    CascadeMux I__1634 (
            .O(N__6530),
            .I(N__6527));
    InMux I__1633 (
            .O(N__6527),
            .I(N__6524));
    LocalMux I__1632 (
            .O(N__6524),
            .I(N__6521));
    Span4Mux_v I__1631 (
            .O(N__6521),
            .I(N__6517));
    InMux I__1630 (
            .O(N__6520),
            .I(N__6514));
    Span4Mux_v I__1629 (
            .O(N__6517),
            .I(N__6511));
    LocalMux I__1628 (
            .O(N__6514),
            .I(N__6508));
    Span4Mux_v I__1627 (
            .O(N__6511),
            .I(N__6502));
    Span4Mux_v I__1626 (
            .O(N__6508),
            .I(N__6502));
    InMux I__1625 (
            .O(N__6507),
            .I(N__6499));
    Sp12to4 I__1624 (
            .O(N__6502),
            .I(N__6494));
    LocalMux I__1623 (
            .O(N__6499),
            .I(N__6494));
    Span12Mux_h I__1622 (
            .O(N__6494),
            .I(N__6491));
    Odrv12 I__1621 (
            .O(N__6491),
            .I(D_UM_AMIGA_in_0));
    InMux I__1620 (
            .O(N__6488),
            .I(N__6485));
    LocalMux I__1619 (
            .O(N__6485),
            .I(N__6482));
    Odrv4 I__1618 (
            .O(N__6482),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ));
    InMux I__1617 (
            .O(N__6479),
            .I(N__6476));
    LocalMux I__1616 (
            .O(N__6476),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa ));
    InMux I__1615 (
            .O(N__6473),
            .I(N__6470));
    LocalMux I__1614 (
            .O(N__6470),
            .I(N__6467));
    Odrv4 I__1613 (
            .O(N__6467),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ));
    InMux I__1612 (
            .O(N__6464),
            .I(N__6460));
    InMux I__1611 (
            .O(N__6463),
            .I(N__6457));
    LocalMux I__1610 (
            .O(N__6460),
            .I(N__6453));
    LocalMux I__1609 (
            .O(N__6457),
            .I(N__6450));
    InMux I__1608 (
            .O(N__6456),
            .I(N__6447));
    Span4Mux_h I__1607 (
            .O(N__6453),
            .I(N__6444));
    Span4Mux_v I__1606 (
            .O(N__6450),
            .I(N__6439));
    LocalMux I__1605 (
            .O(N__6447),
            .I(N__6439));
    Span4Mux_h I__1604 (
            .O(N__6444),
            .I(N__6436));
    Span4Mux_v I__1603 (
            .O(N__6439),
            .I(N__6433));
    Sp12to4 I__1602 (
            .O(N__6436),
            .I(N__6430));
    Sp12to4 I__1601 (
            .O(N__6433),
            .I(N__6427));
    Span12Mux_v I__1600 (
            .O(N__6430),
            .I(N__6424));
    Span12Mux_h I__1599 (
            .O(N__6427),
            .I(N__6421));
    Odrv12 I__1598 (
            .O(N__6424),
            .I(D_UU_AMIGA_in_0));
    Odrv12 I__1597 (
            .O(N__6421),
            .I(D_UU_AMIGA_in_0));
    IoInMux I__1596 (
            .O(N__6416),
            .I(N__6413));
    LocalMux I__1595 (
            .O(N__6413),
            .I(N__6410));
    Span12Mux_s7_v I__1594 (
            .O(N__6410),
            .I(N__6407));
    Span12Mux_h I__1593 (
            .O(N__6407),
            .I(N__6404));
    Odrv12 I__1592 (
            .O(N__6404),
            .I(un1_D_UU_AMIGA_0));
    InMux I__1591 (
            .O(N__6401),
            .I(N__6398));
    LocalMux I__1590 (
            .O(N__6398),
            .I(N__6395));
    Odrv4 I__1589 (
            .O(N__6395),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ));
    CascadeMux I__1588 (
            .O(N__6392),
            .I(N__6389));
    InMux I__1587 (
            .O(N__6389),
            .I(N__6386));
    LocalMux I__1586 (
            .O(N__6386),
            .I(N__6381));
    InMux I__1585 (
            .O(N__6385),
            .I(N__6378));
    InMux I__1584 (
            .O(N__6384),
            .I(N__6375));
    Span4Mux_v I__1583 (
            .O(N__6381),
            .I(N__6372));
    LocalMux I__1582 (
            .O(N__6378),
            .I(N__6367));
    LocalMux I__1581 (
            .O(N__6375),
            .I(N__6367));
    Sp12to4 I__1580 (
            .O(N__6372),
            .I(N__6364));
    Span4Mux_v I__1579 (
            .O(N__6367),
            .I(N__6361));
    Span12Mux_h I__1578 (
            .O(N__6364),
            .I(N__6358));
    Sp12to4 I__1577 (
            .O(N__6361),
            .I(N__6355));
    Span12Mux_v I__1576 (
            .O(N__6358),
            .I(N__6350));
    Span12Mux_h I__1575 (
            .O(N__6355),
            .I(N__6350));
    Odrv12 I__1574 (
            .O(N__6350),
            .I(D_UM_AMIGA_in_5));
    IoInMux I__1573 (
            .O(N__6347),
            .I(N__6344));
    LocalMux I__1572 (
            .O(N__6344),
            .I(N__6341));
    Span4Mux_s1_v I__1571 (
            .O(N__6341),
            .I(N__6338));
    Sp12to4 I__1570 (
            .O(N__6338),
            .I(N__6335));
    Span12Mux_h I__1569 (
            .O(N__6335),
            .I(N__6332));
    Odrv12 I__1568 (
            .O(N__6332),
            .I(un1_D_UM_AMIGA_5));
    InMux I__1567 (
            .O(N__6329),
            .I(N__6323));
    InMux I__1566 (
            .O(N__6328),
            .I(N__6318));
    InMux I__1565 (
            .O(N__6327),
            .I(N__6311));
    InMux I__1564 (
            .O(N__6326),
            .I(N__6311));
    LocalMux I__1563 (
            .O(N__6323),
            .I(N__6308));
    InMux I__1562 (
            .O(N__6322),
            .I(N__6303));
    InMux I__1561 (
            .O(N__6321),
            .I(N__6303));
    LocalMux I__1560 (
            .O(N__6318),
            .I(N__6299));
    InMux I__1559 (
            .O(N__6317),
            .I(N__6296));
    InMux I__1558 (
            .O(N__6316),
            .I(N__6293));
    LocalMux I__1557 (
            .O(N__6311),
            .I(N__6285));
    Span4Mux_h I__1556 (
            .O(N__6308),
            .I(N__6279));
    LocalMux I__1555 (
            .O(N__6303),
            .I(N__6279));
    InMux I__1554 (
            .O(N__6302),
            .I(N__6276));
    Span4Mux_h I__1553 (
            .O(N__6299),
            .I(N__6271));
    LocalMux I__1552 (
            .O(N__6296),
            .I(N__6271));
    LocalMux I__1551 (
            .O(N__6293),
            .I(N__6262));
    InMux I__1550 (
            .O(N__6292),
            .I(N__6257));
    InMux I__1549 (
            .O(N__6291),
            .I(N__6257));
    InMux I__1548 (
            .O(N__6290),
            .I(N__6254));
    InMux I__1547 (
            .O(N__6289),
            .I(N__6251));
    CascadeMux I__1546 (
            .O(N__6288),
            .I(N__6248));
    Span4Mux_v I__1545 (
            .O(N__6285),
            .I(N__6241));
    InMux I__1544 (
            .O(N__6284),
            .I(N__6238));
    Span4Mux_h I__1543 (
            .O(N__6279),
            .I(N__6234));
    LocalMux I__1542 (
            .O(N__6276),
            .I(N__6231));
    Span4Mux_h I__1541 (
            .O(N__6271),
            .I(N__6226));
    InMux I__1540 (
            .O(N__6270),
            .I(N__6221));
    InMux I__1539 (
            .O(N__6269),
            .I(N__6221));
    InMux I__1538 (
            .O(N__6268),
            .I(N__6218));
    InMux I__1537 (
            .O(N__6267),
            .I(N__6213));
    InMux I__1536 (
            .O(N__6266),
            .I(N__6213));
    InMux I__1535 (
            .O(N__6265),
            .I(N__6210));
    Span4Mux_v I__1534 (
            .O(N__6262),
            .I(N__6207));
    LocalMux I__1533 (
            .O(N__6257),
            .I(N__6204));
    LocalMux I__1532 (
            .O(N__6254),
            .I(N__6201));
    LocalMux I__1531 (
            .O(N__6251),
            .I(N__6198));
    InMux I__1530 (
            .O(N__6248),
            .I(N__6195));
    InMux I__1529 (
            .O(N__6247),
            .I(N__6188));
    InMux I__1528 (
            .O(N__6246),
            .I(N__6188));
    InMux I__1527 (
            .O(N__6245),
            .I(N__6188));
    InMux I__1526 (
            .O(N__6244),
            .I(N__6185));
    Span4Mux_v I__1525 (
            .O(N__6241),
            .I(N__6179));
    LocalMux I__1524 (
            .O(N__6238),
            .I(N__6179));
    InMux I__1523 (
            .O(N__6237),
            .I(N__6176));
    Span4Mux_v I__1522 (
            .O(N__6234),
            .I(N__6171));
    Span4Mux_h I__1521 (
            .O(N__6231),
            .I(N__6171));
    InMux I__1520 (
            .O(N__6230),
            .I(N__6168));
    InMux I__1519 (
            .O(N__6229),
            .I(N__6165));
    Sp12to4 I__1518 (
            .O(N__6226),
            .I(N__6158));
    LocalMux I__1517 (
            .O(N__6221),
            .I(N__6158));
    LocalMux I__1516 (
            .O(N__6218),
            .I(N__6155));
    LocalMux I__1515 (
            .O(N__6213),
            .I(N__6152));
    LocalMux I__1514 (
            .O(N__6210),
            .I(N__6149));
    Span4Mux_v I__1513 (
            .O(N__6207),
            .I(N__6144));
    Span4Mux_v I__1512 (
            .O(N__6204),
            .I(N__6144));
    Span4Mux_v I__1511 (
            .O(N__6201),
            .I(N__6139));
    Span4Mux_v I__1510 (
            .O(N__6198),
            .I(N__6139));
    LocalMux I__1509 (
            .O(N__6195),
            .I(N__6134));
    LocalMux I__1508 (
            .O(N__6188),
            .I(N__6134));
    LocalMux I__1507 (
            .O(N__6185),
            .I(N__6131));
    InMux I__1506 (
            .O(N__6184),
            .I(N__6128));
    Span4Mux_h I__1505 (
            .O(N__6179),
            .I(N__6123));
    LocalMux I__1504 (
            .O(N__6176),
            .I(N__6123));
    Span4Mux_v I__1503 (
            .O(N__6171),
            .I(N__6118));
    LocalMux I__1502 (
            .O(N__6168),
            .I(N__6118));
    LocalMux I__1501 (
            .O(N__6165),
            .I(N__6115));
    InMux I__1500 (
            .O(N__6164),
            .I(N__6110));
    InMux I__1499 (
            .O(N__6163),
            .I(N__6110));
    Span12Mux_v I__1498 (
            .O(N__6158),
            .I(N__6106));
    Span12Mux_h I__1497 (
            .O(N__6155),
            .I(N__6101));
    Span12Mux_h I__1496 (
            .O(N__6152),
            .I(N__6101));
    Span4Mux_h I__1495 (
            .O(N__6149),
            .I(N__6098));
    Span4Mux_h I__1494 (
            .O(N__6144),
            .I(N__6089));
    Span4Mux_v I__1493 (
            .O(N__6139),
            .I(N__6089));
    Span4Mux_v I__1492 (
            .O(N__6134),
            .I(N__6089));
    Span4Mux_v I__1491 (
            .O(N__6131),
            .I(N__6089));
    LocalMux I__1490 (
            .O(N__6128),
            .I(N__6086));
    Span4Mux_h I__1489 (
            .O(N__6123),
            .I(N__6077));
    Span4Mux_v I__1488 (
            .O(N__6118),
            .I(N__6077));
    Span4Mux_v I__1487 (
            .O(N__6115),
            .I(N__6077));
    LocalMux I__1486 (
            .O(N__6110),
            .I(N__6077));
    InMux I__1485 (
            .O(N__6109),
            .I(N__6074));
    Odrv12 I__1484 (
            .O(N__6106),
            .I(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ));
    Odrv12 I__1483 (
            .O(N__6101),
            .I(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ));
    Odrv4 I__1482 (
            .O(N__6098),
            .I(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ));
    Odrv4 I__1481 (
            .O(N__6089),
            .I(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ));
    Odrv12 I__1480 (
            .O(N__6086),
            .I(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ));
    Odrv4 I__1479 (
            .O(N__6077),
            .I(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ));
    LocalMux I__1478 (
            .O(N__6074),
            .I(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ));
    InMux I__1477 (
            .O(N__6059),
            .I(N__6056));
    LocalMux I__1476 (
            .O(N__6056),
            .I(N__6053));
    Sp12to4 I__1475 (
            .O(N__6053),
            .I(N__6050));
    Span12Mux_v I__1474 (
            .O(N__6050),
            .I(N__6047));
    Span12Mux_h I__1473 (
            .O(N__6047),
            .I(N__6044));
    Odrv12 I__1472 (
            .O(N__6044),
            .I(D_UU_040_in_6));
    IoInMux I__1471 (
            .O(N__6041),
            .I(N__6037));
    CascadeMux I__1470 (
            .O(N__6040),
            .I(N__6034));
    LocalMux I__1469 (
            .O(N__6037),
            .I(N__6031));
    InMux I__1468 (
            .O(N__6034),
            .I(N__6028));
    Span4Mux_s2_h I__1467 (
            .O(N__6031),
            .I(N__6025));
    LocalMux I__1466 (
            .O(N__6028),
            .I(N__6022));
    Span4Mux_v I__1465 (
            .O(N__6025),
            .I(N__6019));
    Span4Mux_v I__1464 (
            .O(N__6022),
            .I(N__6016));
    Sp12to4 I__1463 (
            .O(N__6019),
            .I(N__6013));
    Span4Mux_v I__1462 (
            .O(N__6016),
            .I(N__6010));
    Span12Mux_h I__1461 (
            .O(N__6013),
            .I(N__6007));
    Sp12to4 I__1460 (
            .O(N__6010),
            .I(N__6004));
    Span12Mux_h I__1459 (
            .O(N__6007),
            .I(N__6001));
    Span12Mux_h I__1458 (
            .O(N__6004),
            .I(N__5998));
    Odrv12 I__1457 (
            .O(N__6001),
            .I(D_LM_040_in_6));
    Odrv12 I__1456 (
            .O(N__5998),
            .I(D_LM_040_in_6));
    InMux I__1455 (
            .O(N__5993),
            .I(N__5989));
    InMux I__1454 (
            .O(N__5992),
            .I(N__5986));
    LocalMux I__1453 (
            .O(N__5989),
            .I(N__5978));
    LocalMux I__1452 (
            .O(N__5986),
            .I(N__5978));
    InMux I__1451 (
            .O(N__5985),
            .I(N__5971));
    InMux I__1450 (
            .O(N__5984),
            .I(N__5971));
    InMux I__1449 (
            .O(N__5983),
            .I(N__5971));
    Span4Mux_h I__1448 (
            .O(N__5978),
            .I(N__5961));
    LocalMux I__1447 (
            .O(N__5971),
            .I(N__5961));
    InMux I__1446 (
            .O(N__5970),
            .I(N__5958));
    InMux I__1445 (
            .O(N__5969),
            .I(N__5950));
    InMux I__1444 (
            .O(N__5968),
            .I(N__5950));
    CascadeMux I__1443 (
            .O(N__5967),
            .I(N__5946));
    CascadeMux I__1442 (
            .O(N__5966),
            .I(N__5942));
    Span4Mux_v I__1441 (
            .O(N__5961),
            .I(N__5935));
    LocalMux I__1440 (
            .O(N__5958),
            .I(N__5935));
    InMux I__1439 (
            .O(N__5957),
            .I(N__5930));
    InMux I__1438 (
            .O(N__5956),
            .I(N__5930));
    InMux I__1437 (
            .O(N__5955),
            .I(N__5927));
    LocalMux I__1436 (
            .O(N__5950),
            .I(N__5923));
    InMux I__1435 (
            .O(N__5949),
            .I(N__5920));
    InMux I__1434 (
            .O(N__5946),
            .I(N__5914));
    InMux I__1433 (
            .O(N__5945),
            .I(N__5914));
    InMux I__1432 (
            .O(N__5942),
            .I(N__5909));
    CascadeMux I__1431 (
            .O(N__5941),
            .I(N__5906));
    CascadeMux I__1430 (
            .O(N__5940),
            .I(N__5903));
    Span4Mux_h I__1429 (
            .O(N__5935),
            .I(N__5898));
    LocalMux I__1428 (
            .O(N__5930),
            .I(N__5898));
    LocalMux I__1427 (
            .O(N__5927),
            .I(N__5895));
    InMux I__1426 (
            .O(N__5926),
            .I(N__5892));
    Span4Mux_h I__1425 (
            .O(N__5923),
            .I(N__5887));
    LocalMux I__1424 (
            .O(N__5920),
            .I(N__5887));
    InMux I__1423 (
            .O(N__5919),
            .I(N__5884));
    LocalMux I__1422 (
            .O(N__5914),
            .I(N__5880));
    InMux I__1421 (
            .O(N__5913),
            .I(N__5877));
    InMux I__1420 (
            .O(N__5912),
            .I(N__5874));
    LocalMux I__1419 (
            .O(N__5909),
            .I(N__5871));
    InMux I__1418 (
            .O(N__5906),
            .I(N__5868));
    InMux I__1417 (
            .O(N__5903),
            .I(N__5865));
    Span4Mux_v I__1416 (
            .O(N__5898),
            .I(N__5861));
    Span4Mux_v I__1415 (
            .O(N__5895),
            .I(N__5854));
    LocalMux I__1414 (
            .O(N__5892),
            .I(N__5854));
    Span4Mux_v I__1413 (
            .O(N__5887),
            .I(N__5846));
    LocalMux I__1412 (
            .O(N__5884),
            .I(N__5846));
    InMux I__1411 (
            .O(N__5883),
            .I(N__5843));
    Span4Mux_v I__1410 (
            .O(N__5880),
            .I(N__5840));
    LocalMux I__1409 (
            .O(N__5877),
            .I(N__5837));
    LocalMux I__1408 (
            .O(N__5874),
            .I(N__5834));
    Span4Mux_v I__1407 (
            .O(N__5871),
            .I(N__5826));
    LocalMux I__1406 (
            .O(N__5868),
            .I(N__5826));
    LocalMux I__1405 (
            .O(N__5865),
            .I(N__5826));
    InMux I__1404 (
            .O(N__5864),
            .I(N__5823));
    Span4Mux_v I__1403 (
            .O(N__5861),
            .I(N__5820));
    InMux I__1402 (
            .O(N__5860),
            .I(N__5817));
    InMux I__1401 (
            .O(N__5859),
            .I(N__5814));
    Span4Mux_v I__1400 (
            .O(N__5854),
            .I(N__5811));
    InMux I__1399 (
            .O(N__5853),
            .I(N__5806));
    InMux I__1398 (
            .O(N__5852),
            .I(N__5806));
    InMux I__1397 (
            .O(N__5851),
            .I(N__5803));
    Span4Mux_v I__1396 (
            .O(N__5846),
            .I(N__5798));
    LocalMux I__1395 (
            .O(N__5843),
            .I(N__5798));
    Span4Mux_h I__1394 (
            .O(N__5840),
            .I(N__5790));
    Span4Mux_v I__1393 (
            .O(N__5837),
            .I(N__5790));
    Span12Mux_h I__1392 (
            .O(N__5834),
            .I(N__5787));
    IoInMux I__1391 (
            .O(N__5833),
            .I(N__5784));
    Span4Mux_v I__1390 (
            .O(N__5826),
            .I(N__5779));
    LocalMux I__1389 (
            .O(N__5823),
            .I(N__5779));
    Sp12to4 I__1388 (
            .O(N__5820),
            .I(N__5770));
    LocalMux I__1387 (
            .O(N__5817),
            .I(N__5770));
    LocalMux I__1386 (
            .O(N__5814),
            .I(N__5770));
    Sp12to4 I__1385 (
            .O(N__5811),
            .I(N__5770));
    LocalMux I__1384 (
            .O(N__5806),
            .I(N__5765));
    LocalMux I__1383 (
            .O(N__5803),
            .I(N__5765));
    Span4Mux_h I__1382 (
            .O(N__5798),
            .I(N__5762));
    InMux I__1381 (
            .O(N__5797),
            .I(N__5757));
    InMux I__1380 (
            .O(N__5796),
            .I(N__5757));
    InMux I__1379 (
            .O(N__5795),
            .I(N__5754));
    Span4Mux_h I__1378 (
            .O(N__5790),
            .I(N__5751));
    Span12Mux_v I__1377 (
            .O(N__5787),
            .I(N__5746));
    LocalMux I__1376 (
            .O(N__5784),
            .I(N__5746));
    Span4Mux_h I__1375 (
            .O(N__5779),
            .I(N__5743));
    Span12Mux_h I__1374 (
            .O(N__5770),
            .I(N__5732));
    Span12Mux_v I__1373 (
            .O(N__5765),
            .I(N__5732));
    Sp12to4 I__1372 (
            .O(N__5762),
            .I(N__5732));
    LocalMux I__1371 (
            .O(N__5757),
            .I(N__5732));
    LocalMux I__1370 (
            .O(N__5754),
            .I(N__5732));
    Odrv4 I__1369 (
            .O(N__5751),
            .I(A_AMIGA_c_1));
    Odrv12 I__1368 (
            .O(N__5746),
            .I(A_AMIGA_c_1));
    Odrv4 I__1367 (
            .O(N__5743),
            .I(A_AMIGA_c_1));
    Odrv12 I__1366 (
            .O(N__5732),
            .I(A_AMIGA_c_1));
    IoInMux I__1365 (
            .O(N__5723),
            .I(N__5720));
    LocalMux I__1364 (
            .O(N__5720),
            .I(N__5717));
    Span12Mux_s10_v I__1363 (
            .O(N__5717),
            .I(N__5714));
    Span12Mux_h I__1362 (
            .O(N__5714),
            .I(N__5711));
    Odrv12 I__1361 (
            .O(N__5711),
            .I(un1_D_UU_040_6));
    CascadeMux I__1360 (
            .O(N__5708),
            .I(N__5705));
    InMux I__1359 (
            .O(N__5705),
            .I(N__5702));
    LocalMux I__1358 (
            .O(N__5702),
            .I(N__5697));
    InMux I__1357 (
            .O(N__5701),
            .I(N__5694));
    InMux I__1356 (
            .O(N__5700),
            .I(N__5691));
    Span4Mux_v I__1355 (
            .O(N__5697),
            .I(N__5686));
    LocalMux I__1354 (
            .O(N__5694),
            .I(N__5686));
    LocalMux I__1353 (
            .O(N__5691),
            .I(N__5683));
    Span4Mux_v I__1352 (
            .O(N__5686),
            .I(N__5678));
    Span4Mux_v I__1351 (
            .O(N__5683),
            .I(N__5678));
    Sp12to4 I__1350 (
            .O(N__5678),
            .I(N__5675));
    Span12Mux_h I__1349 (
            .O(N__5675),
            .I(N__5672));
    Odrv12 I__1348 (
            .O(N__5672),
            .I(D_UU_AMIGA_in_4));
    InMux I__1347 (
            .O(N__5669),
            .I(N__5666));
    LocalMux I__1346 (
            .O(N__5666),
            .I(N__5663));
    Odrv12 I__1345 (
            .O(N__5663),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ));
    IoInMux I__1344 (
            .O(N__5660),
            .I(N__5657));
    LocalMux I__1343 (
            .O(N__5657),
            .I(N__5654));
    Span4Mux_s2_v I__1342 (
            .O(N__5654),
            .I(N__5651));
    Span4Mux_h I__1341 (
            .O(N__5651),
            .I(N__5648));
    Span4Mux_h I__1340 (
            .O(N__5648),
            .I(N__5645));
    Span4Mux_v I__1339 (
            .O(N__5645),
            .I(N__5642));
    Odrv4 I__1338 (
            .O(N__5642),
            .I(un1_D_UU_AMIGA_4));
    InMux I__1337 (
            .O(N__5639),
            .I(N__5636));
    LocalMux I__1336 (
            .O(N__5636),
            .I(N__5633));
    Glb2LocalMux I__1335 (
            .O(N__5633),
            .I(N__5600));
    ClkMux I__1334 (
            .O(N__5632),
            .I(N__5600));
    ClkMux I__1333 (
            .O(N__5631),
            .I(N__5600));
    ClkMux I__1332 (
            .O(N__5630),
            .I(N__5600));
    ClkMux I__1331 (
            .O(N__5629),
            .I(N__5600));
    ClkMux I__1330 (
            .O(N__5628),
            .I(N__5600));
    ClkMux I__1329 (
            .O(N__5627),
            .I(N__5600));
    ClkMux I__1328 (
            .O(N__5626),
            .I(N__5600));
    ClkMux I__1327 (
            .O(N__5625),
            .I(N__5600));
    ClkMux I__1326 (
            .O(N__5624),
            .I(N__5600));
    ClkMux I__1325 (
            .O(N__5623),
            .I(N__5600));
    GlobalMux I__1324 (
            .O(N__5600),
            .I(CLK80));
    IoInMux I__1323 (
            .O(N__5597),
            .I(N__5594));
    LocalMux I__1322 (
            .O(N__5594),
            .I(N__5590));
    IoInMux I__1321 (
            .O(N__5593),
            .I(N__5587));
    IoSpan4Mux I__1320 (
            .O(N__5590),
            .I(N__5584));
    LocalMux I__1319 (
            .O(N__5587),
            .I(N__5580));
    IoSpan4Mux I__1318 (
            .O(N__5584),
            .I(N__5577));
    IoInMux I__1317 (
            .O(N__5583),
            .I(N__5574));
    IoSpan4Mux I__1316 (
            .O(N__5580),
            .I(N__5571));
    Sp12to4 I__1315 (
            .O(N__5577),
            .I(N__5566));
    LocalMux I__1314 (
            .O(N__5574),
            .I(N__5566));
    Span4Mux_s2_h I__1313 (
            .O(N__5571),
            .I(N__5563));
    Span12Mux_s9_v I__1312 (
            .O(N__5566),
            .I(N__5560));
    Sp12to4 I__1311 (
            .O(N__5563),
            .I(N__5557));
    Odrv12 I__1310 (
            .O(N__5560),
            .I(GB_BUFFER_CLK80_THRU_CO));
    Odrv12 I__1309 (
            .O(N__5557),
            .I(GB_BUFFER_CLK80_THRU_CO));
    InMux I__1308 (
            .O(N__5552),
            .I(N__5549));
    LocalMux I__1307 (
            .O(N__5549),
            .I(\U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0 ));
    InMux I__1306 (
            .O(N__5546),
            .I(N__5540));
    InMux I__1305 (
            .O(N__5545),
            .I(N__5537));
    InMux I__1304 (
            .O(N__5544),
            .I(N__5532));
    InMux I__1303 (
            .O(N__5543),
            .I(N__5532));
    LocalMux I__1302 (
            .O(N__5540),
            .I(N__5528));
    LocalMux I__1301 (
            .O(N__5537),
            .I(N__5525));
    LocalMux I__1300 (
            .O(N__5532),
            .I(N__5522));
    ClkMux I__1299 (
            .O(N__5531),
            .I(N__5513));
    Glb2LocalMux I__1298 (
            .O(N__5528),
            .I(N__5513));
    Glb2LocalMux I__1297 (
            .O(N__5525),
            .I(N__5513));
    Glb2LocalMux I__1296 (
            .O(N__5522),
            .I(N__5513));
    GlobalMux I__1295 (
            .O(N__5513),
            .I(CLK40));
    CascadeMux I__1294 (
            .O(N__5510),
            .I(\U111_CYCLE_SM.N_91_cascade_ ));
    InMux I__1293 (
            .O(N__5507),
            .I(N__5504));
    LocalMux I__1292 (
            .O(N__5504),
            .I(N__5497));
    InMux I__1291 (
            .O(N__5503),
            .I(N__5494));
    InMux I__1290 (
            .O(N__5502),
            .I(N__5489));
    InMux I__1289 (
            .O(N__5501),
            .I(N__5489));
    InMux I__1288 (
            .O(N__5500),
            .I(N__5486));
    Odrv4 I__1287 (
            .O(N__5497),
            .I(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ));
    LocalMux I__1286 (
            .O(N__5494),
            .I(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ));
    LocalMux I__1285 (
            .O(N__5489),
            .I(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ));
    LocalMux I__1284 (
            .O(N__5486),
            .I(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ));
    CascadeMux I__1283 (
            .O(N__5477),
            .I(\U111_CYCLE_SM.A_OUT_0_cascade_ ));
    InMux I__1282 (
            .O(N__5474),
            .I(N__5471));
    LocalMux I__1281 (
            .O(N__5471),
            .I(N__5468));
    Span4Mux_v I__1280 (
            .O(N__5468),
            .I(N__5465));
    Sp12to4 I__1279 (
            .O(N__5465),
            .I(N__5462));
    Span12Mux_h I__1278 (
            .O(N__5462),
            .I(N__5459));
    Span12Mux_v I__1277 (
            .O(N__5459),
            .I(N__5455));
    InMux I__1276 (
            .O(N__5458),
            .I(N__5452));
    Odrv12 I__1275 (
            .O(N__5455),
            .I(\U111_CYCLE_SM.A_OUTZ0 ));
    LocalMux I__1274 (
            .O(N__5452),
            .I(\U111_CYCLE_SM.A_OUTZ0 ));
    CascadeMux I__1273 (
            .O(N__5447),
            .I(N__5441));
    InMux I__1272 (
            .O(N__5446),
            .I(N__5434));
    InMux I__1271 (
            .O(N__5445),
            .I(N__5434));
    InMux I__1270 (
            .O(N__5444),
            .I(N__5434));
    InMux I__1269 (
            .O(N__5441),
            .I(N__5431));
    LocalMux I__1268 (
            .O(N__5434),
            .I(N__5426));
    LocalMux I__1267 (
            .O(N__5431),
            .I(N__5426));
    Span4Mux_v I__1266 (
            .O(N__5426),
            .I(N__5422));
    InMux I__1265 (
            .O(N__5425),
            .I(N__5419));
    Sp12to4 I__1264 (
            .O(N__5422),
            .I(N__5414));
    LocalMux I__1263 (
            .O(N__5419),
            .I(N__5414));
    Span12Mux_h I__1262 (
            .O(N__5414),
            .I(N__5411));
    Span12Mux_v I__1261 (
            .O(N__5411),
            .I(N__5408));
    Odrv12 I__1260 (
            .O(N__5408),
            .I(TACKn_c));
    InMux I__1259 (
            .O(N__5405),
            .I(N__5402));
    LocalMux I__1258 (
            .O(N__5402),
            .I(N__5391));
    InMux I__1257 (
            .O(N__5401),
            .I(N__5386));
    InMux I__1256 (
            .O(N__5400),
            .I(N__5386));
    InMux I__1255 (
            .O(N__5399),
            .I(N__5381));
    InMux I__1254 (
            .O(N__5398),
            .I(N__5381));
    InMux I__1253 (
            .O(N__5397),
            .I(N__5372));
    InMux I__1252 (
            .O(N__5396),
            .I(N__5372));
    InMux I__1251 (
            .O(N__5395),
            .I(N__5372));
    InMux I__1250 (
            .O(N__5394),
            .I(N__5372));
    Odrv4 I__1249 (
            .O(N__5391),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1248 (
            .O(N__5386),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1247 (
            .O(N__5381),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1246 (
            .O(N__5372),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    InMux I__1245 (
            .O(N__5363),
            .I(N__5358));
    CascadeMux I__1244 (
            .O(N__5362),
            .I(N__5351));
    CascadeMux I__1243 (
            .O(N__5361),
            .I(N__5347));
    LocalMux I__1242 (
            .O(N__5358),
            .I(N__5343));
    InMux I__1241 (
            .O(N__5357),
            .I(N__5338));
    InMux I__1240 (
            .O(N__5356),
            .I(N__5338));
    InMux I__1239 (
            .O(N__5355),
            .I(N__5333));
    InMux I__1238 (
            .O(N__5354),
            .I(N__5333));
    InMux I__1237 (
            .O(N__5351),
            .I(N__5324));
    InMux I__1236 (
            .O(N__5350),
            .I(N__5324));
    InMux I__1235 (
            .O(N__5347),
            .I(N__5324));
    InMux I__1234 (
            .O(N__5346),
            .I(N__5324));
    Odrv4 I__1233 (
            .O(N__5343),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1232 (
            .O(N__5338),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1231 (
            .O(N__5333),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1230 (
            .O(N__5324),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    CascadeMux I__1229 (
            .O(N__5315),
            .I(N__5306));
    InMux I__1228 (
            .O(N__5314),
            .I(N__5303));
    InMux I__1227 (
            .O(N__5313),
            .I(N__5296));
    InMux I__1226 (
            .O(N__5312),
            .I(N__5296));
    InMux I__1225 (
            .O(N__5311),
            .I(N__5296));
    InMux I__1224 (
            .O(N__5310),
            .I(N__5291));
    InMux I__1223 (
            .O(N__5309),
            .I(N__5291));
    InMux I__1222 (
            .O(N__5306),
            .I(N__5288));
    LocalMux I__1221 (
            .O(N__5303),
            .I(N__5278));
    LocalMux I__1220 (
            .O(N__5296),
            .I(N__5278));
    LocalMux I__1219 (
            .O(N__5291),
            .I(N__5278));
    LocalMux I__1218 (
            .O(N__5288),
            .I(N__5278));
    InMux I__1217 (
            .O(N__5287),
            .I(N__5275));
    Span4Mux_v I__1216 (
            .O(N__5278),
            .I(N__5270));
    LocalMux I__1215 (
            .O(N__5275),
            .I(N__5270));
    Span4Mux_h I__1214 (
            .O(N__5270),
            .I(N__5267));
    Span4Mux_v I__1213 (
            .O(N__5267),
            .I(N__5263));
    InMux I__1212 (
            .O(N__5266),
            .I(N__5260));
    Sp12to4 I__1211 (
            .O(N__5263),
            .I(N__5255));
    LocalMux I__1210 (
            .O(N__5260),
            .I(N__5255));
    Span12Mux_v I__1209 (
            .O(N__5255),
            .I(N__5252));
    Odrv12 I__1208 (
            .O(N__5252),
            .I(RESETn_c));
    CascadeMux I__1207 (
            .O(N__5249),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_ ));
    IoInMux I__1206 (
            .O(N__5246),
            .I(N__5242));
    IoInMux I__1205 (
            .O(N__5245),
            .I(N__5239));
    LocalMux I__1204 (
            .O(N__5242),
            .I(N__5231));
    LocalMux I__1203 (
            .O(N__5239),
            .I(N__5231));
    IoInMux I__1202 (
            .O(N__5238),
            .I(N__5228));
    IoInMux I__1201 (
            .O(N__5237),
            .I(N__5225));
    IoInMux I__1200 (
            .O(N__5236),
            .I(N__5217));
    IoSpan4Mux I__1199 (
            .O(N__5231),
            .I(N__5210));
    LocalMux I__1198 (
            .O(N__5228),
            .I(N__5210));
    LocalMux I__1197 (
            .O(N__5225),
            .I(N__5210));
    IoInMux I__1196 (
            .O(N__5224),
            .I(N__5207));
    IoInMux I__1195 (
            .O(N__5223),
            .I(N__5204));
    IoInMux I__1194 (
            .O(N__5222),
            .I(N__5201));
    IoInMux I__1193 (
            .O(N__5221),
            .I(N__5198));
    IoInMux I__1192 (
            .O(N__5220),
            .I(N__5195));
    LocalMux I__1191 (
            .O(N__5217),
            .I(N__5190));
    IoSpan4Mux I__1190 (
            .O(N__5210),
            .I(N__5175));
    LocalMux I__1189 (
            .O(N__5207),
            .I(N__5175));
    LocalMux I__1188 (
            .O(N__5204),
            .I(N__5175));
    LocalMux I__1187 (
            .O(N__5201),
            .I(N__5175));
    LocalMux I__1186 (
            .O(N__5198),
            .I(N__5175));
    LocalMux I__1185 (
            .O(N__5195),
            .I(N__5175));
    IoInMux I__1184 (
            .O(N__5194),
            .I(N__5172));
    IoInMux I__1183 (
            .O(N__5193),
            .I(N__5169));
    Span4Mux_s3_v I__1182 (
            .O(N__5190),
            .I(N__5166));
    IoInMux I__1181 (
            .O(N__5189),
            .I(N__5162));
    IoInMux I__1180 (
            .O(N__5188),
            .I(N__5159));
    IoSpan4Mux I__1179 (
            .O(N__5175),
            .I(N__5146));
    LocalMux I__1178 (
            .O(N__5172),
            .I(N__5146));
    LocalMux I__1177 (
            .O(N__5169),
            .I(N__5146));
    Span4Mux_h I__1176 (
            .O(N__5166),
            .I(N__5142));
    InMux I__1175 (
            .O(N__5165),
            .I(N__5139));
    LocalMux I__1174 (
            .O(N__5162),
            .I(N__5134));
    LocalMux I__1173 (
            .O(N__5159),
            .I(N__5134));
    IoInMux I__1172 (
            .O(N__5158),
            .I(N__5131));
    IoInMux I__1171 (
            .O(N__5157),
            .I(N__5128));
    IoInMux I__1170 (
            .O(N__5156),
            .I(N__5125));
    IoInMux I__1169 (
            .O(N__5155),
            .I(N__5122));
    IoInMux I__1168 (
            .O(N__5154),
            .I(N__5119));
    IoInMux I__1167 (
            .O(N__5153),
            .I(N__5116));
    IoSpan4Mux I__1166 (
            .O(N__5146),
            .I(N__5109));
    IoInMux I__1165 (
            .O(N__5145),
            .I(N__5106));
    Span4Mux_v I__1164 (
            .O(N__5142),
            .I(N__5100));
    LocalMux I__1163 (
            .O(N__5139),
            .I(N__5100));
    IoSpan4Mux I__1162 (
            .O(N__5134),
            .I(N__5083));
    LocalMux I__1161 (
            .O(N__5131),
            .I(N__5083));
    LocalMux I__1160 (
            .O(N__5128),
            .I(N__5083));
    LocalMux I__1159 (
            .O(N__5125),
            .I(N__5083));
    LocalMux I__1158 (
            .O(N__5122),
            .I(N__5083));
    LocalMux I__1157 (
            .O(N__5119),
            .I(N__5083));
    LocalMux I__1156 (
            .O(N__5116),
            .I(N__5083));
    IoInMux I__1155 (
            .O(N__5115),
            .I(N__5080));
    IoInMux I__1154 (
            .O(N__5114),
            .I(N__5077));
    IoInMux I__1153 (
            .O(N__5113),
            .I(N__5074));
    IoInMux I__1152 (
            .O(N__5112),
            .I(N__5071));
    IoSpan4Mux I__1151 (
            .O(N__5109),
            .I(N__5066));
    LocalMux I__1150 (
            .O(N__5106),
            .I(N__5066));
    IoInMux I__1149 (
            .O(N__5105),
            .I(N__5063));
    Span4Mux_v I__1148 (
            .O(N__5100),
            .I(N__5057));
    IoInMux I__1147 (
            .O(N__5099),
            .I(N__5054));
    InMux I__1146 (
            .O(N__5098),
            .I(N__5051));
    IoSpan4Mux I__1145 (
            .O(N__5083),
            .I(N__5040));
    LocalMux I__1144 (
            .O(N__5080),
            .I(N__5040));
    LocalMux I__1143 (
            .O(N__5077),
            .I(N__5040));
    LocalMux I__1142 (
            .O(N__5074),
            .I(N__5040));
    LocalMux I__1141 (
            .O(N__5071),
            .I(N__5040));
    IoSpan4Mux I__1140 (
            .O(N__5066),
            .I(N__5036));
    LocalMux I__1139 (
            .O(N__5063),
            .I(N__5033));
    IoInMux I__1138 (
            .O(N__5062),
            .I(N__5030));
    IoInMux I__1137 (
            .O(N__5061),
            .I(N__5027));
    IoInMux I__1136 (
            .O(N__5060),
            .I(N__5024));
    Sp12to4 I__1135 (
            .O(N__5057),
            .I(N__5019));
    LocalMux I__1134 (
            .O(N__5054),
            .I(N__5016));
    LocalMux I__1133 (
            .O(N__5051),
            .I(N__5013));
    IoSpan4Mux I__1132 (
            .O(N__5040),
            .I(N__5010));
    IoInMux I__1131 (
            .O(N__5039),
            .I(N__5007));
    IoSpan4Mux I__1130 (
            .O(N__5036),
            .I(N__4996));
    IoSpan4Mux I__1129 (
            .O(N__5033),
            .I(N__4996));
    LocalMux I__1128 (
            .O(N__5030),
            .I(N__4996));
    LocalMux I__1127 (
            .O(N__5027),
            .I(N__4996));
    LocalMux I__1126 (
            .O(N__5024),
            .I(N__4996));
    IoInMux I__1125 (
            .O(N__5023),
            .I(N__4993));
    IoInMux I__1124 (
            .O(N__5022),
            .I(N__4990));
    Span12Mux_h I__1123 (
            .O(N__5019),
            .I(N__4987));
    Span12Mux_s11_v I__1122 (
            .O(N__5016),
            .I(N__4982));
    Span12Mux_h I__1121 (
            .O(N__5013),
            .I(N__4982));
    IoSpan4Mux I__1120 (
            .O(N__5010),
            .I(N__4977));
    LocalMux I__1119 (
            .O(N__5007),
            .I(N__4977));
    IoSpan4Mux I__1118 (
            .O(N__4996),
            .I(N__4972));
    LocalMux I__1117 (
            .O(N__4993),
            .I(N__4972));
    LocalMux I__1116 (
            .O(N__4990),
            .I(N__4969));
    Odrv12 I__1115 (
            .O(N__4987),
            .I(RnW_c));
    Odrv12 I__1114 (
            .O(N__4982),
            .I(RnW_c));
    Odrv4 I__1113 (
            .O(N__4977),
            .I(RnW_c));
    Odrv4 I__1112 (
            .O(N__4972),
            .I(RnW_c));
    Odrv12 I__1111 (
            .O(N__4969),
            .I(RnW_c));
    CascadeMux I__1110 (
            .O(N__4958),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_ ));
    InMux I__1109 (
            .O(N__4955),
            .I(N__4952));
    LocalMux I__1108 (
            .O(N__4952),
            .I(N__4949));
    Odrv4 I__1107 (
            .O(N__4949),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ));
    InMux I__1106 (
            .O(N__4946),
            .I(N__4941));
    InMux I__1105 (
            .O(N__4945),
            .I(N__4938));
    InMux I__1104 (
            .O(N__4944),
            .I(N__4935));
    LocalMux I__1103 (
            .O(N__4941),
            .I(N__4930));
    LocalMux I__1102 (
            .O(N__4938),
            .I(N__4930));
    LocalMux I__1101 (
            .O(N__4935),
            .I(N__4927));
    Span4Mux_v I__1100 (
            .O(N__4930),
            .I(N__4924));
    Sp12to4 I__1099 (
            .O(N__4927),
            .I(N__4921));
    Sp12to4 I__1098 (
            .O(N__4924),
            .I(N__4918));
    Span12Mux_v I__1097 (
            .O(N__4921),
            .I(N__4915));
    Span12Mux_h I__1096 (
            .O(N__4918),
            .I(N__4912));
    Span12Mux_h I__1095 (
            .O(N__4915),
            .I(N__4909));
    Odrv12 I__1094 (
            .O(N__4912),
            .I(D_UU_AMIGA_in_6));
    Odrv12 I__1093 (
            .O(N__4909),
            .I(D_UU_AMIGA_in_6));
    IoInMux I__1092 (
            .O(N__4904),
            .I(N__4901));
    LocalMux I__1091 (
            .O(N__4901),
            .I(N__4898));
    Span4Mux_s1_v I__1090 (
            .O(N__4898),
            .I(N__4895));
    Span4Mux_v I__1089 (
            .O(N__4895),
            .I(N__4892));
    Sp12to4 I__1088 (
            .O(N__4892),
            .I(N__4889));
    Span12Mux_h I__1087 (
            .O(N__4889),
            .I(N__4886));
    Odrv12 I__1086 (
            .O(N__4886),
            .I(un1_D_UU_AMIGA_6));
    InMux I__1085 (
            .O(N__4883),
            .I(N__4880));
    LocalMux I__1084 (
            .O(N__4880),
            .I(N__4877));
    Odrv12 I__1083 (
            .O(N__4877),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ));
    CascadeMux I__1082 (
            .O(N__4874),
            .I(N__4871));
    InMux I__1081 (
            .O(N__4871),
            .I(N__4868));
    LocalMux I__1080 (
            .O(N__4868),
            .I(N__4863));
    InMux I__1079 (
            .O(N__4867),
            .I(N__4860));
    InMux I__1078 (
            .O(N__4866),
            .I(N__4857));
    Span4Mux_v I__1077 (
            .O(N__4863),
            .I(N__4850));
    LocalMux I__1076 (
            .O(N__4860),
            .I(N__4850));
    LocalMux I__1075 (
            .O(N__4857),
            .I(N__4850));
    Span4Mux_v I__1074 (
            .O(N__4850),
            .I(N__4847));
    Sp12to4 I__1073 (
            .O(N__4847),
            .I(N__4844));
    Span12Mux_h I__1072 (
            .O(N__4844),
            .I(N__4841));
    Odrv12 I__1071 (
            .O(N__4841),
            .I(D_UU_AMIGA_in_2));
    IoInMux I__1070 (
            .O(N__4838),
            .I(N__4835));
    LocalMux I__1069 (
            .O(N__4835),
            .I(N__4832));
    Span12Mux_s1_v I__1068 (
            .O(N__4832),
            .I(N__4829));
    Span12Mux_h I__1067 (
            .O(N__4829),
            .I(N__4826));
    Odrv12 I__1066 (
            .O(N__4826),
            .I(un1_D_UU_AMIGA_2));
    IoInMux I__1065 (
            .O(N__4823),
            .I(N__4818));
    IoInMux I__1064 (
            .O(N__4822),
            .I(N__4815));
    IoInMux I__1063 (
            .O(N__4821),
            .I(N__4812));
    LocalMux I__1062 (
            .O(N__4818),
            .I(N__4809));
    LocalMux I__1061 (
            .O(N__4815),
            .I(N__4806));
    LocalMux I__1060 (
            .O(N__4812),
            .I(N__4803));
    Span12Mux_s5_v I__1059 (
            .O(N__4809),
            .I(N__4800));
    Span12Mux_s10_h I__1058 (
            .O(N__4806),
            .I(N__4795));
    Span12Mux_s9_h I__1057 (
            .O(N__4803),
            .I(N__4795));
    Odrv12 I__1056 (
            .O(N__4800),
            .I(GB_BUFFER_CLK40_THRU_CO));
    Odrv12 I__1055 (
            .O(N__4795),
            .I(GB_BUFFER_CLK40_THRU_CO));
    CascadeMux I__1054 (
            .O(N__4790),
            .I(N__4787));
    InMux I__1053 (
            .O(N__4787),
            .I(N__4784));
    LocalMux I__1052 (
            .O(N__4784),
            .I(N__4781));
    Span12Mux_h I__1051 (
            .O(N__4781),
            .I(N__4778));
    Odrv12 I__1050 (
            .O(N__4778),
            .I(D_LM_AMIGA_in_1));
    IoInMux I__1049 (
            .O(N__4775),
            .I(N__4772));
    LocalMux I__1048 (
            .O(N__4772),
            .I(N__4769));
    IoSpan4Mux I__1047 (
            .O(N__4769),
            .I(N__4766));
    Span4Mux_s2_h I__1046 (
            .O(N__4766),
            .I(N__4763));
    Sp12to4 I__1045 (
            .O(N__4763),
            .I(N__4760));
    Span12Mux_h I__1044 (
            .O(N__4760),
            .I(N__4757));
    Odrv12 I__1043 (
            .O(N__4757),
            .I(un1_D_LM_AMIGA_1));
    InMux I__1042 (
            .O(N__4754),
            .I(N__4751));
    LocalMux I__1041 (
            .O(N__4751),
            .I(N__4748));
    Span4Mux_v I__1040 (
            .O(N__4748),
            .I(N__4745));
    Sp12to4 I__1039 (
            .O(N__4745),
            .I(N__4742));
    Span12Mux_h I__1038 (
            .O(N__4742),
            .I(N__4739));
    Odrv12 I__1037 (
            .O(N__4739),
            .I(D_UM_040_in_6));
    IoInMux I__1036 (
            .O(N__4736),
            .I(N__4733));
    LocalMux I__1035 (
            .O(N__4733),
            .I(N__4729));
    CascadeMux I__1034 (
            .O(N__4732),
            .I(N__4726));
    IoSpan4Mux I__1033 (
            .O(N__4729),
            .I(N__4723));
    InMux I__1032 (
            .O(N__4726),
            .I(N__4720));
    IoSpan4Mux I__1031 (
            .O(N__4723),
            .I(N__4717));
    LocalMux I__1030 (
            .O(N__4720),
            .I(N__4714));
    Span4Mux_s2_h I__1029 (
            .O(N__4717),
            .I(N__4711));
    Span4Mux_v I__1028 (
            .O(N__4714),
            .I(N__4708));
    Sp12to4 I__1027 (
            .O(N__4711),
            .I(N__4705));
    Sp12to4 I__1026 (
            .O(N__4708),
            .I(N__4702));
    Span12Mux_h I__1025 (
            .O(N__4705),
            .I(N__4699));
    Span12Mux_h I__1024 (
            .O(N__4702),
            .I(N__4696));
    Span12Mux_h I__1023 (
            .O(N__4699),
            .I(N__4693));
    Span12Mux_v I__1022 (
            .O(N__4696),
            .I(N__4690));
    Odrv12 I__1021 (
            .O(N__4693),
            .I(D_LL_040_in_6));
    Odrv12 I__1020 (
            .O(N__4690),
            .I(D_LL_040_in_6));
    IoInMux I__1019 (
            .O(N__4685),
            .I(N__4682));
    LocalMux I__1018 (
            .O(N__4682),
            .I(N__4679));
    Span12Mux_s2_h I__1017 (
            .O(N__4679),
            .I(N__4676));
    Span12Mux_v I__1016 (
            .O(N__4676),
            .I(N__4673));
    Span12Mux_h I__1015 (
            .O(N__4673),
            .I(N__4670));
    Odrv12 I__1014 (
            .O(N__4670),
            .I(un1_D_UM_040_6));
    CascadeMux I__1013 (
            .O(N__4667),
            .I(N__4663));
    InMux I__1012 (
            .O(N__4666),
            .I(N__4660));
    InMux I__1011 (
            .O(N__4663),
            .I(N__4657));
    LocalMux I__1010 (
            .O(N__4660),
            .I(\U111_CYCLE_SM.TA_ENZ0 ));
    LocalMux I__1009 (
            .O(N__4657),
            .I(\U111_CYCLE_SM.TA_ENZ0 ));
    IoInMux I__1008 (
            .O(N__4652),
            .I(N__4649));
    LocalMux I__1007 (
            .O(N__4649),
            .I(N__4646));
    Span4Mux_s1_v I__1006 (
            .O(N__4646),
            .I(N__4643));
    Span4Mux_v I__1005 (
            .O(N__4643),
            .I(N__4640));
    Span4Mux_v I__1004 (
            .O(N__4640),
            .I(N__4637));
    Span4Mux_v I__1003 (
            .O(N__4637),
            .I(N__4634));
    Odrv4 I__1002 (
            .O(N__4634),
            .I(U111_CYCLE_SM_TAn_0_i));
    InMux I__1001 (
            .O(N__4631),
            .I(N__4628));
    LocalMux I__1000 (
            .O(N__4628),
            .I(N__4625));
    Span4Mux_v I__999 (
            .O(N__4625),
            .I(N__4622));
    Sp12to4 I__998 (
            .O(N__4622),
            .I(N__4619));
    Span12Mux_h I__997 (
            .O(N__4619),
            .I(N__4616));
    Odrv12 I__996 (
            .O(N__4616),
            .I(D_LM_AMIGA_in_4));
    IoInMux I__995 (
            .O(N__4613),
            .I(N__4610));
    LocalMux I__994 (
            .O(N__4610),
            .I(N__4607));
    IoSpan4Mux I__993 (
            .O(N__4607),
            .I(N__4604));
    Span4Mux_s2_h I__992 (
            .O(N__4604),
            .I(N__4601));
    Sp12to4 I__991 (
            .O(N__4601),
            .I(N__4598));
    Span12Mux_h I__990 (
            .O(N__4598),
            .I(N__4595));
    Odrv12 I__989 (
            .O(N__4595),
            .I(un1_D_LM_AMIGA_4));
    InMux I__988 (
            .O(N__4592),
            .I(N__4589));
    LocalMux I__987 (
            .O(N__4589),
            .I(\U111_CYCLE_SM.LW_CYCLE_0 ));
    CascadeMux I__986 (
            .O(N__4586),
            .I(\U111_CYCLE_SM.N_69_0_cascade_ ));
    InMux I__985 (
            .O(N__4583),
            .I(N__4580));
    LocalMux I__984 (
            .O(N__4580),
            .I(\U111_CYCLE_SM.TS_EN_5 ));
    InMux I__983 (
            .O(N__4577),
            .I(N__4574));
    LocalMux I__982 (
            .O(N__4574),
            .I(N__4570));
    CascadeMux I__981 (
            .O(N__4573),
            .I(N__4566));
    Span12Mux_s8_v I__980 (
            .O(N__4570),
            .I(N__4563));
    InMux I__979 (
            .O(N__4569),
            .I(N__4558));
    InMux I__978 (
            .O(N__4566),
            .I(N__4558));
    Span12Mux_v I__977 (
            .O(N__4563),
            .I(N__4555));
    LocalMux I__976 (
            .O(N__4558),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    Odrv12 I__975 (
            .O(N__4555),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    InMux I__974 (
            .O(N__4550),
            .I(N__4547));
    LocalMux I__973 (
            .O(N__4547),
            .I(N__4544));
    Span4Mux_v I__972 (
            .O(N__4544),
            .I(N__4540));
    InMux I__971 (
            .O(N__4543),
            .I(N__4537));
    Sp12to4 I__970 (
            .O(N__4540),
            .I(N__4532));
    LocalMux I__969 (
            .O(N__4537),
            .I(N__4532));
    Span12Mux_h I__968 (
            .O(N__4532),
            .I(N__4529));
    Span12Mux_v I__967 (
            .O(N__4529),
            .I(N__4526));
    Odrv12 I__966 (
            .O(N__4526),
            .I(PORTSIZE_c));
    InMux I__965 (
            .O(N__4523),
            .I(N__4520));
    LocalMux I__964 (
            .O(N__4520),
            .I(N__4516));
    InMux I__963 (
            .O(N__4519),
            .I(N__4513));
    Span4Mux_h I__962 (
            .O(N__4516),
            .I(N__4508));
    LocalMux I__961 (
            .O(N__4513),
            .I(N__4508));
    Span4Mux_v I__960 (
            .O(N__4508),
            .I(N__4505));
    Sp12to4 I__959 (
            .O(N__4505),
            .I(N__4502));
    Span12Mux_h I__958 (
            .O(N__4502),
            .I(N__4499));
    Odrv12 I__957 (
            .O(N__4499),
            .I(SIZ_c_1));
    InMux I__956 (
            .O(N__4496),
            .I(N__4492));
    CascadeMux I__955 (
            .O(N__4495),
            .I(N__4489));
    LocalMux I__954 (
            .O(N__4492),
            .I(N__4486));
    InMux I__953 (
            .O(N__4489),
            .I(N__4483));
    Span4Mux_h I__952 (
            .O(N__4486),
            .I(N__4478));
    LocalMux I__951 (
            .O(N__4483),
            .I(N__4478));
    Span4Mux_v I__950 (
            .O(N__4478),
            .I(N__4475));
    Sp12to4 I__949 (
            .O(N__4475),
            .I(N__4472));
    Span12Mux_h I__948 (
            .O(N__4472),
            .I(N__4469));
    Odrv12 I__947 (
            .O(N__4469),
            .I(SIZ_c_0));
    IoInMux I__946 (
            .O(N__4466),
            .I(N__4462));
    IoInMux I__945 (
            .O(N__4465),
            .I(N__4459));
    LocalMux I__944 (
            .O(N__4462),
            .I(N__4455));
    LocalMux I__943 (
            .O(N__4459),
            .I(N__4452));
    IoInMux I__942 (
            .O(N__4458),
            .I(N__4449));
    Span4Mux_s2_h I__941 (
            .O(N__4455),
            .I(N__4446));
    IoSpan4Mux I__940 (
            .O(N__4452),
            .I(N__4443));
    LocalMux I__939 (
            .O(N__4449),
            .I(N__4440));
    Span4Mux_h I__938 (
            .O(N__4446),
            .I(N__4437));
    IoSpan4Mux I__937 (
            .O(N__4443),
            .I(N__4434));
    Span4Mux_s2_v I__936 (
            .O(N__4440),
            .I(N__4431));
    Span4Mux_v I__935 (
            .O(N__4437),
            .I(N__4428));
    Span4Mux_s2_v I__934 (
            .O(N__4434),
            .I(N__4423));
    Span4Mux_h I__933 (
            .O(N__4431),
            .I(N__4423));
    Sp12to4 I__932 (
            .O(N__4428),
            .I(N__4420));
    Span4Mux_v I__931 (
            .O(N__4423),
            .I(N__4417));
    Odrv12 I__930 (
            .O(N__4420),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__929 (
            .O(N__4417),
            .I(CONSTANT_ONE_NET));
    InMux I__928 (
            .O(N__4412),
            .I(N__4409));
    LocalMux I__927 (
            .O(N__4409),
            .I(N__4406));
    Odrv4 I__926 (
            .O(N__4406),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ));
    CascadeMux I__925 (
            .O(N__4403),
            .I(N__4400));
    InMux I__924 (
            .O(N__4400),
            .I(N__4397));
    LocalMux I__923 (
            .O(N__4397),
            .I(N__4394));
    Span4Mux_v I__922 (
            .O(N__4394),
            .I(N__4389));
    InMux I__921 (
            .O(N__4393),
            .I(N__4386));
    InMux I__920 (
            .O(N__4392),
            .I(N__4383));
    Sp12to4 I__919 (
            .O(N__4389),
            .I(N__4380));
    LocalMux I__918 (
            .O(N__4386),
            .I(N__4375));
    LocalMux I__917 (
            .O(N__4383),
            .I(N__4375));
    Span12Mux_h I__916 (
            .O(N__4380),
            .I(N__4372));
    Span12Mux_v I__915 (
            .O(N__4375),
            .I(N__4369));
    Span12Mux_v I__914 (
            .O(N__4372),
            .I(N__4364));
    Span12Mux_h I__913 (
            .O(N__4369),
            .I(N__4364));
    Odrv12 I__912 (
            .O(N__4364),
            .I(D_UU_AMIGA_in_3));
    IoInMux I__911 (
            .O(N__4361),
            .I(N__4358));
    LocalMux I__910 (
            .O(N__4358),
            .I(N__4355));
    Span4Mux_s3_v I__909 (
            .O(N__4355),
            .I(N__4352));
    Span4Mux_h I__908 (
            .O(N__4352),
            .I(N__4349));
    Span4Mux_v I__907 (
            .O(N__4349),
            .I(N__4346));
    Sp12to4 I__906 (
            .O(N__4346),
            .I(N__4343));
    Span12Mux_h I__905 (
            .O(N__4343),
            .I(N__4340));
    Odrv12 I__904 (
            .O(N__4340),
            .I(un1_D_UU_AMIGA_3));
    InMux I__903 (
            .O(N__4337),
            .I(N__4334));
    LocalMux I__902 (
            .O(N__4334),
            .I(N__4331));
    Span4Mux_v I__901 (
            .O(N__4331),
            .I(N__4328));
    Sp12to4 I__900 (
            .O(N__4328),
            .I(N__4325));
    Span12Mux_h I__899 (
            .O(N__4325),
            .I(N__4322));
    Odrv12 I__898 (
            .O(N__4322),
            .I(D_LL_AMIGA_in_5));
    IoInMux I__897 (
            .O(N__4319),
            .I(N__4316));
    LocalMux I__896 (
            .O(N__4316),
            .I(N__4313));
    Span4Mux_s2_h I__895 (
            .O(N__4313),
            .I(N__4310));
    Span4Mux_v I__894 (
            .O(N__4310),
            .I(N__4307));
    Span4Mux_v I__893 (
            .O(N__4307),
            .I(N__4304));
    Sp12to4 I__892 (
            .O(N__4304),
            .I(N__4301));
    Span12Mux_s9_h I__891 (
            .O(N__4301),
            .I(N__4298));
    Odrv12 I__890 (
            .O(N__4298),
            .I(un1_D_LL_AMIGA_5));
    InMux I__889 (
            .O(N__4295),
            .I(N__4292));
    LocalMux I__888 (
            .O(N__4292),
            .I(N__4289));
    Span12Mux_h I__887 (
            .O(N__4289),
            .I(N__4286));
    Odrv12 I__886 (
            .O(N__4286),
            .I(D_LL_AMIGA_in_7));
    IoInMux I__885 (
            .O(N__4283),
            .I(N__4280));
    LocalMux I__884 (
            .O(N__4280),
            .I(N__4277));
    Span4Mux_s3_h I__883 (
            .O(N__4277),
            .I(N__4274));
    Span4Mux_v I__882 (
            .O(N__4274),
            .I(N__4271));
    Sp12to4 I__881 (
            .O(N__4271),
            .I(N__4268));
    Span12Mux_h I__880 (
            .O(N__4268),
            .I(N__4265));
    Odrv12 I__879 (
            .O(N__4265),
            .I(un1_D_LL_AMIGA_7));
    IoInMux I__878 (
            .O(N__4262),
            .I(N__4259));
    LocalMux I__877 (
            .O(N__4259),
            .I(N__4256));
    Span12Mux_s5_h I__876 (
            .O(N__4256),
            .I(N__4253));
    Span12Mux_h I__875 (
            .O(N__4253),
            .I(N__4250));
    Odrv12 I__874 (
            .O(N__4250),
            .I(un1_D_UM_AMIGA_2));
    SRMux I__873 (
            .O(N__4247),
            .I(N__4244));
    LocalMux I__872 (
            .O(N__4244),
            .I(N__4241));
    Odrv4 I__871 (
            .O(N__4241),
            .I(\U111_CYCLE_SM.RESETn_c_i ));
    InMux I__870 (
            .O(N__4238),
            .I(N__4234));
    InMux I__869 (
            .O(N__4237),
            .I(N__4231));
    LocalMux I__868 (
            .O(N__4234),
            .I(N__4228));
    LocalMux I__867 (
            .O(N__4231),
            .I(N__4225));
    Sp12to4 I__866 (
            .O(N__4228),
            .I(N__4221));
    Span4Mux_v I__865 (
            .O(N__4225),
            .I(N__4218));
    InMux I__864 (
            .O(N__4224),
            .I(N__4215));
    Span12Mux_v I__863 (
            .O(N__4221),
            .I(N__4212));
    Sp12to4 I__862 (
            .O(N__4218),
            .I(N__4207));
    LocalMux I__861 (
            .O(N__4215),
            .I(N__4207));
    Span12Mux_h I__860 (
            .O(N__4212),
            .I(N__4204));
    Span12Mux_h I__859 (
            .O(N__4207),
            .I(N__4201));
    Odrv12 I__858 (
            .O(N__4204),
            .I(D_UM_AMIGA_in_2));
    Odrv12 I__857 (
            .O(N__4201),
            .I(D_UM_AMIGA_in_2));
    InMux I__856 (
            .O(N__4196),
            .I(N__4193));
    LocalMux I__855 (
            .O(N__4193),
            .I(N__4190));
    Odrv4 I__854 (
            .O(N__4190),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ));
    CascadeMux I__853 (
            .O(N__4187),
            .I(\U111_CYCLE_SM.un3_LW_CYCLE_START_cascade_ ));
    CascadeMux I__852 (
            .O(N__4184),
            .I(N__4181));
    InMux I__851 (
            .O(N__4181),
            .I(N__4178));
    LocalMux I__850 (
            .O(N__4178),
            .I(N__4175));
    Span4Mux_h I__849 (
            .O(N__4175),
            .I(N__4172));
    Sp12to4 I__848 (
            .O(N__4172),
            .I(N__4169));
    Odrv12 I__847 (
            .O(N__4169),
            .I(TS_CPUn_c));
    InMux I__846 (
            .O(N__4166),
            .I(N__4163));
    LocalMux I__845 (
            .O(N__4163),
            .I(N__4160));
    Span4Mux_v I__844 (
            .O(N__4160),
            .I(N__4157));
    Sp12to4 I__843 (
            .O(N__4157),
            .I(N__4154));
    Span12Mux_h I__842 (
            .O(N__4154),
            .I(N__4151));
    Odrv12 I__841 (
            .O(N__4151),
            .I(D_UU_040_in_2));
    CascadeMux I__840 (
            .O(N__4148),
            .I(N__4145));
    InMux I__839 (
            .O(N__4145),
            .I(N__4141));
    IoInMux I__838 (
            .O(N__4144),
            .I(N__4138));
    LocalMux I__837 (
            .O(N__4141),
            .I(N__4135));
    LocalMux I__836 (
            .O(N__4138),
            .I(N__4132));
    Sp12to4 I__835 (
            .O(N__4135),
            .I(N__4129));
    Span12Mux_s9_h I__834 (
            .O(N__4132),
            .I(N__4126));
    Span12Mux_v I__833 (
            .O(N__4129),
            .I(N__4123));
    Span12Mux_v I__832 (
            .O(N__4126),
            .I(N__4120));
    Span12Mux_v I__831 (
            .O(N__4123),
            .I(N__4117));
    Span12Mux_h I__830 (
            .O(N__4120),
            .I(N__4114));
    Span12Mux_h I__829 (
            .O(N__4117),
            .I(N__4111));
    Odrv12 I__828 (
            .O(N__4114),
            .I(D_LM_040_in_2));
    Odrv12 I__827 (
            .O(N__4111),
            .I(D_LM_040_in_2));
    IoInMux I__826 (
            .O(N__4106),
            .I(N__4103));
    LocalMux I__825 (
            .O(N__4103),
            .I(N__4100));
    Span12Mux_s6_v I__824 (
            .O(N__4100),
            .I(N__4097));
    Odrv12 I__823 (
            .O(N__4097),
            .I(un1_D_UU_040_2));
    CascadeMux I__822 (
            .O(N__4094),
            .I(N__4091));
    InMux I__821 (
            .O(N__4091),
            .I(N__4088));
    LocalMux I__820 (
            .O(N__4088),
            .I(N__4085));
    Span4Mux_v I__819 (
            .O(N__4085),
            .I(N__4082));
    Span4Mux_h I__818 (
            .O(N__4082),
            .I(N__4079));
    Sp12to4 I__817 (
            .O(N__4079),
            .I(N__4076));
    Span12Mux_h I__816 (
            .O(N__4076),
            .I(N__4073));
    Odrv12 I__815 (
            .O(N__4073),
            .I(D_UU_040_in_0));
    IoInMux I__814 (
            .O(N__4070),
            .I(N__4067));
    LocalMux I__813 (
            .O(N__4067),
            .I(N__4063));
    InMux I__812 (
            .O(N__4066),
            .I(N__4060));
    IoSpan4Mux I__811 (
            .O(N__4063),
            .I(N__4057));
    LocalMux I__810 (
            .O(N__4060),
            .I(N__4054));
    Span4Mux_s2_h I__809 (
            .O(N__4057),
            .I(N__4051));
    Sp12to4 I__808 (
            .O(N__4054),
            .I(N__4048));
    Span4Mux_v I__807 (
            .O(N__4051),
            .I(N__4045));
    Span12Mux_v I__806 (
            .O(N__4048),
            .I(N__4042));
    Sp12to4 I__805 (
            .O(N__4045),
            .I(N__4039));
    Span12Mux_v I__804 (
            .O(N__4042),
            .I(N__4036));
    Span12Mux_s9_h I__803 (
            .O(N__4039),
            .I(N__4033));
    Span12Mux_h I__802 (
            .O(N__4036),
            .I(N__4030));
    Span12Mux_h I__801 (
            .O(N__4033),
            .I(N__4027));
    Odrv12 I__800 (
            .O(N__4030),
            .I(D_LM_040_in_0));
    Odrv12 I__799 (
            .O(N__4027),
            .I(D_LM_040_in_0));
    IoInMux I__798 (
            .O(N__4022),
            .I(N__4019));
    LocalMux I__797 (
            .O(N__4019),
            .I(N__4016));
    IoSpan4Mux I__796 (
            .O(N__4016),
            .I(N__4013));
    IoSpan4Mux I__795 (
            .O(N__4013),
            .I(N__4010));
    Span4Mux_s3_v I__794 (
            .O(N__4010),
            .I(N__4007));
    Odrv4 I__793 (
            .O(N__4007),
            .I(un1_D_UU_040_0));
    IoInMux I__792 (
            .O(N__4004),
            .I(N__4001));
    LocalMux I__791 (
            .O(N__4001),
            .I(N__3997));
    InMux I__790 (
            .O(N__4000),
            .I(N__3994));
    Span4Mux_s2_h I__789 (
            .O(N__3997),
            .I(N__3991));
    LocalMux I__788 (
            .O(N__3994),
            .I(N__3988));
    Span4Mux_v I__787 (
            .O(N__3991),
            .I(N__3985));
    Span12Mux_h I__786 (
            .O(N__3988),
            .I(N__3982));
    Sp12to4 I__785 (
            .O(N__3985),
            .I(N__3979));
    Span12Mux_v I__784 (
            .O(N__3982),
            .I(N__3976));
    Span12Mux_h I__783 (
            .O(N__3979),
            .I(N__3973));
    Span12Mux_v I__782 (
            .O(N__3976),
            .I(N__3970));
    Span12Mux_h I__781 (
            .O(N__3973),
            .I(N__3967));
    Odrv12 I__780 (
            .O(N__3970),
            .I(D_LL_040_in_4));
    Odrv12 I__779 (
            .O(N__3967),
            .I(D_LL_040_in_4));
    CascadeMux I__778 (
            .O(N__3962),
            .I(N__3959));
    InMux I__777 (
            .O(N__3959),
            .I(N__3956));
    LocalMux I__776 (
            .O(N__3956),
            .I(N__3953));
    Span4Mux_v I__775 (
            .O(N__3953),
            .I(N__3950));
    Span4Mux_h I__774 (
            .O(N__3950),
            .I(N__3947));
    Sp12to4 I__773 (
            .O(N__3947),
            .I(N__3944));
    Span12Mux_h I__772 (
            .O(N__3944),
            .I(N__3941));
    Odrv12 I__771 (
            .O(N__3941),
            .I(D_UM_040_in_4));
    IoInMux I__770 (
            .O(N__3938),
            .I(N__3935));
    LocalMux I__769 (
            .O(N__3935),
            .I(N__3932));
    IoSpan4Mux I__768 (
            .O(N__3932),
            .I(N__3929));
    Span4Mux_s2_h I__767 (
            .O(N__3929),
            .I(N__3926));
    Span4Mux_h I__766 (
            .O(N__3926),
            .I(N__3923));
    Span4Mux_h I__765 (
            .O(N__3923),
            .I(N__3920));
    Odrv4 I__764 (
            .O(N__3920),
            .I(un1_D_UM_040_4));
    InMux I__763 (
            .O(N__3917),
            .I(N__3914));
    LocalMux I__762 (
            .O(N__3914),
            .I(N__3911));
    Span12Mux_h I__761 (
            .O(N__3911),
            .I(N__3908));
    Odrv12 I__760 (
            .O(N__3908),
            .I(D_LM_AMIGA_in_2));
    IoInMux I__759 (
            .O(N__3905),
            .I(N__3902));
    LocalMux I__758 (
            .O(N__3902),
            .I(N__3899));
    Span12Mux_s7_h I__757 (
            .O(N__3899),
            .I(N__3896));
    Span12Mux_v I__756 (
            .O(N__3896),
            .I(N__3893));
    Odrv12 I__755 (
            .O(N__3893),
            .I(un1_D_LM_AMIGA_2));
    CascadeMux I__754 (
            .O(N__3890),
            .I(N__3887));
    InMux I__753 (
            .O(N__3887),
            .I(N__3884));
    LocalMux I__752 (
            .O(N__3884),
            .I(N__3881));
    Span12Mux_v I__751 (
            .O(N__3881),
            .I(N__3878));
    Span12Mux_h I__750 (
            .O(N__3878),
            .I(N__3875));
    Odrv12 I__749 (
            .O(N__3875),
            .I(D_LM_AMIGA_in_6));
    IoInMux I__748 (
            .O(N__3872),
            .I(N__3869));
    LocalMux I__747 (
            .O(N__3869),
            .I(N__3866));
    IoSpan4Mux I__746 (
            .O(N__3866),
            .I(N__3863));
    Sp12to4 I__745 (
            .O(N__3863),
            .I(N__3860));
    Span12Mux_s9_h I__744 (
            .O(N__3860),
            .I(N__3857));
    Odrv12 I__743 (
            .O(N__3857),
            .I(un1_D_LM_AMIGA_6));
    CascadeMux I__742 (
            .O(N__3854),
            .I(N__3851));
    InMux I__741 (
            .O(N__3851),
            .I(N__3848));
    LocalMux I__740 (
            .O(N__3848),
            .I(N__3845));
    Span4Mux_v I__739 (
            .O(N__3845),
            .I(N__3842));
    Sp12to4 I__738 (
            .O(N__3842),
            .I(N__3839));
    Span12Mux_s2_v I__737 (
            .O(N__3839),
            .I(N__3836));
    Span12Mux_h I__736 (
            .O(N__3836),
            .I(N__3833));
    Odrv12 I__735 (
            .O(N__3833),
            .I(D_UM_040_in_3));
    IoInMux I__734 (
            .O(N__3830),
            .I(N__3827));
    LocalMux I__733 (
            .O(N__3827),
            .I(N__3823));
    InMux I__732 (
            .O(N__3826),
            .I(N__3820));
    Span4Mux_s3_h I__731 (
            .O(N__3823),
            .I(N__3817));
    LocalMux I__730 (
            .O(N__3820),
            .I(N__3814));
    Sp12to4 I__729 (
            .O(N__3817),
            .I(N__3811));
    Span12Mux_h I__728 (
            .O(N__3814),
            .I(N__3808));
    Span12Mux_v I__727 (
            .O(N__3811),
            .I(N__3805));
    Span12Mux_v I__726 (
            .O(N__3808),
            .I(N__3802));
    Span12Mux_h I__725 (
            .O(N__3805),
            .I(N__3799));
    Span12Mux_v I__724 (
            .O(N__3802),
            .I(N__3796));
    Span12Mux_h I__723 (
            .O(N__3799),
            .I(N__3793));
    Odrv12 I__722 (
            .O(N__3796),
            .I(D_LL_040_in_3));
    Odrv12 I__721 (
            .O(N__3793),
            .I(D_LL_040_in_3));
    IoInMux I__720 (
            .O(N__3788),
            .I(N__3785));
    LocalMux I__719 (
            .O(N__3785),
            .I(N__3782));
    IoSpan4Mux I__718 (
            .O(N__3782),
            .I(N__3779));
    Span4Mux_s3_h I__717 (
            .O(N__3779),
            .I(N__3776));
    Span4Mux_h I__716 (
            .O(N__3776),
            .I(N__3773));
    Span4Mux_h I__715 (
            .O(N__3773),
            .I(N__3770));
    Odrv4 I__714 (
            .O(N__3770),
            .I(un1_D_UM_040_3));
    CascadeMux I__713 (
            .O(N__3767),
            .I(N__3764));
    InMux I__712 (
            .O(N__3764),
            .I(N__3761));
    LocalMux I__711 (
            .O(N__3761),
            .I(N__3758));
    Span4Mux_h I__710 (
            .O(N__3758),
            .I(N__3755));
    Sp12to4 I__709 (
            .O(N__3755),
            .I(N__3752));
    Span12Mux_v I__708 (
            .O(N__3752),
            .I(N__3749));
    Span12Mux_h I__707 (
            .O(N__3749),
            .I(N__3746));
    Odrv12 I__706 (
            .O(N__3746),
            .I(D_UU_040_in_5));
    IoInMux I__705 (
            .O(N__3743),
            .I(N__3740));
    LocalMux I__704 (
            .O(N__3740),
            .I(N__3737));
    IoSpan4Mux I__703 (
            .O(N__3737),
            .I(N__3734));
    Span4Mux_s0_h I__702 (
            .O(N__3734),
            .I(N__3731));
    Span4Mux_v I__701 (
            .O(N__3731),
            .I(N__3727));
    InMux I__700 (
            .O(N__3730),
            .I(N__3724));
    Sp12to4 I__699 (
            .O(N__3727),
            .I(N__3721));
    LocalMux I__698 (
            .O(N__3724),
            .I(N__3718));
    Span12Mux_h I__697 (
            .O(N__3721),
            .I(N__3713));
    Span12Mux_v I__696 (
            .O(N__3718),
            .I(N__3713));
    Span12Mux_h I__695 (
            .O(N__3713),
            .I(N__3710));
    Odrv12 I__694 (
            .O(N__3710),
            .I(D_LM_040_in_5));
    IoInMux I__693 (
            .O(N__3707),
            .I(N__3704));
    LocalMux I__692 (
            .O(N__3704),
            .I(N__3701));
    Span4Mux_s2_h I__691 (
            .O(N__3701),
            .I(N__3698));
    Span4Mux_h I__690 (
            .O(N__3698),
            .I(N__3695));
    Sp12to4 I__689 (
            .O(N__3695),
            .I(N__3692));
    Span12Mux_s7_v I__688 (
            .O(N__3692),
            .I(N__3689));
    Odrv12 I__687 (
            .O(N__3689),
            .I(un1_D_UU_040_5));
    CascadeMux I__686 (
            .O(N__3686),
            .I(N__3683));
    InMux I__685 (
            .O(N__3683),
            .I(N__3680));
    LocalMux I__684 (
            .O(N__3680),
            .I(N__3677));
    Span4Mux_v I__683 (
            .O(N__3677),
            .I(N__3674));
    Span4Mux_h I__682 (
            .O(N__3674),
            .I(N__3671));
    Sp12to4 I__681 (
            .O(N__3671),
            .I(N__3668));
    Span12Mux_h I__680 (
            .O(N__3668),
            .I(N__3665));
    Odrv12 I__679 (
            .O(N__3665),
            .I(D_UM_040_in_5));
    IoInMux I__678 (
            .O(N__3662),
            .I(N__3658));
    InMux I__677 (
            .O(N__3661),
            .I(N__3655));
    LocalMux I__676 (
            .O(N__3658),
            .I(N__3652));
    LocalMux I__675 (
            .O(N__3655),
            .I(N__3649));
    IoSpan4Mux I__674 (
            .O(N__3652),
            .I(N__3646));
    Span4Mux_v I__673 (
            .O(N__3649),
            .I(N__3643));
    Span4Mux_s3_h I__672 (
            .O(N__3646),
            .I(N__3640));
    Sp12to4 I__671 (
            .O(N__3643),
            .I(N__3637));
    Sp12to4 I__670 (
            .O(N__3640),
            .I(N__3634));
    Span12Mux_h I__669 (
            .O(N__3637),
            .I(N__3631));
    Span12Mux_v I__668 (
            .O(N__3634),
            .I(N__3628));
    Span12Mux_v I__667 (
            .O(N__3631),
            .I(N__3625));
    Span12Mux_h I__666 (
            .O(N__3628),
            .I(N__3622));
    Span12Mux_v I__665 (
            .O(N__3625),
            .I(N__3617));
    Span12Mux_h I__664 (
            .O(N__3622),
            .I(N__3617));
    Odrv12 I__663 (
            .O(N__3617),
            .I(D_LL_040_in_5));
    IoInMux I__662 (
            .O(N__3614),
            .I(N__3611));
    LocalMux I__661 (
            .O(N__3611),
            .I(N__3608));
    IoSpan4Mux I__660 (
            .O(N__3608),
            .I(N__3605));
    Sp12to4 I__659 (
            .O(N__3605),
            .I(N__3602));
    Span12Mux_s6_v I__658 (
            .O(N__3602),
            .I(N__3599));
    Odrv12 I__657 (
            .O(N__3599),
            .I(un1_D_UM_040_5));
    CascadeMux I__656 (
            .O(N__3596),
            .I(N__3593));
    InMux I__655 (
            .O(N__3593),
            .I(N__3590));
    LocalMux I__654 (
            .O(N__3590),
            .I(N__3587));
    Span4Mux_v I__653 (
            .O(N__3587),
            .I(N__3584));
    Sp12to4 I__652 (
            .O(N__3584),
            .I(N__3581));
    Odrv12 I__651 (
            .O(N__3581),
            .I(D_LL_AMIGA_in_6));
    IoInMux I__650 (
            .O(N__3578),
            .I(N__3575));
    LocalMux I__649 (
            .O(N__3575),
            .I(N__3572));
    Span4Mux_s2_h I__648 (
            .O(N__3572),
            .I(N__3569));
    Span4Mux_v I__647 (
            .O(N__3569),
            .I(N__3566));
    Span4Mux_v I__646 (
            .O(N__3566),
            .I(N__3563));
    Sp12to4 I__645 (
            .O(N__3563),
            .I(N__3560));
    Span12Mux_s11_h I__644 (
            .O(N__3560),
            .I(N__3557));
    Odrv12 I__643 (
            .O(N__3557),
            .I(un1_D_LL_AMIGA_6));
    InMux I__642 (
            .O(N__3554),
            .I(N__3551));
    LocalMux I__641 (
            .O(N__3551),
            .I(N__3548));
    Span4Mux_v I__640 (
            .O(N__3548),
            .I(N__3545));
    Sp12to4 I__639 (
            .O(N__3545),
            .I(N__3542));
    Odrv12 I__638 (
            .O(N__3542),
            .I(D_LM_AMIGA_in_5));
    IoInMux I__637 (
            .O(N__3539),
            .I(N__3536));
    LocalMux I__636 (
            .O(N__3536),
            .I(N__3533));
    IoSpan4Mux I__635 (
            .O(N__3533),
            .I(N__3530));
    Sp12to4 I__634 (
            .O(N__3530),
            .I(N__3527));
    Span12Mux_s9_h I__633 (
            .O(N__3527),
            .I(N__3524));
    Span12Mux_h I__632 (
            .O(N__3524),
            .I(N__3521));
    Odrv12 I__631 (
            .O(N__3521),
            .I(un1_D_LM_AMIGA_5));
    CascadeMux I__630 (
            .O(N__3518),
            .I(N__3515));
    InMux I__629 (
            .O(N__3515),
            .I(N__3512));
    LocalMux I__628 (
            .O(N__3512),
            .I(N__3509));
    Span4Mux_v I__627 (
            .O(N__3509),
            .I(N__3506));
    Sp12to4 I__626 (
            .O(N__3506),
            .I(N__3503));
    Odrv12 I__625 (
            .O(N__3503),
            .I(D_LM_AMIGA_in_7));
    IoInMux I__624 (
            .O(N__3500),
            .I(N__3497));
    LocalMux I__623 (
            .O(N__3497),
            .I(N__3494));
    Span12Mux_s4_h I__622 (
            .O(N__3494),
            .I(N__3491));
    Span12Mux_h I__621 (
            .O(N__3491),
            .I(N__3488));
    Odrv12 I__620 (
            .O(N__3488),
            .I(un1_D_LM_AMIGA_7));
    IoInMux I__619 (
            .O(N__3485),
            .I(N__3482));
    LocalMux I__618 (
            .O(N__3482),
            .I(N__3479));
    Odrv12 I__617 (
            .O(N__3479),
            .I(TSn_c));
    InMux I__616 (
            .O(N__3476),
            .I(N__3473));
    LocalMux I__615 (
            .O(N__3473),
            .I(N__3470));
    Span4Mux_v I__614 (
            .O(N__3470),
            .I(N__3467));
    Span4Mux_h I__613 (
            .O(N__3467),
            .I(N__3464));
    Span4Mux_h I__612 (
            .O(N__3464),
            .I(N__3461));
    Odrv4 I__611 (
            .O(N__3461),
            .I(D_LL_AMIGA_in_0));
    IoInMux I__610 (
            .O(N__3458),
            .I(N__3455));
    LocalMux I__609 (
            .O(N__3455),
            .I(N__3452));
    IoSpan4Mux I__608 (
            .O(N__3452),
            .I(N__3449));
    IoSpan4Mux I__607 (
            .O(N__3449),
            .I(N__3446));
    Sp12to4 I__606 (
            .O(N__3446),
            .I(N__3443));
    Span12Mux_s9_h I__605 (
            .O(N__3443),
            .I(N__3440));
    Odrv12 I__604 (
            .O(N__3440),
            .I(un1_D_LL_AMIGA_0));
    InMux I__603 (
            .O(N__3437),
            .I(N__3434));
    LocalMux I__602 (
            .O(N__3434),
            .I(N__3431));
    Span4Mux_v I__601 (
            .O(N__3431),
            .I(N__3428));
    Sp12to4 I__600 (
            .O(N__3428),
            .I(N__3425));
    Span12Mux_h I__599 (
            .O(N__3425),
            .I(N__3422));
    Odrv12 I__598 (
            .O(N__3422),
            .I(D_UU_040_in_4));
    IoInMux I__597 (
            .O(N__3419),
            .I(N__3416));
    LocalMux I__596 (
            .O(N__3416),
            .I(N__3413));
    Span4Mux_s1_h I__595 (
            .O(N__3413),
            .I(N__3409));
    InMux I__594 (
            .O(N__3412),
            .I(N__3406));
    Sp12to4 I__593 (
            .O(N__3409),
            .I(N__3403));
    LocalMux I__592 (
            .O(N__3406),
            .I(N__3400));
    Span12Mux_v I__591 (
            .O(N__3403),
            .I(N__3397));
    Span12Mux_h I__590 (
            .O(N__3400),
            .I(N__3394));
    Span12Mux_h I__589 (
            .O(N__3397),
            .I(N__3391));
    Span12Mux_v I__588 (
            .O(N__3394),
            .I(N__3388));
    Span12Mux_h I__587 (
            .O(N__3391),
            .I(N__3385));
    Span12Mux_h I__586 (
            .O(N__3388),
            .I(N__3382));
    Odrv12 I__585 (
            .O(N__3385),
            .I(D_LM_040_in_4));
    Odrv12 I__584 (
            .O(N__3382),
            .I(D_LM_040_in_4));
    IoInMux I__583 (
            .O(N__3377),
            .I(N__3374));
    LocalMux I__582 (
            .O(N__3374),
            .I(N__3371));
    Span4Mux_s2_v I__581 (
            .O(N__3371),
            .I(N__3368));
    Span4Mux_h I__580 (
            .O(N__3368),
            .I(N__3365));
    Span4Mux_v I__579 (
            .O(N__3365),
            .I(N__3362));
    Odrv4 I__578 (
            .O(N__3362),
            .I(un1_D_UU_040_4));
    InMux I__577 (
            .O(N__3359),
            .I(N__3356));
    LocalMux I__576 (
            .O(N__3356),
            .I(N__3353));
    Span4Mux_v I__575 (
            .O(N__3353),
            .I(N__3350));
    Sp12to4 I__574 (
            .O(N__3350),
            .I(N__3347));
    Span12Mux_h I__573 (
            .O(N__3347),
            .I(N__3344));
    Odrv12 I__572 (
            .O(N__3344),
            .I(D_LL_AMIGA_in_1));
    IoInMux I__571 (
            .O(N__3341),
            .I(N__3338));
    LocalMux I__570 (
            .O(N__3338),
            .I(N__3335));
    IoSpan4Mux I__569 (
            .O(N__3335),
            .I(N__3332));
    IoSpan4Mux I__568 (
            .O(N__3332),
            .I(N__3329));
    Span4Mux_s2_h I__567 (
            .O(N__3329),
            .I(N__3326));
    Sp12to4 I__566 (
            .O(N__3326),
            .I(N__3323));
    Span12Mux_s11_h I__565 (
            .O(N__3323),
            .I(N__3320));
    Odrv12 I__564 (
            .O(N__3320),
            .I(un1_D_LL_AMIGA_1));
    InMux I__563 (
            .O(N__3317),
            .I(N__3314));
    LocalMux I__562 (
            .O(N__3314),
            .I(N__3311));
    Span4Mux_v I__561 (
            .O(N__3311),
            .I(N__3308));
    Sp12to4 I__560 (
            .O(N__3308),
            .I(N__3305));
    Span12Mux_h I__559 (
            .O(N__3305),
            .I(N__3302));
    Odrv12 I__558 (
            .O(N__3302),
            .I(D_LL_AMIGA_in_2));
    IoInMux I__557 (
            .O(N__3299),
            .I(N__3296));
    LocalMux I__556 (
            .O(N__3296),
            .I(N__3293));
    IoSpan4Mux I__555 (
            .O(N__3293),
            .I(N__3290));
    Sp12to4 I__554 (
            .O(N__3290),
            .I(N__3287));
    Span12Mux_s7_h I__553 (
            .O(N__3287),
            .I(N__3284));
    Span12Mux_h I__552 (
            .O(N__3284),
            .I(N__3281));
    Odrv12 I__551 (
            .O(N__3281),
            .I(un1_D_LL_AMIGA_2));
    InMux I__550 (
            .O(N__3278),
            .I(N__3275));
    LocalMux I__549 (
            .O(N__3275),
            .I(N__3272));
    Span4Mux_v I__548 (
            .O(N__3272),
            .I(N__3269));
    Sp12to4 I__547 (
            .O(N__3269),
            .I(N__3266));
    Span12Mux_h I__546 (
            .O(N__3266),
            .I(N__3263));
    Odrv12 I__545 (
            .O(N__3263),
            .I(D_LM_AMIGA_in_0));
    IoInMux I__544 (
            .O(N__3260),
            .I(N__3257));
    LocalMux I__543 (
            .O(N__3257),
            .I(N__3254));
    Span12Mux_s7_h I__542 (
            .O(N__3254),
            .I(N__3251));
    Span12Mux_h I__541 (
            .O(N__3251),
            .I(N__3248));
    Odrv12 I__540 (
            .O(N__3248),
            .I(un1_D_LM_AMIGA_0));
    CascadeMux I__539 (
            .O(N__3245),
            .I(N__3242));
    InMux I__538 (
            .O(N__3242),
            .I(N__3239));
    LocalMux I__537 (
            .O(N__3239),
            .I(N__3236));
    Span12Mux_h I__536 (
            .O(N__3236),
            .I(N__3233));
    Span12Mux_h I__535 (
            .O(N__3233),
            .I(N__3230));
    Odrv12 I__534 (
            .O(N__3230),
            .I(D_UM_040_in_2));
    InMux I__533 (
            .O(N__3227),
            .I(N__3223));
    IoInMux I__532 (
            .O(N__3226),
            .I(N__3220));
    LocalMux I__531 (
            .O(N__3223),
            .I(N__3217));
    LocalMux I__530 (
            .O(N__3220),
            .I(N__3214));
    Span4Mux_v I__529 (
            .O(N__3217),
            .I(N__3211));
    Span4Mux_s1_h I__528 (
            .O(N__3214),
            .I(N__3208));
    Sp12to4 I__527 (
            .O(N__3211),
            .I(N__3205));
    Sp12to4 I__526 (
            .O(N__3208),
            .I(N__3202));
    Span12Mux_h I__525 (
            .O(N__3205),
            .I(N__3199));
    Span12Mux_v I__524 (
            .O(N__3202),
            .I(N__3196));
    Span12Mux_v I__523 (
            .O(N__3199),
            .I(N__3193));
    Span12Mux_h I__522 (
            .O(N__3196),
            .I(N__3190));
    Span12Mux_h I__521 (
            .O(N__3193),
            .I(N__3187));
    Span12Mux_h I__520 (
            .O(N__3190),
            .I(N__3184));
    Odrv12 I__519 (
            .O(N__3187),
            .I(D_LL_040_in_2));
    Odrv12 I__518 (
            .O(N__3184),
            .I(D_LL_040_in_2));
    IoInMux I__517 (
            .O(N__3179),
            .I(N__3176));
    LocalMux I__516 (
            .O(N__3176),
            .I(N__3173));
    Span4Mux_s3_h I__515 (
            .O(N__3173),
            .I(N__3170));
    Span4Mux_v I__514 (
            .O(N__3170),
            .I(N__3167));
    Odrv4 I__513 (
            .O(N__3167),
            .I(un1_D_UM_040_2));
    InMux I__512 (
            .O(N__3164),
            .I(N__3160));
    IoInMux I__511 (
            .O(N__3163),
            .I(N__3157));
    LocalMux I__510 (
            .O(N__3160),
            .I(N__3154));
    LocalMux I__509 (
            .O(N__3157),
            .I(N__3151));
    Sp12to4 I__508 (
            .O(N__3154),
            .I(N__3148));
    Span4Mux_s3_h I__507 (
            .O(N__3151),
            .I(N__3145));
    Span12Mux_v I__506 (
            .O(N__3148),
            .I(N__3142));
    Sp12to4 I__505 (
            .O(N__3145),
            .I(N__3139));
    Span12Mux_v I__504 (
            .O(N__3142),
            .I(N__3136));
    Span12Mux_v I__503 (
            .O(N__3139),
            .I(N__3133));
    Span12Mux_h I__502 (
            .O(N__3136),
            .I(N__3130));
    Span12Mux_h I__501 (
            .O(N__3133),
            .I(N__3127));
    Span12Mux_h I__500 (
            .O(N__3130),
            .I(N__3124));
    Span12Mux_h I__499 (
            .O(N__3127),
            .I(N__3121));
    Odrv12 I__498 (
            .O(N__3124),
            .I(D_LL_040_in_1));
    Odrv12 I__497 (
            .O(N__3121),
            .I(D_LL_040_in_1));
    CascadeMux I__496 (
            .O(N__3116),
            .I(N__3113));
    InMux I__495 (
            .O(N__3113),
            .I(N__3110));
    LocalMux I__494 (
            .O(N__3110),
            .I(N__3107));
    Span4Mux_h I__493 (
            .O(N__3107),
            .I(N__3104));
    Sp12to4 I__492 (
            .O(N__3104),
            .I(N__3101));
    Span12Mux_v I__491 (
            .O(N__3101),
            .I(N__3098));
    Span12Mux_h I__490 (
            .O(N__3098),
            .I(N__3095));
    Odrv12 I__489 (
            .O(N__3095),
            .I(D_UM_040_in_1));
    IoInMux I__488 (
            .O(N__3092),
            .I(N__3089));
    LocalMux I__487 (
            .O(N__3089),
            .I(N__3086));
    Span4Mux_s2_h I__486 (
            .O(N__3086),
            .I(N__3083));
    Span4Mux_h I__485 (
            .O(N__3083),
            .I(N__3080));
    Odrv4 I__484 (
            .O(N__3080),
            .I(un1_D_UM_040_1));
    IoInMux I__483 (
            .O(N__3077),
            .I(N__3073));
    InMux I__482 (
            .O(N__3076),
            .I(N__3070));
    LocalMux I__481 (
            .O(N__3073),
            .I(N__3067));
    LocalMux I__480 (
            .O(N__3070),
            .I(N__3064));
    IoSpan4Mux I__479 (
            .O(N__3067),
            .I(N__3061));
    Sp12to4 I__478 (
            .O(N__3064),
            .I(N__3058));
    Span4Mux_s3_h I__477 (
            .O(N__3061),
            .I(N__3055));
    Span12Mux_v I__476 (
            .O(N__3058),
            .I(N__3052));
    Sp12to4 I__475 (
            .O(N__3055),
            .I(N__3049));
    Span12Mux_v I__474 (
            .O(N__3052),
            .I(N__3046));
    Span12Mux_v I__473 (
            .O(N__3049),
            .I(N__3043));
    Span12Mux_h I__472 (
            .O(N__3046),
            .I(N__3040));
    Span12Mux_h I__471 (
            .O(N__3043),
            .I(N__3037));
    Span12Mux_h I__470 (
            .O(N__3040),
            .I(N__3034));
    Span12Mux_h I__469 (
            .O(N__3037),
            .I(N__3031));
    Odrv12 I__468 (
            .O(N__3034),
            .I(D_LL_040_in_7));
    Odrv12 I__467 (
            .O(N__3031),
            .I(D_LL_040_in_7));
    CascadeMux I__466 (
            .O(N__3026),
            .I(N__3023));
    InMux I__465 (
            .O(N__3023),
            .I(N__3020));
    LocalMux I__464 (
            .O(N__3020),
            .I(N__3017));
    Span4Mux_v I__463 (
            .O(N__3017),
            .I(N__3014));
    Span4Mux_v I__462 (
            .O(N__3014),
            .I(N__3011));
    Sp12to4 I__461 (
            .O(N__3011),
            .I(N__3008));
    Span12Mux_h I__460 (
            .O(N__3008),
            .I(N__3005));
    Span12Mux_h I__459 (
            .O(N__3005),
            .I(N__3002));
    Odrv12 I__458 (
            .O(N__3002),
            .I(D_UM_040_in_7));
    IoInMux I__457 (
            .O(N__2999),
            .I(N__2996));
    LocalMux I__456 (
            .O(N__2996),
            .I(N__2993));
    Span4Mux_s1_h I__455 (
            .O(N__2993),
            .I(N__2990));
    Span4Mux_h I__454 (
            .O(N__2990),
            .I(N__2987));
    Span4Mux_v I__453 (
            .O(N__2987),
            .I(N__2984));
    Odrv4 I__452 (
            .O(N__2984),
            .I(un1_D_UM_040_7));
    InMux I__451 (
            .O(N__2981),
            .I(N__2978));
    LocalMux I__450 (
            .O(N__2978),
            .I(N__2975));
    Sp12to4 I__449 (
            .O(N__2975),
            .I(N__2972));
    Span12Mux_v I__448 (
            .O(N__2972),
            .I(N__2969));
    Span12Mux_h I__447 (
            .O(N__2969),
            .I(N__2966));
    Span12Mux_h I__446 (
            .O(N__2966),
            .I(N__2963));
    Odrv12 I__445 (
            .O(N__2963),
            .I(D_UU_040_in_1));
    CascadeMux I__444 (
            .O(N__2960),
            .I(N__2957));
    InMux I__443 (
            .O(N__2957),
            .I(N__2953));
    IoInMux I__442 (
            .O(N__2956),
            .I(N__2950));
    LocalMux I__441 (
            .O(N__2953),
            .I(N__2947));
    LocalMux I__440 (
            .O(N__2950),
            .I(N__2944));
    Sp12to4 I__439 (
            .O(N__2947),
            .I(N__2941));
    Span4Mux_s3_h I__438 (
            .O(N__2944),
            .I(N__2938));
    Span12Mux_v I__437 (
            .O(N__2941),
            .I(N__2935));
    Sp12to4 I__436 (
            .O(N__2938),
            .I(N__2932));
    Span12Mux_v I__435 (
            .O(N__2935),
            .I(N__2929));
    Span12Mux_v I__434 (
            .O(N__2932),
            .I(N__2926));
    Span12Mux_h I__433 (
            .O(N__2929),
            .I(N__2923));
    Span12Mux_h I__432 (
            .O(N__2926),
            .I(N__2920));
    Span12Mux_h I__431 (
            .O(N__2923),
            .I(N__2917));
    Span12Mux_h I__430 (
            .O(N__2920),
            .I(N__2914));
    Odrv12 I__429 (
            .O(N__2917),
            .I(D_LM_040_in_1));
    Odrv12 I__428 (
            .O(N__2914),
            .I(D_LM_040_in_1));
    IoInMux I__427 (
            .O(N__2909),
            .I(N__2906));
    LocalMux I__426 (
            .O(N__2906),
            .I(N__2903));
    Span4Mux_s2_h I__425 (
            .O(N__2903),
            .I(N__2900));
    Span4Mux_h I__424 (
            .O(N__2900),
            .I(N__2897));
    Odrv4 I__423 (
            .O(N__2897),
            .I(un1_D_UU_040_1));
    InMux I__422 (
            .O(N__2894),
            .I(N__2891));
    LocalMux I__421 (
            .O(N__2891),
            .I(N__2888));
    Odrv12 I__420 (
            .O(N__2888),
            .I(D_LM_AMIGA_in_3));
    IoInMux I__419 (
            .O(N__2885),
            .I(N__2882));
    LocalMux I__418 (
            .O(N__2882),
            .I(N__2879));
    Span4Mux_s2_h I__417 (
            .O(N__2879),
            .I(N__2876));
    Sp12to4 I__416 (
            .O(N__2876),
            .I(N__2873));
    Span12Mux_v I__415 (
            .O(N__2873),
            .I(N__2870));
    Span12Mux_h I__414 (
            .O(N__2870),
            .I(N__2867));
    Odrv12 I__413 (
            .O(N__2867),
            .I(un1_D_LM_AMIGA_3));
    IoInMux I__412 (
            .O(N__2864),
            .I(N__2861));
    LocalMux I__411 (
            .O(N__2861),
            .I(N__2858));
    IoSpan4Mux I__410 (
            .O(N__2858),
            .I(N__2854));
    InMux I__409 (
            .O(N__2857),
            .I(N__2851));
    Span4Mux_s2_h I__408 (
            .O(N__2854),
            .I(N__2848));
    LocalMux I__407 (
            .O(N__2851),
            .I(N__2845));
    Sp12to4 I__406 (
            .O(N__2848),
            .I(N__2842));
    Span4Mux_v I__405 (
            .O(N__2845),
            .I(N__2839));
    Span12Mux_h I__404 (
            .O(N__2842),
            .I(N__2836));
    Sp12to4 I__403 (
            .O(N__2839),
            .I(N__2833));
    Span12Mux_h I__402 (
            .O(N__2836),
            .I(N__2830));
    Span12Mux_h I__401 (
            .O(N__2833),
            .I(N__2827));
    Odrv12 I__400 (
            .O(N__2830),
            .I(D_LM_040_in_7));
    Odrv12 I__399 (
            .O(N__2827),
            .I(D_LM_040_in_7));
    CascadeMux I__398 (
            .O(N__2822),
            .I(N__2819));
    InMux I__397 (
            .O(N__2819),
            .I(N__2816));
    LocalMux I__396 (
            .O(N__2816),
            .I(N__2813));
    Span4Mux_v I__395 (
            .O(N__2813),
            .I(N__2810));
    Sp12to4 I__394 (
            .O(N__2810),
            .I(N__2807));
    Span12Mux_h I__393 (
            .O(N__2807),
            .I(N__2804));
    Span12Mux_h I__392 (
            .O(N__2804),
            .I(N__2801));
    Odrv12 I__391 (
            .O(N__2801),
            .I(D_UU_040_in_7));
    IoInMux I__390 (
            .O(N__2798),
            .I(N__2795));
    LocalMux I__389 (
            .O(N__2795),
            .I(N__2792));
    Span4Mux_s2_v I__388 (
            .O(N__2792),
            .I(N__2789));
    Span4Mux_h I__387 (
            .O(N__2789),
            .I(N__2786));
    Span4Mux_v I__386 (
            .O(N__2786),
            .I(N__2783));
    Odrv4 I__385 (
            .O(N__2783),
            .I(un1_D_UU_040_7));
    IoInMux I__384 (
            .O(N__2780),
            .I(N__2777));
    LocalMux I__383 (
            .O(N__2777),
            .I(N__2773));
    InMux I__382 (
            .O(N__2776),
            .I(N__2770));
    IoSpan4Mux I__381 (
            .O(N__2773),
            .I(N__2767));
    LocalMux I__380 (
            .O(N__2770),
            .I(N__2764));
    IoSpan4Mux I__379 (
            .O(N__2767),
            .I(N__2761));
    Span4Mux_v I__378 (
            .O(N__2764),
            .I(N__2758));
    Span4Mux_s2_h I__377 (
            .O(N__2761),
            .I(N__2755));
    Sp12to4 I__376 (
            .O(N__2758),
            .I(N__2752));
    Sp12to4 I__375 (
            .O(N__2755),
            .I(N__2749));
    Span12Mux_v I__374 (
            .O(N__2752),
            .I(N__2746));
    Span12Mux_h I__373 (
            .O(N__2749),
            .I(N__2743));
    Span12Mux_h I__372 (
            .O(N__2746),
            .I(N__2740));
    Span12Mux_h I__371 (
            .O(N__2743),
            .I(N__2737));
    Odrv12 I__370 (
            .O(N__2740),
            .I(D_LM_040_in_3));
    Odrv12 I__369 (
            .O(N__2737),
            .I(D_LM_040_in_3));
    CascadeMux I__368 (
            .O(N__2732),
            .I(N__2729));
    InMux I__367 (
            .O(N__2729),
            .I(N__2726));
    LocalMux I__366 (
            .O(N__2726),
            .I(N__2723));
    Span4Mux_v I__365 (
            .O(N__2723),
            .I(N__2720));
    Sp12to4 I__364 (
            .O(N__2720),
            .I(N__2717));
    Span12Mux_h I__363 (
            .O(N__2717),
            .I(N__2714));
    Span12Mux_h I__362 (
            .O(N__2714),
            .I(N__2711));
    Odrv12 I__361 (
            .O(N__2711),
            .I(D_UU_040_in_3));
    IoInMux I__360 (
            .O(N__2708),
            .I(N__2705));
    LocalMux I__359 (
            .O(N__2705),
            .I(N__2702));
    IoSpan4Mux I__358 (
            .O(N__2702),
            .I(N__2699));
    Span4Mux_s2_v I__357 (
            .O(N__2699),
            .I(N__2696));
    Span4Mux_v I__356 (
            .O(N__2696),
            .I(N__2693));
    Odrv4 I__355 (
            .O(N__2693),
            .I(un1_D_UU_040_3));
    IoInMux I__354 (
            .O(N__2690),
            .I(N__2686));
    IoInMux I__353 (
            .O(N__2689),
            .I(N__2683));
    LocalMux I__352 (
            .O(N__2686),
            .I(N__2676));
    LocalMux I__351 (
            .O(N__2683),
            .I(N__2676));
    IoInMux I__350 (
            .O(N__2682),
            .I(N__2673));
    IoInMux I__349 (
            .O(N__2681),
            .I(N__2670));
    IoSpan4Mux I__348 (
            .O(N__2676),
            .I(N__2661));
    LocalMux I__347 (
            .O(N__2673),
            .I(N__2661));
    LocalMux I__346 (
            .O(N__2670),
            .I(N__2661));
    IoInMux I__345 (
            .O(N__2669),
            .I(N__2658));
    IoInMux I__344 (
            .O(N__2668),
            .I(N__2655));
    IoSpan4Mux I__343 (
            .O(N__2661),
            .I(N__2648));
    LocalMux I__342 (
            .O(N__2658),
            .I(N__2648));
    LocalMux I__341 (
            .O(N__2655),
            .I(N__2648));
    IoSpan4Mux I__340 (
            .O(N__2648),
            .I(N__2639));
    IoInMux I__339 (
            .O(N__2647),
            .I(N__2636));
    IoInMux I__338 (
            .O(N__2646),
            .I(N__2626));
    IoInMux I__337 (
            .O(N__2645),
            .I(N__2623));
    IoInMux I__336 (
            .O(N__2644),
            .I(N__2620));
    IoInMux I__335 (
            .O(N__2643),
            .I(N__2617));
    IoInMux I__334 (
            .O(N__2642),
            .I(N__2614));
    IoSpan4Mux I__333 (
            .O(N__2639),
            .I(N__2609));
    LocalMux I__332 (
            .O(N__2636),
            .I(N__2609));
    IoInMux I__331 (
            .O(N__2635),
            .I(N__2606));
    IoInMux I__330 (
            .O(N__2634),
            .I(N__2603));
    IoInMux I__329 (
            .O(N__2633),
            .I(N__2600));
    IoInMux I__328 (
            .O(N__2632),
            .I(N__2597));
    IoInMux I__327 (
            .O(N__2631),
            .I(N__2590));
    IoInMux I__326 (
            .O(N__2630),
            .I(N__2587));
    IoInMux I__325 (
            .O(N__2629),
            .I(N__2584));
    LocalMux I__324 (
            .O(N__2626),
            .I(N__2575));
    LocalMux I__323 (
            .O(N__2623),
            .I(N__2575));
    LocalMux I__322 (
            .O(N__2620),
            .I(N__2575));
    LocalMux I__321 (
            .O(N__2617),
            .I(N__2575));
    LocalMux I__320 (
            .O(N__2614),
            .I(N__2570));
    IoSpan4Mux I__319 (
            .O(N__2609),
            .I(N__2556));
    LocalMux I__318 (
            .O(N__2606),
            .I(N__2556));
    LocalMux I__317 (
            .O(N__2603),
            .I(N__2556));
    LocalMux I__316 (
            .O(N__2600),
            .I(N__2556));
    LocalMux I__315 (
            .O(N__2597),
            .I(N__2556));
    IoInMux I__314 (
            .O(N__2596),
            .I(N__2553));
    IoInMux I__313 (
            .O(N__2595),
            .I(N__2550));
    IoInMux I__312 (
            .O(N__2594),
            .I(N__2547));
    IoInMux I__311 (
            .O(N__2593),
            .I(N__2544));
    LocalMux I__310 (
            .O(N__2590),
            .I(N__2535));
    LocalMux I__309 (
            .O(N__2587),
            .I(N__2535));
    LocalMux I__308 (
            .O(N__2584),
            .I(N__2535));
    IoSpan4Mux I__307 (
            .O(N__2575),
            .I(N__2535));
    IoInMux I__306 (
            .O(N__2574),
            .I(N__2532));
    IoInMux I__305 (
            .O(N__2573),
            .I(N__2529));
    IoSpan4Mux I__304 (
            .O(N__2570),
            .I(N__2526));
    IoInMux I__303 (
            .O(N__2569),
            .I(N__2522));
    IoInMux I__302 (
            .O(N__2568),
            .I(N__2519));
    IoInMux I__301 (
            .O(N__2567),
            .I(N__2516));
    IoSpan4Mux I__300 (
            .O(N__2556),
            .I(N__2508));
    LocalMux I__299 (
            .O(N__2553),
            .I(N__2508));
    LocalMux I__298 (
            .O(N__2550),
            .I(N__2508));
    LocalMux I__297 (
            .O(N__2547),
            .I(N__2497));
    LocalMux I__296 (
            .O(N__2544),
            .I(N__2497));
    IoSpan4Mux I__295 (
            .O(N__2535),
            .I(N__2497));
    LocalMux I__294 (
            .O(N__2532),
            .I(N__2497));
    LocalMux I__293 (
            .O(N__2529),
            .I(N__2497));
    Span4Mux_s3_v I__292 (
            .O(N__2526),
            .I(N__2494));
    IoInMux I__291 (
            .O(N__2525),
            .I(N__2491));
    LocalMux I__290 (
            .O(N__2522),
            .I(N__2484));
    LocalMux I__289 (
            .O(N__2519),
            .I(N__2484));
    LocalMux I__288 (
            .O(N__2516),
            .I(N__2481));
    IoInMux I__287 (
            .O(N__2515),
            .I(N__2478));
    IoSpan4Mux I__286 (
            .O(N__2508),
            .I(N__2473));
    IoSpan4Mux I__285 (
            .O(N__2497),
            .I(N__2473));
    Span4Mux_v I__284 (
            .O(N__2494),
            .I(N__2468));
    LocalMux I__283 (
            .O(N__2491),
            .I(N__2468));
    IoInMux I__282 (
            .O(N__2490),
            .I(N__2465));
    IoInMux I__281 (
            .O(N__2489),
            .I(N__2462));
    Span12Mux_s9_h I__280 (
            .O(N__2484),
            .I(N__2459));
    Span12Mux_s9_h I__279 (
            .O(N__2481),
            .I(N__2456));
    LocalMux I__278 (
            .O(N__2478),
            .I(N__2453));
    Span4Mux_s2_h I__277 (
            .O(N__2473),
            .I(N__2450));
    Span4Mux_s3_v I__276 (
            .O(N__2468),
            .I(N__2447));
    LocalMux I__275 (
            .O(N__2465),
            .I(N__2442));
    LocalMux I__274 (
            .O(N__2462),
            .I(N__2442));
    Span12Mux_v I__273 (
            .O(N__2459),
            .I(N__2439));
    Span12Mux_v I__272 (
            .O(N__2456),
            .I(N__2434));
    Span12Mux_s9_h I__271 (
            .O(N__2453),
            .I(N__2434));
    Span4Mux_h I__270 (
            .O(N__2450),
            .I(N__2429));
    Span4Mux_v I__269 (
            .O(N__2447),
            .I(N__2429));
    Span12Mux_s2_h I__268 (
            .O(N__2442),
            .I(N__2426));
    Odrv12 I__267 (
            .O(N__2439),
            .I(RnW_c_i_0));
    Odrv12 I__266 (
            .O(N__2434),
            .I(RnW_c_i_0));
    Odrv4 I__265 (
            .O(N__2429),
            .I(RnW_c_i_0));
    Odrv12 I__264 (
            .O(N__2426),
            .I(RnW_c_i_0));
    InMux I__263 (
            .O(N__2417),
            .I(N__2414));
    LocalMux I__262 (
            .O(N__2414),
            .I(N__2411));
    Span4Mux_h I__261 (
            .O(N__2411),
            .I(N__2408));
    Span4Mux_v I__260 (
            .O(N__2408),
            .I(N__2405));
    Odrv4 I__259 (
            .O(N__2405),
            .I(A_040_c_0));
    IoInMux I__258 (
            .O(N__2402),
            .I(N__2399));
    LocalMux I__257 (
            .O(N__2399),
            .I(N__2396));
    Span4Mux_s2_v I__256 (
            .O(N__2396),
            .I(N__2393));
    Span4Mux_v I__255 (
            .O(N__2393),
            .I(N__2390));
    Odrv4 I__254 (
            .O(N__2390),
            .I(A_AMIGA_c_0));
    InMux I__253 (
            .O(N__2387),
            .I(N__2384));
    LocalMux I__252 (
            .O(N__2384),
            .I(N__2381));
    Span12Mux_h I__251 (
            .O(N__2381),
            .I(N__2378));
    Odrv12 I__250 (
            .O(N__2378),
            .I(A_040_c_1));
    CascadeMux I__249 (
            .O(N__2375),
            .I(A_AMIGA_c_1_cascade_));
    InMux I__248 (
            .O(N__2372),
            .I(N__2369));
    LocalMux I__247 (
            .O(N__2369),
            .I(N__2366));
    Span4Mux_v I__246 (
            .O(N__2366),
            .I(N__2363));
    Sp12to4 I__245 (
            .O(N__2363),
            .I(N__2360));
    Odrv12 I__244 (
            .O(N__2360),
            .I(D_LL_AMIGA_in_3));
    IoInMux I__243 (
            .O(N__2357),
            .I(N__2354));
    LocalMux I__242 (
            .O(N__2354),
            .I(N__2351));
    Span4Mux_s1_h I__241 (
            .O(N__2351),
            .I(N__2348));
    Sp12to4 I__240 (
            .O(N__2348),
            .I(N__2345));
    Span12Mux_s6_v I__239 (
            .O(N__2345),
            .I(N__2342));
    Span12Mux_h I__238 (
            .O(N__2342),
            .I(N__2339));
    Odrv12 I__237 (
            .O(N__2339),
            .I(un1_D_LL_AMIGA_3));
    CascadeMux I__236 (
            .O(N__2336),
            .I(N__2333));
    InMux I__235 (
            .O(N__2333),
            .I(N__2330));
    LocalMux I__234 (
            .O(N__2330),
            .I(N__2327));
    Span4Mux_v I__233 (
            .O(N__2327),
            .I(N__2324));
    Span4Mux_h I__232 (
            .O(N__2324),
            .I(N__2321));
    Odrv4 I__231 (
            .O(N__2321),
            .I(D_LL_AMIGA_in_4));
    IoInMux I__230 (
            .O(N__2318),
            .I(N__2315));
    LocalMux I__229 (
            .O(N__2315),
            .I(N__2312));
    Sp12to4 I__228 (
            .O(N__2312),
            .I(N__2309));
    Span12Mux_h I__227 (
            .O(N__2309),
            .I(N__2306));
    Span12Mux_h I__226 (
            .O(N__2306),
            .I(N__2303));
    Odrv12 I__225 (
            .O(N__2303),
            .I(un1_D_LL_AMIGA_4));
    InMux I__224 (
            .O(N__2300),
            .I(N__2297));
    LocalMux I__223 (
            .O(N__2297),
            .I(N__2294));
    Sp12to4 I__222 (
            .O(N__2294),
            .I(N__2291));
    Span12Mux_v I__221 (
            .O(N__2291),
            .I(N__2288));
    Span12Mux_h I__220 (
            .O(N__2288),
            .I(N__2285));
    Span12Mux_h I__219 (
            .O(N__2285),
            .I(N__2282));
    Odrv12 I__218 (
            .O(N__2282),
            .I(D_UM_040_in_0));
    CascadeMux I__217 (
            .O(N__2279),
            .I(N__2276));
    InMux I__216 (
            .O(N__2276),
            .I(N__2272));
    IoInMux I__215 (
            .O(N__2275),
            .I(N__2269));
    LocalMux I__214 (
            .O(N__2272),
            .I(N__2266));
    LocalMux I__213 (
            .O(N__2269),
            .I(N__2263));
    Span4Mux_v I__212 (
            .O(N__2266),
            .I(N__2260));
    IoSpan4Mux I__211 (
            .O(N__2263),
            .I(N__2257));
    Sp12to4 I__210 (
            .O(N__2260),
            .I(N__2254));
    Span4Mux_s2_h I__209 (
            .O(N__2257),
            .I(N__2251));
    Span12Mux_h I__208 (
            .O(N__2254),
            .I(N__2248));
    Sp12to4 I__207 (
            .O(N__2251),
            .I(N__2245));
    Span12Mux_v I__206 (
            .O(N__2248),
            .I(N__2242));
    Span12Mux_h I__205 (
            .O(N__2245),
            .I(N__2239));
    Span12Mux_h I__204 (
            .O(N__2242),
            .I(N__2236));
    Span12Mux_h I__203 (
            .O(N__2239),
            .I(N__2233));
    Odrv12 I__202 (
            .O(N__2236),
            .I(D_LL_040_in_0));
    Odrv12 I__201 (
            .O(N__2233),
            .I(D_LL_040_in_0));
    IoInMux I__200 (
            .O(N__2228),
            .I(N__2225));
    LocalMux I__199 (
            .O(N__2225),
            .I(N__2222));
    IoSpan4Mux I__198 (
            .O(N__2222),
            .I(N__2219));
    Span4Mux_s1_h I__197 (
            .O(N__2219),
            .I(N__2216));
    Span4Mux_h I__196 (
            .O(N__2216),
            .I(N__2213));
    Odrv4 I__195 (
            .O(N__2213),
            .I(un1_D_UM_040_0));
    INV \INVU111_CYCLE_SM.UU_LATCHED_nesr_5C  (
            .O(\INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net ),
            .I(N__5626));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_1C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_1C_net ),
            .I(N__5629));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net ),
            .I(N__5631));
    INV \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C  (
            .O(\INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net ),
            .I(N__5623));
    INV \INVU111_CYCLE_SM.CYCLE_STATE_0C  (
            .O(\INVU111_CYCLE_SM.CYCLE_STATE_0C_net ),
            .I(N__5624));
    INV \INVU111_CYCLE_SM.LW_CYCLEC  (
            .O(\INVU111_CYCLE_SM.LW_CYCLEC_net ),
            .I(N__5627));
    INV \INVU111_CYCLE_SM.UU_LATCHED_nesr_6C  (
            .O(\INVU111_CYCLE_SM.UU_LATCHED_nesr_6C_net ),
            .I(N__5625));
    INV \INVU111_CYCLE_SM.LW_CYCLE_STARTC  (
            .O(\INVU111_CYCLE_SM.LW_CYCLE_STARTC_net ),
            .I(N__5628));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_2C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_2C_net ),
            .I(N__5630));
    INV \INVU111_CYCLE_SM.TA_ENC  (
            .O(\INVU111_CYCLE_SM.TA_ENC_net ),
            .I(N__5632));
    INV \INVU111_CYCLE_SM.TSnC  (
            .O(\INVU111_CYCLE_SM.TSnC_net ),
            .I(N__5531));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_0  (
            .in0(N__7346),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2417),
            .lcout(A_AMIGA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_3  (
            .in0(N__2387),
            .in1(N__5474),
            .in2(_gnd_net_),
            .in3(N__7345),
            .lcout(A_AMIGA_c_1),
            .ltout(A_AMIGA_c_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_3_1_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_3_1_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_3_1_4 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_3_1_4  (
            .in0(N__7082),
            .in1(N__6328),
            .in2(N__2375),
            .in3(N__2372),
            .lcout(un1_D_LL_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_3_3_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_3_3_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_3_3_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_3_3_5  (
            .in0(N__6329),
            .in1(N__6842),
            .in2(N__2336),
            .in3(N__5795),
            .lcout(un1_D_LL_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_3_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_3_10_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_3_10_3  (
            .in0(N__6326),
            .in1(N__2300),
            .in2(N__2279),
            .in3(N__5796),
            .lcout(un1_D_UM_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_3_10_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_3_10_6 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_3_10_6  (
            .in0(N__5797),
            .in1(N__6327),
            .in2(N__3245),
            .in3(N__3227),
            .lcout(un1_D_UM_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_3_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_3_15_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_3_15_0  (
            .in0(N__3164),
            .in1(N__6284),
            .in2(N__3116),
            .in3(N__5851),
            .lcout(un1_D_UM_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_3_18_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_3_18_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_3_18_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_3_18_0  (
            .in0(N__3076),
            .in1(N__6266),
            .in2(N__3026),
            .in3(N__5852),
            .lcout(un1_D_UM_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_3_18_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_3_18_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_3_18_2 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_3_18_2  (
            .in0(N__2981),
            .in1(N__6267),
            .in2(N__2960),
            .in3(N__5853),
            .lcout(un1_D_UU_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_5_11_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_5_11_7 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_5_11_7  (
            .in0(N__5883),
            .in1(N__6316),
            .in2(N__4403),
            .in3(N__2894),
            .lcout(un1_D_LM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_5_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_5_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_5_20_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_5_20_3  (
            .in0(N__6292),
            .in1(N__2857),
            .in2(N__2822),
            .in3(N__5957),
            .lcout(un1_D_UU_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_5_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_5_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_5_20_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_5_20_7  (
            .in0(N__6291),
            .in1(N__2776),
            .in2(N__2732),
            .in3(N__5956),
            .lcout(un1_D_UU_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RnW_c_sbtinv_LC_6_19_3.C_ON=1'b0;
    defparam RnW_c_sbtinv_LC_6_19_3.SEQ_MODE=4'b0000;
    defparam RnW_c_sbtinv_LC_6_19_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 RnW_c_sbtinv_LC_6_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5165),
            .lcout(RnW_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_7_6_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_7_6_6 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_7_6_6  (
            .in0(N__6268),
            .in1(N__6586),
            .in2(N__3596),
            .in3(N__5913),
            .lcout(un1_D_LL_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_7_15_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_7_15_7 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_7_15_7  (
            .in0(N__3554),
            .in1(N__6237),
            .in2(N__7393),
            .in3(N__5919),
            .lcout(un1_D_LM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_7_17_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_7_17_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_7_17_3  (
            .in0(N__6681),
            .in1(N__6184),
            .in2(N__3518),
            .in3(N__5949),
            .lcout(un1_D_LM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TSn_LC_8_1_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TSn_LC_8_1_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TSn_LC_8_1_2 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U111_CYCLE_SM.TSn_LC_8_1_2  (
            .in0(N__5266),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4577),
            .lcout(TSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TSnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_8_1_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_8_1_5 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_8_1_5  (
            .in0(N__6317),
            .in1(N__3476),
            .in2(N__6530),
            .in3(N__5864),
            .lcout(un1_D_LL_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_8_20_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_8_20_6 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_8_20_6  (
            .in0(N__3437),
            .in1(N__3412),
            .in2(N__6288),
            .in3(N__5970),
            .lcout(un1_D_UU_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_9_3_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_9_3_0 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_9_3_0  (
            .in0(N__6998),
            .in1(N__6321),
            .in2(N__5940),
            .in3(N__3359),
            .lcout(un1_D_LL_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_9_3_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_9_3_5 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_9_3_5  (
            .in0(N__6322),
            .in1(N__4238),
            .in2(N__5941),
            .in3(N__3317),
            .lcout(un1_D_LL_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_9_7_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_9_7_4 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_9_7_4  (
            .in0(N__6302),
            .in1(N__6464),
            .in2(N__5966),
            .in3(N__3278),
            .lcout(un1_D_LM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_9_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_9_20_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_9_20_3  (
            .in0(N__6245),
            .in1(N__4166),
            .in2(N__4148),
            .in3(N__5983),
            .lcout(un1_D_UU_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_9_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_9_20_4 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_9_20_4  (
            .in0(N__5985),
            .in1(N__6247),
            .in2(N__4094),
            .in3(N__4066),
            .lcout(un1_D_UU_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_9_20_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_9_20_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_9_20_5  (
            .in0(N__6246),
            .in1(N__4000),
            .in2(N__3962),
            .in3(N__5984),
            .lcout(un1_D_UM_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_10_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_10_12_5 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_10_12_5  (
            .in0(N__5859),
            .in1(N__6230),
            .in2(N__4874),
            .in3(N__3917),
            .lcout(un1_D_LM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_10_16_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_10_16_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_10_16_7  (
            .in0(N__6109),
            .in1(N__4945),
            .in2(N__3890),
            .in3(N__5912),
            .lcout(un1_D_LM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_10_19_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_10_19_1 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_10_19_1  (
            .in0(N__5969),
            .in1(N__6164),
            .in2(N__3854),
            .in3(N__3826),
            .lcout(un1_D_UM_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_10_19_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_10_19_3 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_10_19_3  (
            .in0(N__5968),
            .in1(N__6163),
            .in2(N__3767),
            .in3(N__3730),
            .lcout(un1_D_UU_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_10_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_10_20_3 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_10_20_3  (
            .in0(N__5992),
            .in1(N__6229),
            .in2(N__3686),
            .in3(N__3661),
            .lcout(un1_D_UM_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_0 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_0  (
            .in0(N__4337),
            .in1(N__6269),
            .in2(N__6392),
            .in3(N__5945),
            .lcout(un1_D_LL_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_11_6_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_11_6_1 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_11_6_1  (
            .in0(N__6270),
            .in1(N__6770),
            .in2(N__5967),
            .in3(N__4295),
            .lcout(un1_D_LL_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_EN_RNO_0_LC_11_12_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_EN_RNO_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_EN_RNO_0_LC_11_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U111_CYCLE_SM.TA_EN_RNO_0_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5287),
            .lcout(\U111_CYCLE_SM.RESETn_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_11_12_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_11_12_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_11_12_2  (
            .in0(N__4196),
            .in1(N__4237),
            .in2(_gnd_net_),
            .in3(N__7304),
            .lcout(un1_D_UM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_EN_LC_11_13_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_EN_LC_11_13_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.TA_EN_LC_11_13_3 .LUT_INIT=16'b1111000011011100;
    LogicCell40 \U111_CYCLE_SM.TA_EN_LC_11_13_3  (
            .in0(N__5507),
            .in1(N__5363),
            .in2(N__4667),
            .in3(N__5405),
            .lcout(\U111_CYCLE_SM.TA_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TA_ENC_net ),
            .ce(),
            .sr(N__4247));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_11_14_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_11_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4224),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_2C_net ),
            .ce(N__7190),
            .sr(N__7143));
    defparam \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_11_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_11_15_0 .LUT_INIT=16'b1001000000000000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_11_15_0  (
            .in0(N__4496),
            .in1(N__4523),
            .in2(N__4573),
            .in3(N__4543),
            .lcout(),
            .ltout(\U111_CYCLE_SM.un3_LW_CYCLE_START_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_START_LC_11_15_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_LC_11_15_1 .LUT_INIT=16'b1010001010100000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_START_LC_11_15_1  (
            .in0(N__5309),
            .in1(N__7252),
            .in2(N__4187),
            .in3(N__5503),
            .lcout(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.LW_CYCLE_STARTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_11_15_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_11_15_2 .LUT_INIT=16'b0000001011001110;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_1_LC_11_15_2  (
            .in0(N__5544),
            .in1(N__5355),
            .in2(N__4184),
            .in3(N__5400),
            .lcout(\U111_CYCLE_SM.TS_EN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_15_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_15_6 .LUT_INIT=16'b1100110010111011;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_15_6  (
            .in0(N__5543),
            .in1(N__5354),
            .in2(_gnd_net_),
            .in3(N__5401),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_69_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_LC_11_15_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TS_EN_LC_11_15_7 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \U111_CYCLE_SM.TS_EN_LC_11_15_7  (
            .in0(N__5310),
            .in1(N__4569),
            .in2(N__4586),
            .in3(N__4583),
            .lcout(\U111_CYCLE_SM.TS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.LW_CYCLE_STARTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_11_16_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_11_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4946),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_6C_net ),
            .ce(N__7191),
            .sr(N__7139));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_16_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_16_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_16_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_16_3  (
            .in0(N__4867),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_6C_net ),
            .ce(N__7191),
            .sr(N__7139));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_11_16_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_11_16_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_11_16_7  (
            .in0(N__4393),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_6C_net ),
            .ce(N__7191),
            .sr(N__7139));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI2RET_LC_11_17_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI2RET_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI2RET_LC_11_17_1 .LUT_INIT=16'b0000000011010111;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI2RET_LC_11_17_1  (
            .in0(N__4550),
            .in1(N__4519),
            .in2(N__4495),
            .in3(N__7331),
            .lcout(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_11_17_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_17_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_17_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_11_18_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_11_18_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_11_18_1  (
            .in0(N__7333),
            .in1(N__4412),
            .in2(_gnd_net_),
            .in3(N__4392),
            .lcout(un1_D_UU_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_11_18_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_11_18_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_11_18_3  (
            .in0(N__7334),
            .in1(N__4955),
            .in2(_gnd_net_),
            .in3(N__4944),
            .lcout(un1_D_UU_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_18_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_18_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_18_7  (
            .in0(N__7332),
            .in1(N__4883),
            .in2(_gnd_net_),
            .in3(N__4866),
            .lcout(un1_D_UU_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_2.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5546),
            .lcout(GB_BUFFER_CLK40_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_12_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_12_10_3 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_12_10_3  (
            .in0(N__5926),
            .in1(N__6290),
            .in2(N__4790),
            .in3(N__6909),
            .lcout(un1_D_LM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_12_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_12_12_5 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_12_12_5  (
            .in0(N__4754),
            .in1(N__6289),
            .in2(N__4732),
            .in3(N__5860),
            .lcout(un1_D_UM_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_EN_RNI1DSB_LC_12_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_EN_RNI1DSB_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_EN_RNI1DSB_LC_12_13_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U111_CYCLE_SM.TA_EN_RNI1DSB_LC_12_13_0  (
            .in0(N__4666),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5425),
            .lcout(U111_CYCLE_SM_TAn_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_12_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_12_13_1 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_12_13_1  (
            .in0(N__4631),
            .in1(N__6265),
            .in2(N__5708),
            .in3(N__5955),
            .lcout(un1_D_LM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_LC_12_14_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_CYCLE_LC_12_14_0 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_LC_12_14_0  (
            .in0(N__5357),
            .in1(N__4592),
            .in2(N__5315),
            .in3(N__5552),
            .lcout(\U111_CYCLE_SM.LW_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.LW_CYCLEC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_12_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_12_14_5 .LUT_INIT=16'b1010001010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_12_14_5  (
            .in0(N__7251),
            .in1(N__5356),
            .in2(N__5447),
            .in3(N__5399),
            .lcout(\U111_CYCLE_SM.LW_CYCLE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_12_14_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_12_14_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__5500),
            .in2(_gnd_net_),
            .in3(N__5398),
            .lcout(\U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_15_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_15_0  (
            .in0(N__5350),
            .in1(N__5502),
            .in2(_gnd_net_),
            .in3(N__5545),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_91_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_15_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_15_1 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_15_1  (
            .in0(N__5444),
            .in1(N__5312),
            .in2(N__5510),
            .in3(N__5397),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.CYCLE_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A_OUT_RNO_0_LC_12_15_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A_OUT_RNO_0_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A_OUT_RNO_0_LC_12_15_2 .LUT_INIT=16'b1111101101010000;
    LogicCell40 \U111_CYCLE_SM.A_OUT_RNO_0_LC_12_15_2  (
            .in0(N__5395),
            .in1(N__5501),
            .in2(N__5361),
            .in3(N__5458),
            .lcout(),
            .ltout(\U111_CYCLE_SM.A_OUT_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A_OUT_LC_12_15_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A_OUT_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.A_OUT_LC_12_15_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U111_CYCLE_SM.A_OUT_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5477),
            .in3(N__5311),
            .lcout(\U111_CYCLE_SM.A_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.CYCLE_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_15_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_15_4 .LUT_INIT=16'b1101001000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_15_4  (
            .in0(N__5396),
            .in1(N__5445),
            .in2(N__5362),
            .in3(N__5314),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.CYCLE_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_12_15_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_12_15_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_12_15_5  (
            .in0(N__5446),
            .in1(N__5394),
            .in2(_gnd_net_),
            .in3(N__5346),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa ),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_12_15_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_12_15_6 .LUT_INIT=16'b0101010111110101;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_12_15_6  (
            .in0(N__5313),
            .in1(_gnd_net_),
            .in2(N__5249),
            .in3(N__5098),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0 ),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_12_15_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_12_15_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4958),
            .in3(N__6479),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_12_16_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_12_16_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_12_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5701),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net ),
            .ce(N__7188),
            .sr(N__7138));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_12_16_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_12_16_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_12_16_5  (
            .in0(N__6463),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net ),
            .ce(N__7188),
            .sr(N__7138));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_12_16_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_12_16_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_12_16_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_12_16_7  (
            .in0(N__6385),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net ),
            .ce(N__7188),
            .sr(N__7138));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_12_18_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_12_18_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_12_18_1  (
            .in0(N__7316),
            .in1(N__6473),
            .in2(_gnd_net_),
            .in3(N__6456),
            .lcout(un1_D_UU_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_12_18_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_12_18_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_12_18_7  (
            .in0(N__7315),
            .in1(N__6401),
            .in2(_gnd_net_),
            .in3(N__6384),
            .lcout(un1_D_UM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_12_20_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_12_20_0 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_12_20_0  (
            .in0(N__6244),
            .in1(N__6059),
            .in2(N__6040),
            .in3(N__5993),
            .lcout(un1_D_UU_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_12_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_12_20_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_12_20_4  (
            .in0(N__5700),
            .in1(N__5669),
            .in2(_gnd_net_),
            .in3(N__7317),
            .lcout(un1_D_UU_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_12_4.C_ON=1'b0;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_12_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_12_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_12_4 (
            .in0(N__5639),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_CLK80_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_13_12_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_13_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_13_12_6  (
            .in0(N__6488),
            .in1(N__6507),
            .in2(_gnd_net_),
            .in3(N__7286),
            .lcout(un1_D_UM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_13_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_13_12_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_13_12_7  (
            .in0(N__7287),
            .in1(N__6539),
            .in2(_gnd_net_),
            .in3(N__6582),
            .lcout(un1_D_UM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_13_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_13_14_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_13_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6587),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net ),
            .ce(N__7192),
            .sr(N__7144));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_13_14_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_13_14_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_13_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6520),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net ),
            .ce(N__7192),
            .sr(N__7144));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_13_15_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_13_15_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_13_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6996),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_1C_net ),
            .ce(N__7189),
            .sr(N__7125));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_13_15_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_13_15_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_13_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6769),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_1C_net ),
            .ce(N__7189),
            .sr(N__7125));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_13_16_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_13_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7394),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net ),
            .ce(N__7193),
            .sr(N__7145));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_13_16_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_13_16_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_13_16_2  (
            .in0(N__7081),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net ),
            .ce(N__7193),
            .sr(N__7145));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_13_16_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_13_16_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_13_16_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_13_16_4  (
            .in0(N__6838),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net ),
            .ce(N__7193),
            .sr(N__7145));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_13_16_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_13_16_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_13_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6683),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net ),
            .ce(N__7193),
            .sr(N__7145));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_13_16_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_13_16_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_13_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6914),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net ),
            .ce(N__7193),
            .sr(N__7145));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_13_17_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_13_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_13_17_2  (
            .in0(N__7322),
            .in1(N__7088),
            .in2(_gnd_net_),
            .in3(N__7080),
            .lcout(un1_D_UM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_13_17_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_13_17_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_13_17_3  (
            .in0(N__6997),
            .in1(N__6953),
            .in2(_gnd_net_),
            .in3(N__7321),
            .lcout(un1_D_UM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_13_18_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_13_18_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_13_18_4  (
            .in0(N__7323),
            .in1(N__6923),
            .in2(_gnd_net_),
            .in3(N__6910),
            .lcout(un1_D_UU_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_13_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_13_19_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_13_19_2  (
            .in0(N__7324),
            .in1(N__6851),
            .in2(_gnd_net_),
            .in3(N__6831),
            .lcout(un1_D_UM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_13_19_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_13_19_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_13_19_3  (
            .in0(N__6762),
            .in1(N__6722),
            .in2(_gnd_net_),
            .in3(N__7325),
            .lcout(un1_D_UM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_13_20_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_13_20_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_13_20_0  (
            .in0(N__7339),
            .in1(N__6692),
            .in2(_gnd_net_),
            .in3(N__6682),
            .lcout(un1_D_UU_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_13_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_13_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_13_20_3  (
            .in0(N__7403),
            .in1(N__7389),
            .in2(_gnd_net_),
            .in3(N__7338),
            .lcout(un1_D_UU_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U111_TOP

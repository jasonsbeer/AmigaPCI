// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 30 2025 11:26:14

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    CMA,
    DRA,
    SIZ,
    A,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    DBRn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    output [10:0] CMA;
    input [9:0] DRA;
    input [1:0] SIZ;
    input [20:0] A;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input DBRn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__11659;
    wire N__11658;
    wire N__11657;
    wire N__11650;
    wire N__11649;
    wire N__11648;
    wire N__11641;
    wire N__11640;
    wire N__11639;
    wire N__11632;
    wire N__11631;
    wire N__11630;
    wire N__11623;
    wire N__11622;
    wire N__11621;
    wire N__11614;
    wire N__11613;
    wire N__11612;
    wire N__11605;
    wire N__11604;
    wire N__11603;
    wire N__11596;
    wire N__11595;
    wire N__11594;
    wire N__11587;
    wire N__11586;
    wire N__11585;
    wire N__11578;
    wire N__11577;
    wire N__11576;
    wire N__11569;
    wire N__11568;
    wire N__11567;
    wire N__11560;
    wire N__11559;
    wire N__11558;
    wire N__11551;
    wire N__11550;
    wire N__11549;
    wire N__11542;
    wire N__11541;
    wire N__11540;
    wire N__11533;
    wire N__11532;
    wire N__11531;
    wire N__11524;
    wire N__11523;
    wire N__11522;
    wire N__11515;
    wire N__11514;
    wire N__11513;
    wire N__11506;
    wire N__11505;
    wire N__11504;
    wire N__11497;
    wire N__11496;
    wire N__11495;
    wire N__11488;
    wire N__11487;
    wire N__11486;
    wire N__11479;
    wire N__11478;
    wire N__11477;
    wire N__11470;
    wire N__11469;
    wire N__11468;
    wire N__11461;
    wire N__11460;
    wire N__11459;
    wire N__11452;
    wire N__11451;
    wire N__11450;
    wire N__11443;
    wire N__11442;
    wire N__11441;
    wire N__11434;
    wire N__11433;
    wire N__11432;
    wire N__11425;
    wire N__11424;
    wire N__11423;
    wire N__11416;
    wire N__11415;
    wire N__11414;
    wire N__11407;
    wire N__11406;
    wire N__11405;
    wire N__11398;
    wire N__11397;
    wire N__11396;
    wire N__11389;
    wire N__11388;
    wire N__11387;
    wire N__11380;
    wire N__11379;
    wire N__11378;
    wire N__11371;
    wire N__11370;
    wire N__11369;
    wire N__11362;
    wire N__11361;
    wire N__11360;
    wire N__11353;
    wire N__11352;
    wire N__11351;
    wire N__11344;
    wire N__11343;
    wire N__11342;
    wire N__11335;
    wire N__11334;
    wire N__11333;
    wire N__11326;
    wire N__11325;
    wire N__11324;
    wire N__11317;
    wire N__11316;
    wire N__11315;
    wire N__11308;
    wire N__11307;
    wire N__11306;
    wire N__11299;
    wire N__11298;
    wire N__11297;
    wire N__11290;
    wire N__11289;
    wire N__11288;
    wire N__11281;
    wire N__11280;
    wire N__11279;
    wire N__11272;
    wire N__11271;
    wire N__11270;
    wire N__11263;
    wire N__11262;
    wire N__11261;
    wire N__11254;
    wire N__11253;
    wire N__11252;
    wire N__11245;
    wire N__11244;
    wire N__11243;
    wire N__11236;
    wire N__11235;
    wire N__11234;
    wire N__11227;
    wire N__11226;
    wire N__11225;
    wire N__11218;
    wire N__11217;
    wire N__11216;
    wire N__11209;
    wire N__11208;
    wire N__11207;
    wire N__11200;
    wire N__11199;
    wire N__11198;
    wire N__11191;
    wire N__11190;
    wire N__11189;
    wire N__11182;
    wire N__11181;
    wire N__11180;
    wire N__11173;
    wire N__11172;
    wire N__11171;
    wire N__11164;
    wire N__11163;
    wire N__11162;
    wire N__11155;
    wire N__11154;
    wire N__11153;
    wire N__11146;
    wire N__11145;
    wire N__11144;
    wire N__11137;
    wire N__11136;
    wire N__11135;
    wire N__11128;
    wire N__11127;
    wire N__11126;
    wire N__11119;
    wire N__11118;
    wire N__11117;
    wire N__11110;
    wire N__11109;
    wire N__11108;
    wire N__11101;
    wire N__11100;
    wire N__11099;
    wire N__11092;
    wire N__11091;
    wire N__11090;
    wire N__11083;
    wire N__11082;
    wire N__11081;
    wire N__11074;
    wire N__11073;
    wire N__11072;
    wire N__11065;
    wire N__11064;
    wire N__11063;
    wire N__11056;
    wire N__11055;
    wire N__11054;
    wire N__11047;
    wire N__11046;
    wire N__11045;
    wire N__11038;
    wire N__11037;
    wire N__11036;
    wire N__11029;
    wire N__11028;
    wire N__11027;
    wire N__11020;
    wire N__11019;
    wire N__11018;
    wire N__11011;
    wire N__11010;
    wire N__11009;
    wire N__11002;
    wire N__11001;
    wire N__11000;
    wire N__10993;
    wire N__10992;
    wire N__10991;
    wire N__10984;
    wire N__10983;
    wire N__10982;
    wire N__10975;
    wire N__10974;
    wire N__10973;
    wire N__10966;
    wire N__10965;
    wire N__10964;
    wire N__10957;
    wire N__10956;
    wire N__10955;
    wire N__10948;
    wire N__10947;
    wire N__10946;
    wire N__10939;
    wire N__10938;
    wire N__10937;
    wire N__10930;
    wire N__10929;
    wire N__10928;
    wire N__10921;
    wire N__10920;
    wire N__10919;
    wire N__10912;
    wire N__10911;
    wire N__10910;
    wire N__10903;
    wire N__10902;
    wire N__10901;
    wire N__10894;
    wire N__10893;
    wire N__10892;
    wire N__10885;
    wire N__10884;
    wire N__10883;
    wire N__10876;
    wire N__10875;
    wire N__10874;
    wire N__10867;
    wire N__10866;
    wire N__10865;
    wire N__10848;
    wire N__10847;
    wire N__10846;
    wire N__10845;
    wire N__10844;
    wire N__10843;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10830;
    wire N__10823;
    wire N__10822;
    wire N__10821;
    wire N__10820;
    wire N__10819;
    wire N__10818;
    wire N__10817;
    wire N__10816;
    wire N__10815;
    wire N__10814;
    wire N__10813;
    wire N__10812;
    wire N__10809;
    wire N__10808;
    wire N__10807;
    wire N__10806;
    wire N__10805;
    wire N__10804;
    wire N__10803;
    wire N__10802;
    wire N__10801;
    wire N__10800;
    wire N__10799;
    wire N__10798;
    wire N__10795;
    wire N__10792;
    wire N__10791;
    wire N__10790;
    wire N__10789;
    wire N__10788;
    wire N__10787;
    wire N__10786;
    wire N__10785;
    wire N__10784;
    wire N__10783;
    wire N__10780;
    wire N__10777;
    wire N__10776;
    wire N__10775;
    wire N__10774;
    wire N__10773;
    wire N__10772;
    wire N__10771;
    wire N__10770;
    wire N__10769;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10666;
    wire N__10663;
    wire N__10660;
    wire N__10657;
    wire N__10654;
    wire N__10653;
    wire N__10650;
    wire N__10647;
    wire N__10644;
    wire N__10641;
    wire N__10636;
    wire N__10629;
    wire N__10628;
    wire N__10625;
    wire N__10624;
    wire N__10621;
    wire N__10620;
    wire N__10617;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10603;
    wire N__10600;
    wire N__10597;
    wire N__10596;
    wire N__10593;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10581;
    wire N__10576;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10562;
    wire N__10559;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10545;
    wire N__10544;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10534;
    wire N__10531;
    wire N__10530;
    wire N__10525;
    wire N__10522;
    wire N__10519;
    wire N__10518;
    wire N__10511;
    wire N__10508;
    wire N__10503;
    wire N__10500;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10476;
    wire N__10473;
    wire N__10470;
    wire N__10467;
    wire N__10464;
    wire N__10461;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10443;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10419;
    wire N__10416;
    wire N__10415;
    wire N__10414;
    wire N__10409;
    wire N__10408;
    wire N__10405;
    wire N__10402;
    wire N__10399;
    wire N__10396;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10374;
    wire N__10371;
    wire N__10370;
    wire N__10369;
    wire N__10366;
    wire N__10363;
    wire N__10362;
    wire N__10359;
    wire N__10354;
    wire N__10351;
    wire N__10344;
    wire N__10341;
    wire N__10338;
    wire N__10335;
    wire N__10332;
    wire N__10329;
    wire N__10326;
    wire N__10323;
    wire N__10320;
    wire N__10319;
    wire N__10314;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10306;
    wire N__10301;
    wire N__10298;
    wire N__10293;
    wire N__10290;
    wire N__10287;
    wire N__10284;
    wire N__10283;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10275;
    wire N__10272;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10230;
    wire N__10227;
    wire N__10224;
    wire N__10221;
    wire N__10218;
    wire N__10215;
    wire N__10212;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10200;
    wire N__10197;
    wire N__10196;
    wire N__10195;
    wire N__10194;
    wire N__10191;
    wire N__10188;
    wire N__10185;
    wire N__10182;
    wire N__10173;
    wire N__10170;
    wire N__10167;
    wire N__10166;
    wire N__10165;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10152;
    wire N__10149;
    wire N__10142;
    wire N__10137;
    wire N__10134;
    wire N__10131;
    wire N__10128;
    wire N__10125;
    wire N__10122;
    wire N__10119;
    wire N__10118;
    wire N__10115;
    wire N__10114;
    wire N__10111;
    wire N__10108;
    wire N__10105;
    wire N__10102;
    wire N__10097;
    wire N__10094;
    wire N__10093;
    wire N__10090;
    wire N__10087;
    wire N__10084;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10059;
    wire N__10056;
    wire N__10053;
    wire N__10050;
    wire N__10049;
    wire N__10048;
    wire N__10045;
    wire N__10044;
    wire N__10043;
    wire N__10042;
    wire N__10041;
    wire N__10040;
    wire N__10039;
    wire N__10036;
    wire N__10035;
    wire N__10034;
    wire N__10033;
    wire N__10032;
    wire N__10031;
    wire N__10028;
    wire N__10027;
    wire N__10026;
    wire N__10023;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10011;
    wire N__10008;
    wire N__10001;
    wire N__9994;
    wire N__9993;
    wire N__9992;
    wire N__9989;
    wire N__9984;
    wire N__9981;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9967;
    wire N__9964;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9945;
    wire N__9944;
    wire N__9939;
    wire N__9936;
    wire N__9933;
    wire N__9930;
    wire N__9923;
    wire N__9918;
    wire N__9915;
    wire N__9910;
    wire N__9907;
    wire N__9902;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9883;
    wire N__9880;
    wire N__9877;
    wire N__9874;
    wire N__9867;
    wire N__9864;
    wire N__9861;
    wire N__9858;
    wire N__9857;
    wire N__9856;
    wire N__9855;
    wire N__9854;
    wire N__9853;
    wire N__9852;
    wire N__9851;
    wire N__9834;
    wire N__9831;
    wire N__9828;
    wire N__9827;
    wire N__9826;
    wire N__9825;
    wire N__9824;
    wire N__9823;
    wire N__9822;
    wire N__9821;
    wire N__9820;
    wire N__9819;
    wire N__9818;
    wire N__9817;
    wire N__9816;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9780;
    wire N__9777;
    wire N__9774;
    wire N__9771;
    wire N__9768;
    wire N__9765;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9751;
    wire N__9750;
    wire N__9749;
    wire N__9744;
    wire N__9741;
    wire N__9738;
    wire N__9735;
    wire N__9734;
    wire N__9733;
    wire N__9730;
    wire N__9727;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9705;
    wire N__9702;
    wire N__9699;
    wire N__9696;
    wire N__9693;
    wire N__9684;
    wire N__9681;
    wire N__9678;
    wire N__9675;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9663;
    wire N__9660;
    wire N__9659;
    wire N__9658;
    wire N__9657;
    wire N__9656;
    wire N__9655;
    wire N__9654;
    wire N__9653;
    wire N__9652;
    wire N__9651;
    wire N__9650;
    wire N__9649;
    wire N__9648;
    wire N__9647;
    wire N__9646;
    wire N__9645;
    wire N__9644;
    wire N__9643;
    wire N__9642;
    wire N__9641;
    wire N__9640;
    wire N__9639;
    wire N__9638;
    wire N__9637;
    wire N__9636;
    wire N__9635;
    wire N__9634;
    wire N__9633;
    wire N__9632;
    wire N__9631;
    wire N__9630;
    wire N__9629;
    wire N__9626;
    wire N__9625;
    wire N__9624;
    wire N__9623;
    wire N__9622;
    wire N__9621;
    wire N__9620;
    wire N__9619;
    wire N__9618;
    wire N__9617;
    wire N__9616;
    wire N__9531;
    wire N__9528;
    wire N__9527;
    wire N__9522;
    wire N__9519;
    wire N__9516;
    wire N__9513;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9501;
    wire N__9498;
    wire N__9495;
    wire N__9492;
    wire N__9489;
    wire N__9486;
    wire N__9483;
    wire N__9480;
    wire N__9477;
    wire N__9474;
    wire N__9471;
    wire N__9468;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9458;
    wire N__9457;
    wire N__9454;
    wire N__9451;
    wire N__9448;
    wire N__9445;
    wire N__9444;
    wire N__9439;
    wire N__9436;
    wire N__9433;
    wire N__9430;
    wire N__9427;
    wire N__9424;
    wire N__9421;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9405;
    wire N__9402;
    wire N__9399;
    wire N__9396;
    wire N__9393;
    wire N__9392;
    wire N__9391;
    wire N__9390;
    wire N__9389;
    wire N__9388;
    wire N__9387;
    wire N__9384;
    wire N__9383;
    wire N__9380;
    wire N__9379;
    wire N__9378;
    wire N__9375;
    wire N__9372;
    wire N__9371;
    wire N__9370;
    wire N__9369;
    wire N__9366;
    wire N__9365;
    wire N__9360;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9346;
    wire N__9341;
    wire N__9340;
    wire N__9337;
    wire N__9332;
    wire N__9329;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9307;
    wire N__9306;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9294;
    wire N__9293;
    wire N__9290;
    wire N__9285;
    wire N__9282;
    wire N__9279;
    wire N__9274;
    wire N__9271;
    wire N__9266;
    wire N__9263;
    wire N__9258;
    wire N__9253;
    wire N__9246;
    wire N__9241;
    wire N__9236;
    wire N__9227;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9203;
    wire N__9202;
    wire N__9201;
    wire N__9200;
    wire N__9199;
    wire N__9196;
    wire N__9195;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9181;
    wire N__9180;
    wire N__9177;
    wire N__9176;
    wire N__9175;
    wire N__9174;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9154;
    wire N__9153;
    wire N__9150;
    wire N__9149;
    wire N__9144;
    wire N__9137;
    wire N__9136;
    wire N__9135;
    wire N__9130;
    wire N__9129;
    wire N__9128;
    wire N__9127;
    wire N__9122;
    wire N__9113;
    wire N__9108;
    wire N__9105;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9090;
    wire N__9087;
    wire N__9082;
    wire N__9079;
    wire N__9078;
    wire N__9075;
    wire N__9072;
    wire N__9069;
    wire N__9066;
    wire N__9063;
    wire N__9048;
    wire N__9045;
    wire N__9042;
    wire N__9037;
    wire N__9032;
    wire N__9029;
    wire N__9018;
    wire N__9015;
    wire N__9012;
    wire N__9009;
    wire N__9006;
    wire N__9003;
    wire N__9000;
    wire N__8997;
    wire N__8994;
    wire N__8991;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8955;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8943;
    wire N__8940;
    wire N__8939;
    wire N__8938;
    wire N__8937;
    wire N__8934;
    wire N__8929;
    wire N__8926;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8910;
    wire N__8909;
    wire N__8904;
    wire N__8901;
    wire N__8898;
    wire N__8895;
    wire N__8892;
    wire N__8889;
    wire N__8886;
    wire N__8883;
    wire N__8880;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8862;
    wire N__8859;
    wire N__8856;
    wire N__8853;
    wire N__8850;
    wire N__8849;
    wire N__8848;
    wire N__8847;
    wire N__8844;
    wire N__8843;
    wire N__8842;
    wire N__8835;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8823;
    wire N__8822;
    wire N__8817;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8793;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8777;
    wire N__8772;
    wire N__8771;
    wire N__8770;
    wire N__8769;
    wire N__8768;
    wire N__8767;
    wire N__8766;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8746;
    wire N__8741;
    wire N__8736;
    wire N__8733;
    wire N__8732;
    wire N__8729;
    wire N__8728;
    wire N__8725;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8704;
    wire N__8701;
    wire N__8698;
    wire N__8695;
    wire N__8690;
    wire N__8685;
    wire N__8684;
    wire N__8683;
    wire N__8682;
    wire N__8679;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8668;
    wire N__8665;
    wire N__8662;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8640;
    wire N__8639;
    wire N__8634;
    wire N__8629;
    wire N__8626;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8610;
    wire N__8607;
    wire N__8606;
    wire N__8605;
    wire N__8602;
    wire N__8599;
    wire N__8598;
    wire N__8597;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8587;
    wire N__8580;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8557;
    wire N__8552;
    wire N__8547;
    wire N__8544;
    wire N__8541;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8529;
    wire N__8526;
    wire N__8523;
    wire N__8520;
    wire N__8517;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8466;
    wire N__8465;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8457;
    wire N__8454;
    wire N__8451;
    wire N__8448;
    wire N__8445;
    wire N__8442;
    wire N__8439;
    wire N__8436;
    wire N__8433;
    wire N__8432;
    wire N__8429;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8406;
    wire N__8405;
    wire N__8404;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8390;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8373;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8328;
    wire N__8325;
    wire N__8322;
    wire N__8319;
    wire N__8316;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8304;
    wire N__8301;
    wire N__8298;
    wire N__8295;
    wire N__8292;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8282;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8269;
    wire N__8268;
    wire N__8267;
    wire N__8266;
    wire N__8263;
    wire N__8260;
    wire N__8255;
    wire N__8250;
    wire N__8241;
    wire N__8238;
    wire N__8237;
    wire N__8236;
    wire N__8235;
    wire N__8234;
    wire N__8231;
    wire N__8230;
    wire N__8227;
    wire N__8226;
    wire N__8223;
    wire N__8220;
    wire N__8219;
    wire N__8216;
    wire N__8213;
    wire N__8210;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8169;
    wire N__8166;
    wire N__8163;
    wire N__8160;
    wire N__8157;
    wire N__8154;
    wire N__8151;
    wire N__8148;
    wire N__8145;
    wire N__8144;
    wire N__8143;
    wire N__8140;
    wire N__8137;
    wire N__8134;
    wire N__8127;
    wire N__8124;
    wire N__8121;
    wire N__8118;
    wire N__8115;
    wire N__8112;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8097;
    wire N__8094;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8084;
    wire N__8083;
    wire N__8082;
    wire N__8081;
    wire N__8080;
    wire N__8077;
    wire N__8074;
    wire N__8073;
    wire N__8070;
    wire N__8067;
    wire N__8064;
    wire N__8061;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8036;
    wire N__8031;
    wire N__8026;
    wire N__8023;
    wire N__8016;
    wire N__8015;
    wire N__8010;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7977;
    wire N__7974;
    wire N__7971;
    wire N__7968;
    wire N__7965;
    wire N__7962;
    wire N__7959;
    wire N__7956;
    wire N__7953;
    wire N__7950;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7917;
    wire N__7914;
    wire N__7911;
    wire N__7908;
    wire N__7905;
    wire N__7902;
    wire N__7899;
    wire N__7896;
    wire N__7893;
    wire N__7890;
    wire N__7887;
    wire N__7884;
    wire N__7881;
    wire N__7878;
    wire N__7875;
    wire N__7872;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7851;
    wire N__7848;
    wire N__7845;
    wire N__7842;
    wire N__7839;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7819;
    wire N__7816;
    wire N__7813;
    wire N__7810;
    wire N__7803;
    wire N__7800;
    wire N__7797;
    wire N__7794;
    wire N__7791;
    wire N__7788;
    wire N__7785;
    wire N__7782;
    wire N__7781;
    wire N__7780;
    wire N__7779;
    wire N__7778;
    wire N__7777;
    wire N__7774;
    wire N__7771;
    wire N__7768;
    wire N__7765;
    wire N__7762;
    wire N__7759;
    wire N__7758;
    wire N__7757;
    wire N__7756;
    wire N__7755;
    wire N__7754;
    wire N__7753;
    wire N__7752;
    wire N__7751;
    wire N__7750;
    wire N__7749;
    wire N__7748;
    wire N__7747;
    wire N__7746;
    wire N__7745;
    wire N__7744;
    wire N__7743;
    wire N__7742;
    wire N__7741;
    wire N__7736;
    wire N__7729;
    wire N__7726;
    wire N__7721;
    wire N__7718;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7699;
    wire N__7696;
    wire N__7693;
    wire N__7684;
    wire N__7681;
    wire N__7678;
    wire N__7673;
    wire N__7660;
    wire N__7657;
    wire N__7654;
    wire N__7647;
    wire N__7646;
    wire N__7645;
    wire N__7644;
    wire N__7641;
    wire N__7638;
    wire N__7631;
    wire N__7626;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7610;
    wire N__7601;
    wire N__7598;
    wire N__7595;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7581;
    wire N__7578;
    wire N__7575;
    wire N__7572;
    wire N__7569;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7551;
    wire N__7548;
    wire N__7545;
    wire N__7542;
    wire N__7539;
    wire N__7536;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7485;
    wire N__7482;
    wire N__7479;
    wire N__7476;
    wire N__7473;
    wire N__7472;
    wire N__7471;
    wire N__7468;
    wire N__7465;
    wire N__7462;
    wire N__7459;
    wire N__7454;
    wire N__7449;
    wire N__7448;
    wire N__7445;
    wire N__7444;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7432;
    wire N__7427;
    wire N__7422;
    wire N__7421;
    wire N__7420;
    wire N__7419;
    wire N__7416;
    wire N__7413;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7405;
    wire N__7404;
    wire N__7399;
    wire N__7396;
    wire N__7393;
    wire N__7392;
    wire N__7389;
    wire N__7384;
    wire N__7379;
    wire N__7376;
    wire N__7373;
    wire N__7362;
    wire N__7359;
    wire N__7356;
    wire N__7353;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7341;
    wire N__7338;
    wire N__7335;
    wire N__7332;
    wire N__7329;
    wire N__7326;
    wire N__7323;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7311;
    wire N__7308;
    wire N__7305;
    wire N__7302;
    wire N__7299;
    wire N__7296;
    wire N__7293;
    wire N__7290;
    wire N__7287;
    wire N__7284;
    wire N__7281;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7273;
    wire N__7272;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7257;
    wire N__7248;
    wire N__7247;
    wire N__7246;
    wire N__7245;
    wire N__7242;
    wire N__7241;
    wire N__7238;
    wire N__7237;
    wire N__7236;
    wire N__7235;
    wire N__7230;
    wire N__7229;
    wire N__7226;
    wire N__7225;
    wire N__7224;
    wire N__7223;
    wire N__7218;
    wire N__7217;
    wire N__7216;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7191;
    wire N__7188;
    wire N__7183;
    wire N__7180;
    wire N__7161;
    wire N__7160;
    wire N__7159;
    wire N__7156;
    wire N__7155;
    wire N__7152;
    wire N__7149;
    wire N__7148;
    wire N__7147;
    wire N__7146;
    wire N__7145;
    wire N__7142;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7127;
    wire N__7124;
    wire N__7123;
    wire N__7122;
    wire N__7121;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7109;
    wire N__7102;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7074;
    wire N__7071;
    wire N__7068;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7058;
    wire N__7057;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7047;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7037;
    wire N__7036;
    wire N__7033;
    wire N__7030;
    wire N__7029;
    wire N__7024;
    wire N__7019;
    wire N__7014;
    wire N__7011;
    wire N__7002;
    wire N__6999;
    wire N__6998;
    wire N__6995;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6985;
    wire N__6984;
    wire N__6981;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6963;
    wire N__6962;
    wire N__6957;
    wire N__6954;
    wire N__6951;
    wire N__6948;
    wire N__6945;
    wire N__6942;
    wire N__6939;
    wire N__6936;
    wire N__6933;
    wire N__6930;
    wire N__6927;
    wire N__6924;
    wire N__6921;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6885;
    wire N__6882;
    wire N__6879;
    wire N__6876;
    wire N__6873;
    wire N__6870;
    wire N__6867;
    wire N__6866;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6856;
    wire N__6853;
    wire N__6850;
    wire N__6849;
    wire N__6846;
    wire N__6841;
    wire N__6838;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6815;
    wire N__6810;
    wire N__6807;
    wire N__6806;
    wire N__6805;
    wire N__6802;
    wire N__6799;
    wire N__6796;
    wire N__6793;
    wire N__6790;
    wire N__6787;
    wire N__6784;
    wire N__6781;
    wire N__6778;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6753;
    wire N__6750;
    wire N__6749;
    wire N__6748;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6740;
    wire N__6739;
    wire N__6738;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6726;
    wire N__6723;
    wire N__6720;
    wire N__6715;
    wire N__6702;
    wire N__6701;
    wire N__6700;
    wire N__6697;
    wire N__6694;
    wire N__6691;
    wire N__6684;
    wire N__6683;
    wire N__6680;
    wire N__6677;
    wire N__6676;
    wire N__6675;
    wire N__6674;
    wire N__6669;
    wire N__6664;
    wire N__6663;
    wire N__6662;
    wire N__6661;
    wire N__6658;
    wire N__6657;
    wire N__6656;
    wire N__6651;
    wire N__6650;
    wire N__6649;
    wire N__6646;
    wire N__6645;
    wire N__6642;
    wire N__6641;
    wire N__6636;
    wire N__6635;
    wire N__6634;
    wire N__6633;
    wire N__6630;
    wire N__6627;
    wire N__6624;
    wire N__6619;
    wire N__6616;
    wire N__6613;
    wire N__6608;
    wire N__6605;
    wire N__6600;
    wire N__6597;
    wire N__6576;
    wire N__6575;
    wire N__6574;
    wire N__6573;
    wire N__6572;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6564;
    wire N__6563;
    wire N__6562;
    wire N__6561;
    wire N__6558;
    wire N__6555;
    wire N__6554;
    wire N__6551;
    wire N__6550;
    wire N__6549;
    wire N__6542;
    wire N__6539;
    wire N__6538;
    wire N__6535;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6483;
    wire N__6480;
    wire N__6477;
    wire N__6474;
    wire N__6471;
    wire N__6468;
    wire N__6467;
    wire N__6462;
    wire N__6459;
    wire N__6456;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6441;
    wire N__6438;
    wire N__6435;
    wire N__6432;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6420;
    wire N__6417;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6375;
    wire N__6374;
    wire N__6371;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6357;
    wire N__6354;
    wire N__6351;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6336;
    wire N__6333;
    wire N__6330;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6315;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6303;
    wire N__6302;
    wire N__6299;
    wire N__6296;
    wire N__6291;
    wire N__6290;
    wire N__6287;
    wire N__6286;
    wire N__6283;
    wire N__6280;
    wire N__6277;
    wire N__6274;
    wire N__6267;
    wire N__6264;
    wire N__6261;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6251;
    wire N__6250;
    wire N__6247;
    wire N__6244;
    wire N__6241;
    wire N__6238;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6218;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6201;
    wire N__6200;
    wire N__6199;
    wire N__6196;
    wire N__6193;
    wire N__6190;
    wire N__6183;
    wire N__6180;
    wire N__6179;
    wire N__6178;
    wire N__6175;
    wire N__6172;
    wire N__6169;
    wire N__6162;
    wire N__6161;
    wire N__6158;
    wire N__6157;
    wire N__6156;
    wire N__6153;
    wire N__6150;
    wire N__6147;
    wire N__6146;
    wire N__6143;
    wire N__6138;
    wire N__6135;
    wire N__6134;
    wire N__6133;
    wire N__6130;
    wire N__6129;
    wire N__6128;
    wire N__6125;
    wire N__6120;
    wire N__6117;
    wire N__6114;
    wire N__6111;
    wire N__6106;
    wire N__6093;
    wire N__6090;
    wire N__6087;
    wire N__6086;
    wire N__6085;
    wire N__6082;
    wire N__6081;
    wire N__6080;
    wire N__6075;
    wire N__6072;
    wire N__6067;
    wire N__6060;
    wire N__6059;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6051;
    wire N__6050;
    wire N__6049;
    wire N__6048;
    wire N__6045;
    wire N__6040;
    wire N__6037;
    wire N__6036;
    wire N__6035;
    wire N__6032;
    wire N__6029;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6006;
    wire N__6003;
    wire N__5988;
    wire N__5985;
    wire N__5982;
    wire N__5979;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5967;
    wire N__5964;
    wire N__5961;
    wire N__5960;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5947;
    wire N__5940;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5930;
    wire N__5929;
    wire N__5928;
    wire N__5927;
    wire N__5926;
    wire N__5925;
    wire N__5924;
    wire N__5915;
    wire N__5910;
    wire N__5905;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5886;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5874;
    wire N__5871;
    wire N__5868;
    wire N__5865;
    wire N__5862;
    wire N__5859;
    wire N__5856;
    wire N__5853;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5829;
    wire N__5826;
    wire N__5823;
    wire N__5820;
    wire N__5817;
    wire N__5816;
    wire N__5815;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5802;
    wire N__5797;
    wire N__5794;
    wire N__5787;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5754;
    wire N__5751;
    wire N__5748;
    wire N__5745;
    wire N__5742;
    wire N__5739;
    wire N__5736;
    wire N__5735;
    wire N__5732;
    wire N__5731;
    wire N__5730;
    wire N__5727;
    wire N__5724;
    wire N__5723;
    wire N__5720;
    wire N__5717;
    wire N__5712;
    wire N__5709;
    wire N__5700;
    wire N__5697;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5685;
    wire N__5682;
    wire N__5679;
    wire N__5676;
    wire N__5673;
    wire N__5670;
    wire N__5669;
    wire N__5668;
    wire N__5667;
    wire N__5666;
    wire N__5665;
    wire N__5664;
    wire N__5663;
    wire N__5662;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5648;
    wire N__5647;
    wire N__5646;
    wire N__5645;
    wire N__5642;
    wire N__5637;
    wire N__5632;
    wire N__5629;
    wire N__5624;
    wire N__5617;
    wire N__5604;
    wire N__5601;
    wire N__5598;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5580;
    wire N__5577;
    wire N__5576;
    wire N__5575;
    wire N__5574;
    wire N__5571;
    wire N__5566;
    wire N__5563;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5532;
    wire N__5529;
    wire N__5528;
    wire N__5525;
    wire N__5524;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5512;
    wire N__5505;
    wire N__5502;
    wire N__5499;
    wire N__5496;
    wire N__5493;
    wire N__5490;
    wire N__5487;
    wire N__5484;
    wire N__5481;
    wire N__5478;
    wire N__5475;
    wire N__5474;
    wire N__5473;
    wire N__5472;
    wire N__5467;
    wire N__5462;
    wire N__5457;
    wire N__5456;
    wire N__5453;
    wire N__5450;
    wire N__5445;
    wire N__5444;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5434;
    wire N__5429;
    wire N__5424;
    wire N__5421;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5409;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5397;
    wire N__5394;
    wire N__5391;
    wire N__5388;
    wire N__5385;
    wire N__5382;
    wire N__5381;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5364;
    wire N__5361;
    wire N__5358;
    wire N__5355;
    wire N__5354;
    wire N__5353;
    wire N__5350;
    wire N__5345;
    wire N__5340;
    wire N__5339;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5310;
    wire N__5307;
    wire N__5304;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5292;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5280;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5265;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5253;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5241;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5229;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5217;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5205;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5187;
    wire N__5184;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5168;
    wire N__5165;
    wire N__5162;
    wire N__5157;
    wire N__5156;
    wire N__5155;
    wire N__5152;
    wire N__5151;
    wire N__5148;
    wire N__5145;
    wire N__5142;
    wire N__5139;
    wire N__5130;
    wire N__5127;
    wire N__5124;
    wire N__5121;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5070;
    wire N__5069;
    wire N__5068;
    wire N__5067;
    wire N__5066;
    wire N__5065;
    wire N__5064;
    wire N__5049;
    wire N__5046;
    wire N__5043;
    wire N__5040;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5010;
    wire N__5009;
    wire N__5008;
    wire N__5005;
    wire N__5004;
    wire N__4999;
    wire N__4996;
    wire N__4993;
    wire N__4990;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4902;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4881;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4854;
    wire N__4851;
    wire N__4848;
    wire N__4847;
    wire N__4846;
    wire N__4843;
    wire N__4838;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4743;
    wire N__4740;
    wire N__4737;
    wire N__4734;
    wire N__4733;
    wire N__4732;
    wire N__4731;
    wire N__4728;
    wire N__4727;
    wire N__4726;
    wire N__4725;
    wire N__4724;
    wire N__4723;
    wire N__4722;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4697;
    wire N__4688;
    wire N__4677;
    wire N__4674;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4593;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4575;
    wire N__4572;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4560;
    wire N__4559;
    wire N__4558;
    wire N__4555;
    wire N__4550;
    wire N__4545;
    wire N__4542;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4494;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4482;
    wire N__4479;
    wire N__4476;
    wire N__4473;
    wire N__4470;
    wire N__4467;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4431;
    wire N__4430;
    wire N__4429;
    wire N__4424;
    wire N__4421;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4401;
    wire N__4400;
    wire N__4399;
    wire N__4398;
    wire N__4397;
    wire N__4396;
    wire N__4393;
    wire N__4388;
    wire N__4385;
    wire N__4380;
    wire N__4371;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4322;
    wire N__4319;
    wire N__4318;
    wire N__4317;
    wire N__4316;
    wire N__4315;
    wire N__4314;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4299;
    wire N__4292;
    wire N__4281;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4245;
    wire N__4242;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4227;
    wire N__4226;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4212;
    wire N__4209;
    wire N__4208;
    wire N__4207;
    wire N__4204;
    wire N__4199;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4187;
    wire N__4186;
    wire N__4185;
    wire N__4184;
    wire N__4183;
    wire N__4180;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4158;
    wire N__4155;
    wire N__4154;
    wire N__4153;
    wire N__4152;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4119;
    wire N__4118;
    wire N__4117;
    wire N__4114;
    wire N__4113;
    wire N__4112;
    wire N__4109;
    wire N__4108;
    wire N__4105;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4091;
    wire N__4080;
    wire N__4077;
    wire N__4074;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4047;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4035;
    wire N__4032;
    wire N__4029;
    wire N__4026;
    wire N__4023;
    wire N__4020;
    wire N__4017;
    wire N__4014;
    wire N__4011;
    wire N__4008;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3987;
    wire N__3984;
    wire N__3981;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_PLL_i_i;
    wire N_812_i;
    wire TACK_EN_i_ess;
    wire DBRn_c_i_0;
    wire \U712_REG_SM.N_266_cascade_ ;
    wire \U712_REG_SM.N_269_cascade_ ;
    wire \U712_REG_SM.N_233 ;
    wire \U712_REG_SM.N_191_cascade_ ;
    wire C3_c;
    wire \U712_REG_SM.N_85 ;
    wire \U712_REG_SM.N_263 ;
    wire \U712_REG_SM.N_209 ;
    wire \U712_REG_SM.STATE_COUNTc_1_0_cascade_ ;
    wire \U712_REG_SM.N_272_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_1 ;
    wire \U712_REG_SM.STATE_COUNT_srsts_i_0_a5_0_0_0 ;
    wire \U712_REG_SM.N_207 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.N_191 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_0 ;
    wire \U712_REG_SM.DS_EN_RNOZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire DBRn_c;
    wire DBR_SYNCZ0Z_0;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire VBENn_c;
    wire \U712_CYCLE_TERM.TACK_STATEZ1Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a5_0_0_0 ;
    wire REGSPACEn_c;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_i_i_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_i_i_0_cascade_ ;
    wire \U712_CHIP_RAM.N_23 ;
    wire \U712_REG_SM.N_219 ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.N_261 ;
    wire \U712_BYTE_ENABLE.N_215_cascade_ ;
    wire N_167_i;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire ASn_c;
    wire \U712_REG_SM.N_219_0_0 ;
    wire A_c_6;
    wire A_c_13;
    wire DBDIR_c;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire TACK_OUTn;
    wire N_165_i;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_a5_0Z0Z_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0 ;
    wire RAMSPACEn_c;
    wire TSn_c;
    wire \U712_CHIP_RAM.N_279_cascade_ ;
    wire \U712_CHIP_RAM.N_187_cascade_ ;
    wire \U712_CHIP_RAM.N_316_cascade_ ;
    wire \U712_CHIP_RAM.N_316 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a5_1 ;
    wire \U712_CHIP_RAM.N_283_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ;
    wire \U712_CHIP_RAM.N_258 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_ ;
    wire N_235;
    wire RnW_c;
    wire AWEn_c;
    wire \U712_CHIP_RAM.N_222 ;
    wire \U712_BYTE_ENABLE.N_217 ;
    wire DMA_LATCH_EN_c;
    wire A_c_11;
    wire A_c_4;
    wire A_c_3;
    wire A_c_10;
    wire bfn_10_9_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire \U712_CHIP_RAM.REFRESH5lto1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH5lto2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.N_340 ;
    wire \U712_CHIP_RAM.N_340_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_ ;
    wire \U712_CHIP_RAM.N_97 ;
    wire LATCH_CLK_c;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.N_312 ;
    wire \U712_CHIP_RAM.N_206_cascade_ ;
    wire \U712_CHIP_RAM.N_329 ;
    wire \U712_CHIP_RAM.BANK0_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_323_cascade_ ;
    wire \U712_CHIP_RAM.N_374 ;
    wire \U712_CHIP_RAM.N_378 ;
    wire \U712_CHIP_RAM.N_184 ;
    wire \U712_CHIP_RAM.N_335_cascade_ ;
    wire \U712_CHIP_RAM.N_280 ;
    wire \U712_CHIP_RAM.N_284 ;
    wire \U712_CHIP_RAM.N_284_cascade_ ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_CHIP_RAM.N_218 ;
    wire \U712_CHIP_RAM.N_218_cascade_ ;
    wire \U712_CHIP_RAM.N_259 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a2_0_a5_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_i_a5_0_1_cascade_ ;
    wire \U712_CHIP_RAM.N_257_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_i_0 ;
    wire \U712_CHIP_RAM.N_338_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_284_2 ;
    wire \U712_CHIP_RAM.N_253 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.N_284_2_cascade_ ;
    wire \U712_CHIP_RAM.N_254 ;
    wire \U712_CHIP_RAM.N_322 ;
    wire \U712_CHIP_RAM.N_206 ;
    wire \U712_CHIP_RAM.N_338 ;
    wire \U712_CHIP_RAM.N_256 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire A_c_5;
    wire A_c_12;
    wire A_c_16;
    wire A_c_18;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.N_211_i_0_en_cascade_ ;
    wire \U712_CYCLE_TERM.N_211_i_0_en_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0 ;
    wire \U712_CHIP_RAM.N_339_cascade_ ;
    wire \U712_CHIP_RAM.N_335 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_1_cascade_ ;
    wire \U712_CHIP_RAM.N_296 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire bfn_11_12_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.N_181 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire A_c_20;
    wire \U712_CHIP_RAM.N_289_cascade_ ;
    wire \U712_CHIP_RAM.N_288 ;
    wire BANK0_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a5_0 ;
    wire \U712_CHIP_RAM.N_186 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0 ;
    wire \U712_CHIP_RAM.N_341 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ;
    wire \U712_CHIP_RAM.N_331 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.N_331_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ;
    wire \U712_CHIP_RAM.N_337 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.un3_DMA_CYCLE_START ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire CONSTANT_ONE_NET;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CMA_c_2;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire A_c_9;
    wire A_c_2;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire A_c_7;
    wire CLK40_PLL_i;
    wire CLK40_PLL_i_i;
    wire \U712_CHIP_RAM.N_327 ;
    wire \U712_CHIP_RAM.N_339 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire REG_TACK;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire WRITE_CYCLEm;
    wire CPU_TACKm;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0 ;
    wire N_118_i;
    wire N_119_i;
    wire \U712_CHIP_RAM.N_323 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.CPU_TACK_7_iv_i_a5_0_1_0 ;
    wire \U712_CHIP_RAM.N_287 ;
    wire DMA_CYCLEm;
    wire DBENn_c;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_a5_0Z0Z_0 ;
    wire \U712_BYTE_ENABLE.UUBE ;
    wire \U712_BYTE_ENABLE.N_216 ;
    wire RESETn_c;
    wire RESETn_c_i;
    wire N_163;
    wire A_c_17;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.N_146 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5_cascade_ ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire A_c_14;
    wire \U712_CHIP_RAM.CMA_5_0_8_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire \U712_CHIP_RAM.un1_CMA28_0_i ;
    wire A_c_15;
    wire A_c_8;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.CLK_EN_6_0_a5_2 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0 ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire DS_ENm;
    wire U712_BYTE_ENABLE_un1_UDSn_i;
    wire WEn_c;
    wire CASn_c;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire CPU_CYCLEm;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire U712_BYTE_ENABLE_UUBE_i;
    wire N_215_i;
    wire N_217_i;
    wire A_c_1;
    wire A_c_0;
    wire SIZ_c_0;
    wire SIZ_c_1;
    wire N_216_i;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire CLK80_PLL;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_AZ0Z20 ;
    wire \INVU712_CHIP_RAM.DMA_A20C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire DRA_c_5;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire DRA_c_4;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire DRA_c_7;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_9;
    wire RAS0n_c;
    wire AGNUS_REV_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire REG_CYCLEm;
    wire CASUn_c;
    wire CASLn_c;
    wire DRDENn_c;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__3939),
            .RESETB(N__6459),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__11659),
            .DIN(N__11658),
            .DOUT(N__11657),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__11659),
            .PADOUT(N__11658),
            .PADIN(N__11657),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7002),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11650),
            .DIN(N__11649),
            .DOUT(N__11648),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11650),
            .PADOUT(N__11649),
            .PADIN(N__11648),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__11641),
            .DIN(N__11640),
            .DOUT(N__11639),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__11641),
            .PADOUT(N__11640),
            .PADIN(N__11639),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8514),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__11632),
            .DIN(N__11631),
            .DOUT(N__11630),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__11632),
            .PADOUT(N__11631),
            .PADIN(N__11630),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5034),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__11623),
            .DIN(N__11622),
            .DOUT(N__11621),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__11623),
            .PADOUT(N__11622),
            .PADIN(N__11621),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__11614),
            .DIN(N__11613),
            .DOUT(N__11612),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__11614),
            .PADOUT(N__11613),
            .PADIN(N__11612),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__11605),
            .DIN(N__11604),
            .DOUT(N__11603),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__11605),
            .PADOUT(N__11604),
            .PADIN(N__11603),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__11596),
            .DIN(N__11595),
            .DOUT(N__11594),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__11596),
            .PADOUT(N__11595),
            .PADIN(N__11594),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__11587),
            .DIN(N__11586),
            .DOUT(N__11585),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__11587),
            .PADOUT(N__11586),
            .PADIN(N__11585),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11578),
            .DIN(N__11577),
            .DOUT(N__11576),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11578),
            .PADOUT(N__11577),
            .PADIN(N__11576),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__11569),
            .DIN(N__11568),
            .DOUT(N__11567),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__11569),
            .PADOUT(N__11568),
            .PADIN(N__11567),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7914),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__11560),
            .DIN(N__11559),
            .DOUT(N__11558),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__11560),
            .PADOUT(N__11559),
            .PADIN(N__11558),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8895),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__11551),
            .DIN(N__11550),
            .DOUT(N__11549),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__11551),
            .PADOUT(N__11550),
            .PADIN(N__11549),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__11542),
            .DIN(N__11541),
            .DOUT(N__11540),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__11542),
            .PADOUT(N__11541),
            .PADIN(N__11540),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__11533),
            .DIN(N__11532),
            .DOUT(N__11531),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__11533),
            .PADOUT(N__11532),
            .PADIN(N__11531),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__11524),
            .DIN(N__11523),
            .DOUT(N__11522),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__11524),
            .PADOUT(N__11523),
            .PADIN(N__11522),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4239),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__11515),
            .DIN(N__11514),
            .DOUT(N__11513),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__11515),
            .PADOUT(N__11514),
            .PADIN(N__11513),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11506),
            .DIN(N__11505),
            .DOUT(N__11504),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11506),
            .PADOUT(N__11505),
            .PADIN(N__11504),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__11497),
            .DIN(N__11496),
            .DOUT(N__11495),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__11497),
            .PADOUT(N__11496),
            .PADIN(N__11495),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7935),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__11488),
            .DIN(N__11487),
            .DOUT(N__11486),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__11488),
            .PADOUT(N__11487),
            .PADIN(N__11486),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__11479),
            .DIN(N__11478),
            .DOUT(N__11477),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__11479),
            .PADOUT(N__11478),
            .PADIN(N__11477),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8496),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11470),
            .DIN(N__11469),
            .DOUT(N__11468),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11470),
            .PADOUT(N__11469),
            .PADIN(N__11468),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__11461),
            .DIN(N__11460),
            .DOUT(N__11459),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__11461),
            .PADOUT(N__11460),
            .PADIN(N__11459),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8880),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__11452),
            .DIN(N__11451),
            .DOUT(N__11450),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__11452),
            .PADOUT(N__11451),
            .PADIN(N__11450),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11443),
            .DIN(N__11442),
            .DOUT(N__11441),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11443),
            .PADOUT(N__11442),
            .PADIN(N__11441),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__11434),
            .DIN(N__11433),
            .DOUT(N__11432),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__11434),
            .PADOUT(N__11433),
            .PADIN(N__11432),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11425),
            .DIN(N__11424),
            .DOUT(N__11423),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11425),
            .PADOUT(N__11424),
            .PADIN(N__11423),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__11416),
            .DIN(N__11415),
            .DOUT(N__11414),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__11416),
            .PADOUT(N__11415),
            .PADIN(N__11414),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__11407),
            .DIN(N__11406),
            .DOUT(N__11405),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__11407),
            .PADOUT(N__11406),
            .PADIN(N__11405),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4923),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__11398),
            .DIN(N__11397),
            .DOUT(N__11396),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__11398),
            .PADOUT(N__11397),
            .PADIN(N__11396),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11389),
            .DIN(N__11388),
            .DOUT(N__11387),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11389),
            .PADOUT(N__11388),
            .PADIN(N__11387),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11380),
            .DIN(N__11379),
            .DOUT(N__11378),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11380),
            .PADOUT(N__11379),
            .PADIN(N__11378),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11371),
            .DIN(N__11370),
            .DOUT(N__11369),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11371),
            .PADOUT(N__11370),
            .PADIN(N__11369),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__11362),
            .DIN(N__11361),
            .DOUT(N__11360),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__11362),
            .PADOUT(N__11361),
            .PADIN(N__11360),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6810),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__11353),
            .DIN(N__11352),
            .DOUT(N__11351),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__11353),
            .PADOUT(N__11352),
            .PADIN(N__11351),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__11344),
            .DIN(N__11343),
            .DOUT(N__11342),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__11344),
            .PADOUT(N__11343),
            .PADIN(N__11342),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9684),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__11335),
            .DIN(N__11334),
            .DOUT(N__11333),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__11335),
            .PADOUT(N__11334),
            .PADIN(N__11333),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__11326),
            .DIN(N__11325),
            .DOUT(N__11324),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__11326),
            .PADOUT(N__11325),
            .PADIN(N__11324),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6327),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__11317),
            .DIN(N__11316),
            .DOUT(N__11315),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__11317),
            .PADOUT(N__11316),
            .PADIN(N__11315),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6806),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11308),
            .DIN(N__11307),
            .DOUT(N__11306),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11308),
            .PADOUT(N__11307),
            .PADIN(N__11306),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3954),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__11299),
            .DIN(N__11298),
            .DOUT(N__11297),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__11299),
            .PADOUT(N__11298),
            .PADIN(N__11297),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__11290),
            .DIN(N__11289),
            .DOUT(N__11288),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__11290),
            .PADOUT(N__11289),
            .PADIN(N__11288),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4677),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11281),
            .DIN(N__11280),
            .DOUT(N__11279),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11281),
            .PADOUT(N__11280),
            .PADIN(N__11279),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6399),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11272),
            .DIN(N__11271),
            .DOUT(N__11270),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11272),
            .PADOUT(N__11271),
            .PADIN(N__11270),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11263),
            .DIN(N__11262),
            .DOUT(N__11261),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11263),
            .PADOUT(N__11262),
            .PADIN(N__11261),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11254),
            .DIN(N__11253),
            .DOUT(N__11252),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11254),
            .PADOUT(N__11253),
            .PADIN(N__11252),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__11245),
            .DIN(N__11244),
            .DOUT(N__11243),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__11245),
            .PADOUT(N__11244),
            .PADIN(N__11243),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__11236),
            .DIN(N__11235),
            .DOUT(N__11234),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__11236),
            .PADOUT(N__11235),
            .PADIN(N__11234),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8328),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11227),
            .DIN(N__11226),
            .DOUT(N__11225),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11227),
            .PADOUT(N__11226),
            .PADIN(N__11225),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11218),
            .DIN(N__11217),
            .DOUT(N__11216),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11218),
            .PADOUT(N__11217),
            .PADIN(N__11216),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6805),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__11209),
            .DIN(N__11208),
            .DOUT(N__11207),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__11209),
            .PADOUT(N__11208),
            .PADIN(N__11207),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8304),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11200),
            .DIN(N__11199),
            .DOUT(N__11198),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11200),
            .PADOUT(N__11199),
            .PADIN(N__11198),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10476),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11191),
            .DIN(N__11190),
            .DOUT(N__11189),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11191),
            .PADOUT(N__11190),
            .PADIN(N__11189),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4746),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11182),
            .DIN(N__11181),
            .DOUT(N__11180),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11182),
            .PADOUT(N__11181),
            .PADIN(N__11180),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8106),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__11173),
            .DIN(N__11172),
            .DOUT(N__11171),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__11173),
            .PADOUT(N__11172),
            .PADIN(N__11171),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4673),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11164),
            .DIN(N__11163),
            .DOUT(N__11162),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11164),
            .PADOUT(N__11163),
            .PADIN(N__11162),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__11155),
            .DIN(N__11154),
            .DOUT(N__11153),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__11155),
            .PADOUT(N__11154),
            .PADIN(N__11153),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__11146),
            .DIN(N__11145),
            .DOUT(N__11144),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__11146),
            .PADOUT(N__11145),
            .PADIN(N__11144),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4521),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__11137),
            .DIN(N__11136),
            .DOUT(N__11135),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__11137),
            .PADOUT(N__11136),
            .PADIN(N__11135),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8535),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__11128),
            .DIN(N__11127),
            .DOUT(N__11126),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__11128),
            .PADOUT(N__11127),
            .PADIN(N__11126),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4587),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__11119),
            .DIN(N__11118),
            .DOUT(N__11117),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__11119),
            .PADOUT(N__11118),
            .PADIN(N__11117),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7308),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__11110),
            .DIN(N__11109),
            .DOUT(N__11108),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__11110),
            .PADOUT(N__11109),
            .PADIN(N__11108),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__11101),
            .DIN(N__11100),
            .DOUT(N__11099),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__11101),
            .PADOUT(N__11100),
            .PADIN(N__11099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11092),
            .DIN(N__11091),
            .DOUT(N__11090),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11092),
            .PADOUT(N__11091),
            .PADIN(N__11090),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11083),
            .DIN(N__11082),
            .DOUT(N__11081),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11083),
            .PADOUT(N__11082),
            .PADIN(N__11081),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__11074),
            .DIN(N__11073),
            .DOUT(N__11072),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__11074),
            .PADOUT(N__11073),
            .PADIN(N__11072),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6435),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__11065),
            .DIN(N__11064),
            .DOUT(N__11063),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__11065),
            .PADOUT(N__11064),
            .PADIN(N__11063),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8865),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__11056),
            .DIN(N__11055),
            .DOUT(N__11054),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__11056),
            .PADOUT(N__11055),
            .PADIN(N__11054),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__11047),
            .DIN(N__11046),
            .DOUT(N__11045),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__11047),
            .PADOUT(N__11046),
            .PADIN(N__11045),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7332),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__11038),
            .DIN(N__11037),
            .DOUT(N__11036),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__11038),
            .PADOUT(N__11037),
            .PADIN(N__11036),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4014),
            .DIN0(),
            .DOUT0(N__4545),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__11029),
            .DIN(N__11028),
            .DOUT(N__11027),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__11029),
            .PADOUT(N__11028),
            .PADIN(N__11027),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6417),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__11020),
            .DIN(N__11019),
            .DOUT(N__11018),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__11020),
            .PADOUT(N__11019),
            .PADIN(N__11018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__11011),
            .DIN(N__11010),
            .DOUT(N__11009),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__11011),
            .PADOUT(N__11010),
            .PADIN(N__11009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__11002),
            .DIN(N__11001),
            .DOUT(N__11000),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__11002),
            .PADOUT(N__11001),
            .PADIN(N__11000),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7542),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__10993),
            .DIN(N__10992),
            .DOUT(N__10991),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__10993),
            .PADOUT(N__10992),
            .PADIN(N__10991),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__10984),
            .DIN(N__10983),
            .DOUT(N__10982),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__10984),
            .PADOUT(N__10983),
            .PADIN(N__10982),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__10975),
            .DIN(N__10974),
            .DOUT(N__10973),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__10975),
            .PADOUT(N__10974),
            .PADIN(N__10973),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__10966),
            .DIN(N__10965),
            .DOUT(N__10964),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__10966),
            .PADOUT(N__10965),
            .PADIN(N__10964),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__10957),
            .DIN(N__10956),
            .DOUT(N__10955),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__10957),
            .PADOUT(N__10956),
            .PADIN(N__10955),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7500),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__10948),
            .DIN(N__10947),
            .DOUT(N__10946),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__10948),
            .PADOUT(N__10947),
            .PADIN(N__10946),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7803),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__10939),
            .DIN(N__10938),
            .DOUT(N__10937),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__10939),
            .PADOUT(N__10938),
            .PADIN(N__10937),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9783),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__10930),
            .DIN(N__10929),
            .DOUT(N__10928),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__10930),
            .PADOUT(N__10929),
            .PADIN(N__10928),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7881),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__10921),
            .DIN(N__10920),
            .DOUT(N__10919),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__10921),
            .PADOUT(N__10920),
            .PADIN(N__10919),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__10912),
            .DIN(N__10911),
            .DOUT(N__10910),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__10912),
            .PADOUT(N__10911),
            .PADIN(N__10910),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__10903),
            .DIN(N__10902),
            .DOUT(N__10901),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__10903),
            .PADOUT(N__10902),
            .PADIN(N__10901),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8169),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__10894),
            .DIN(N__10893),
            .DOUT(N__10892),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__10894),
            .PADOUT(N__10893),
            .PADIN(N__10892),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__10885),
            .DIN(N__10884),
            .DOUT(N__10883),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__10885),
            .PADOUT(N__10884),
            .PADIN(N__10883),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__10876),
            .DIN(N__10875),
            .DOUT(N__10874),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__10876),
            .PADOUT(N__10875),
            .PADIN(N__10874),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5178),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__10867),
            .DIN(N__10866),
            .DOUT(N__10865),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__10867),
            .PADOUT(N__10866),
            .PADIN(N__10865),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7578),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2647 (
            .O(N__10848),
            .I(N__10839));
    InMux I__2646 (
            .O(N__10847),
            .I(N__10836));
    InMux I__2645 (
            .O(N__10846),
            .I(N__10833));
    InMux I__2644 (
            .O(N__10845),
            .I(N__10830));
    InMux I__2643 (
            .O(N__10844),
            .I(N__10823));
    InMux I__2642 (
            .O(N__10843),
            .I(N__10823));
    InMux I__2641 (
            .O(N__10842),
            .I(N__10823));
    LocalMux I__2640 (
            .O(N__10839),
            .I(N__10809));
    LocalMux I__2639 (
            .O(N__10836),
            .I(N__10795));
    LocalMux I__2638 (
            .O(N__10833),
            .I(N__10792));
    LocalMux I__2637 (
            .O(N__10830),
            .I(N__10780));
    LocalMux I__2636 (
            .O(N__10823),
            .I(N__10777));
    SRMux I__2635 (
            .O(N__10822),
            .I(N__10680));
    SRMux I__2634 (
            .O(N__10821),
            .I(N__10680));
    SRMux I__2633 (
            .O(N__10820),
            .I(N__10680));
    SRMux I__2632 (
            .O(N__10819),
            .I(N__10680));
    SRMux I__2631 (
            .O(N__10818),
            .I(N__10680));
    SRMux I__2630 (
            .O(N__10817),
            .I(N__10680));
    SRMux I__2629 (
            .O(N__10816),
            .I(N__10680));
    SRMux I__2628 (
            .O(N__10815),
            .I(N__10680));
    SRMux I__2627 (
            .O(N__10814),
            .I(N__10680));
    SRMux I__2626 (
            .O(N__10813),
            .I(N__10680));
    SRMux I__2625 (
            .O(N__10812),
            .I(N__10680));
    Glb2LocalMux I__2624 (
            .O(N__10809),
            .I(N__10680));
    SRMux I__2623 (
            .O(N__10808),
            .I(N__10680));
    SRMux I__2622 (
            .O(N__10807),
            .I(N__10680));
    SRMux I__2621 (
            .O(N__10806),
            .I(N__10680));
    SRMux I__2620 (
            .O(N__10805),
            .I(N__10680));
    SRMux I__2619 (
            .O(N__10804),
            .I(N__10680));
    SRMux I__2618 (
            .O(N__10803),
            .I(N__10680));
    SRMux I__2617 (
            .O(N__10802),
            .I(N__10680));
    SRMux I__2616 (
            .O(N__10801),
            .I(N__10680));
    SRMux I__2615 (
            .O(N__10800),
            .I(N__10680));
    SRMux I__2614 (
            .O(N__10799),
            .I(N__10680));
    SRMux I__2613 (
            .O(N__10798),
            .I(N__10680));
    Glb2LocalMux I__2612 (
            .O(N__10795),
            .I(N__10680));
    Glb2LocalMux I__2611 (
            .O(N__10792),
            .I(N__10680));
    SRMux I__2610 (
            .O(N__10791),
            .I(N__10680));
    SRMux I__2609 (
            .O(N__10790),
            .I(N__10680));
    SRMux I__2608 (
            .O(N__10789),
            .I(N__10680));
    SRMux I__2607 (
            .O(N__10788),
            .I(N__10680));
    SRMux I__2606 (
            .O(N__10787),
            .I(N__10680));
    SRMux I__2605 (
            .O(N__10786),
            .I(N__10680));
    SRMux I__2604 (
            .O(N__10785),
            .I(N__10680));
    SRMux I__2603 (
            .O(N__10784),
            .I(N__10680));
    SRMux I__2602 (
            .O(N__10783),
            .I(N__10680));
    Glb2LocalMux I__2601 (
            .O(N__10780),
            .I(N__10680));
    Glb2LocalMux I__2600 (
            .O(N__10777),
            .I(N__10680));
    SRMux I__2599 (
            .O(N__10776),
            .I(N__10680));
    SRMux I__2598 (
            .O(N__10775),
            .I(N__10680));
    SRMux I__2597 (
            .O(N__10774),
            .I(N__10680));
    SRMux I__2596 (
            .O(N__10773),
            .I(N__10680));
    SRMux I__2595 (
            .O(N__10772),
            .I(N__10680));
    SRMux I__2594 (
            .O(N__10771),
            .I(N__10680));
    SRMux I__2593 (
            .O(N__10770),
            .I(N__10680));
    SRMux I__2592 (
            .O(N__10769),
            .I(N__10680));
    GlobalMux I__2591 (
            .O(N__10680),
            .I(N__10677));
    gio2CtrlBuf I__2590 (
            .O(N__10677),
            .I(RESETn_c_i_g));
    InMux I__2589 (
            .O(N__10674),
            .I(N__10670));
    InMux I__2588 (
            .O(N__10673),
            .I(N__10667));
    LocalMux I__2587 (
            .O(N__10670),
            .I(N__10663));
    LocalMux I__2586 (
            .O(N__10667),
            .I(N__10660));
    InMux I__2585 (
            .O(N__10666),
            .I(N__10657));
    Span12Mux_v I__2584 (
            .O(N__10663),
            .I(N__10654));
    Span4Mux_h I__2583 (
            .O(N__10660),
            .I(N__10650));
    LocalMux I__2582 (
            .O(N__10657),
            .I(N__10647));
    Span12Mux_h I__2581 (
            .O(N__10654),
            .I(N__10644));
    InMux I__2580 (
            .O(N__10653),
            .I(N__10641));
    Span4Mux_v I__2579 (
            .O(N__10650),
            .I(N__10636));
    Span4Mux_h I__2578 (
            .O(N__10647),
            .I(N__10636));
    Odrv12 I__2577 (
            .O(N__10644),
            .I(REG_CYCLEm));
    LocalMux I__2576 (
            .O(N__10641),
            .I(REG_CYCLEm));
    Odrv4 I__2575 (
            .O(N__10636),
            .I(REG_CYCLEm));
    InMux I__2574 (
            .O(N__10629),
            .I(N__10625));
    CascadeMux I__2573 (
            .O(N__10628),
            .I(N__10621));
    LocalMux I__2572 (
            .O(N__10625),
            .I(N__10617));
    InMux I__2571 (
            .O(N__10624),
            .I(N__10614));
    InMux I__2570 (
            .O(N__10621),
            .I(N__10611));
    CascadeMux I__2569 (
            .O(N__10620),
            .I(N__10608));
    Span4Mux_v I__2568 (
            .O(N__10617),
            .I(N__10603));
    LocalMux I__2567 (
            .O(N__10614),
            .I(N__10603));
    LocalMux I__2566 (
            .O(N__10611),
            .I(N__10600));
    InMux I__2565 (
            .O(N__10608),
            .I(N__10597));
    Span4Mux_v I__2564 (
            .O(N__10603),
            .I(N__10593));
    Span4Mux_v I__2563 (
            .O(N__10600),
            .I(N__10588));
    LocalMux I__2562 (
            .O(N__10597),
            .I(N__10588));
    InMux I__2561 (
            .O(N__10596),
            .I(N__10585));
    Span4Mux_h I__2560 (
            .O(N__10593),
            .I(N__10582));
    Span4Mux_v I__2559 (
            .O(N__10588),
            .I(N__10576));
    LocalMux I__2558 (
            .O(N__10585),
            .I(N__10576));
    Span4Mux_h I__2557 (
            .O(N__10582),
            .I(N__10573));
    InMux I__2556 (
            .O(N__10581),
            .I(N__10570));
    Sp12to4 I__2555 (
            .O(N__10576),
            .I(N__10567));
    Span4Mux_h I__2554 (
            .O(N__10573),
            .I(N__10562));
    LocalMux I__2553 (
            .O(N__10570),
            .I(N__10562));
    Span12Mux_v I__2552 (
            .O(N__10567),
            .I(N__10559));
    Span4Mux_h I__2551 (
            .O(N__10562),
            .I(N__10556));
    Span12Mux_h I__2550 (
            .O(N__10559),
            .I(N__10553));
    Span4Mux_v I__2549 (
            .O(N__10556),
            .I(N__10550));
    Odrv12 I__2548 (
            .O(N__10553),
            .I(CASUn_c));
    Odrv4 I__2547 (
            .O(N__10550),
            .I(CASUn_c));
    CascadeMux I__2546 (
            .O(N__10545),
            .I(N__10540));
    InMux I__2545 (
            .O(N__10544),
            .I(N__10537));
    InMux I__2544 (
            .O(N__10543),
            .I(N__10534));
    InMux I__2543 (
            .O(N__10540),
            .I(N__10531));
    LocalMux I__2542 (
            .O(N__10537),
            .I(N__10525));
    LocalMux I__2541 (
            .O(N__10534),
            .I(N__10525));
    LocalMux I__2540 (
            .O(N__10531),
            .I(N__10522));
    InMux I__2539 (
            .O(N__10530),
            .I(N__10519));
    Span4Mux_v I__2538 (
            .O(N__10525),
            .I(N__10511));
    Span4Mux_v I__2537 (
            .O(N__10522),
            .I(N__10511));
    LocalMux I__2536 (
            .O(N__10519),
            .I(N__10511));
    InMux I__2535 (
            .O(N__10518),
            .I(N__10508));
    Span4Mux_h I__2534 (
            .O(N__10511),
            .I(N__10503));
    LocalMux I__2533 (
            .O(N__10508),
            .I(N__10503));
    Span4Mux_v I__2532 (
            .O(N__10503),
            .I(N__10500));
    Span4Mux_v I__2531 (
            .O(N__10500),
            .I(N__10496));
    InMux I__2530 (
            .O(N__10499),
            .I(N__10493));
    Sp12to4 I__2529 (
            .O(N__10496),
            .I(N__10490));
    LocalMux I__2528 (
            .O(N__10493),
            .I(N__10487));
    Span12Mux_h I__2527 (
            .O(N__10490),
            .I(N__10484));
    Span12Mux_v I__2526 (
            .O(N__10487),
            .I(N__10481));
    Odrv12 I__2525 (
            .O(N__10484),
            .I(CASLn_c));
    Odrv12 I__2524 (
            .O(N__10481),
            .I(CASLn_c));
    IoInMux I__2523 (
            .O(N__10476),
            .I(N__10473));
    LocalMux I__2522 (
            .O(N__10473),
            .I(N__10470));
    Span12Mux_s7_v I__2521 (
            .O(N__10470),
            .I(N__10467));
    Odrv12 I__2520 (
            .O(N__10467),
            .I(DRDENn_c));
    InMux I__2519 (
            .O(N__10464),
            .I(N__10461));
    LocalMux I__2518 (
            .O(N__10461),
            .I(N__10457));
    InMux I__2517 (
            .O(N__10460),
            .I(N__10454));
    Span12Mux_h I__2516 (
            .O(N__10457),
            .I(N__10451));
    LocalMux I__2515 (
            .O(N__10454),
            .I(N__10448));
    Odrv12 I__2514 (
            .O(N__10451),
            .I(DBRn_c_i));
    Odrv4 I__2513 (
            .O(N__10448),
            .I(DBRn_c_i));
    InMux I__2512 (
            .O(N__10443),
            .I(N__10439));
    InMux I__2511 (
            .O(N__10442),
            .I(N__10436));
    LocalMux I__2510 (
            .O(N__10439),
            .I(N__10433));
    LocalMux I__2509 (
            .O(N__10436),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    Odrv12 I__2508 (
            .O(N__10433),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    InMux I__2507 (
            .O(N__10428),
            .I(N__10425));
    LocalMux I__2506 (
            .O(N__10425),
            .I(N__10422));
    Span4Mux_v I__2505 (
            .O(N__10422),
            .I(N__10419));
    Odrv4 I__2504 (
            .O(N__10419),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2503 (
            .O(N__10416),
            .I(N__10409));
    InMux I__2502 (
            .O(N__10415),
            .I(N__10409));
    InMux I__2501 (
            .O(N__10414),
            .I(N__10405));
    LocalMux I__2500 (
            .O(N__10409),
            .I(N__10402));
    InMux I__2499 (
            .O(N__10408),
            .I(N__10399));
    LocalMux I__2498 (
            .O(N__10405),
            .I(N__10396));
    Span4Mux_v I__2497 (
            .O(N__10402),
            .I(N__10391));
    LocalMux I__2496 (
            .O(N__10399),
            .I(N__10391));
    Span4Mux_v I__2495 (
            .O(N__10396),
            .I(N__10388));
    Span4Mux_h I__2494 (
            .O(N__10391),
            .I(N__10385));
    Span4Mux_v I__2493 (
            .O(N__10388),
            .I(N__10382));
    Span4Mux_v I__2492 (
            .O(N__10385),
            .I(N__10379));
    Sp12to4 I__2491 (
            .O(N__10382),
            .I(N__10374));
    Sp12to4 I__2490 (
            .O(N__10379),
            .I(N__10374));
    Odrv12 I__2489 (
            .O(N__10374),
            .I(DRA_c_5));
    InMux I__2488 (
            .O(N__10371),
            .I(N__10366));
    InMux I__2487 (
            .O(N__10370),
            .I(N__10363));
    InMux I__2486 (
            .O(N__10369),
            .I(N__10359));
    LocalMux I__2485 (
            .O(N__10366),
            .I(N__10354));
    LocalMux I__2484 (
            .O(N__10363),
            .I(N__10354));
    InMux I__2483 (
            .O(N__10362),
            .I(N__10351));
    LocalMux I__2482 (
            .O(N__10359),
            .I(N__10344));
    Span4Mux_v I__2481 (
            .O(N__10354),
            .I(N__10344));
    LocalMux I__2480 (
            .O(N__10351),
            .I(N__10344));
    Span4Mux_h I__2479 (
            .O(N__10344),
            .I(N__10341));
    Span4Mux_v I__2478 (
            .O(N__10341),
            .I(N__10338));
    Sp12to4 I__2477 (
            .O(N__10338),
            .I(N__10335));
    Odrv12 I__2476 (
            .O(N__10335),
            .I(DRA_c_6));
    InMux I__2475 (
            .O(N__10332),
            .I(N__10329));
    LocalMux I__2474 (
            .O(N__10329),
            .I(N__10326));
    Span4Mux_h I__2473 (
            .O(N__10326),
            .I(N__10323));
    Odrv4 I__2472 (
            .O(N__10323),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2471 (
            .O(N__10320),
            .I(N__10314));
    InMux I__2470 (
            .O(N__10319),
            .I(N__10314));
    LocalMux I__2469 (
            .O(N__10314),
            .I(N__10310));
    InMux I__2468 (
            .O(N__10313),
            .I(N__10307));
    Span4Mux_h I__2467 (
            .O(N__10310),
            .I(N__10301));
    LocalMux I__2466 (
            .O(N__10307),
            .I(N__10301));
    InMux I__2465 (
            .O(N__10306),
            .I(N__10298));
    Sp12to4 I__2464 (
            .O(N__10301),
            .I(N__10293));
    LocalMux I__2463 (
            .O(N__10298),
            .I(N__10293));
    Span12Mux_v I__2462 (
            .O(N__10293),
            .I(N__10290));
    Span12Mux_h I__2461 (
            .O(N__10290),
            .I(N__10287));
    Odrv12 I__2460 (
            .O(N__10287),
            .I(DRA_c_4));
    InMux I__2459 (
            .O(N__10284),
            .I(N__10279));
    InMux I__2458 (
            .O(N__10283),
            .I(N__10276));
    InMux I__2457 (
            .O(N__10282),
            .I(N__10272));
    LocalMux I__2456 (
            .O(N__10279),
            .I(N__10267));
    LocalMux I__2455 (
            .O(N__10276),
            .I(N__10267));
    InMux I__2454 (
            .O(N__10275),
            .I(N__10264));
    LocalMux I__2453 (
            .O(N__10272),
            .I(N__10261));
    Span4Mux_v I__2452 (
            .O(N__10267),
            .I(N__10256));
    LocalMux I__2451 (
            .O(N__10264),
            .I(N__10256));
    Span4Mux_v I__2450 (
            .O(N__10261),
            .I(N__10253));
    Span4Mux_h I__2449 (
            .O(N__10256),
            .I(N__10250));
    Span4Mux_v I__2448 (
            .O(N__10253),
            .I(N__10247));
    Span4Mux_v I__2447 (
            .O(N__10250),
            .I(N__10244));
    Sp12to4 I__2446 (
            .O(N__10247),
            .I(N__10239));
    Sp12to4 I__2445 (
            .O(N__10244),
            .I(N__10239));
    Odrv12 I__2444 (
            .O(N__10239),
            .I(DRA_c_3));
    InMux I__2443 (
            .O(N__10236),
            .I(N__10233));
    LocalMux I__2442 (
            .O(N__10233),
            .I(N__10230));
    Span4Mux_h I__2441 (
            .O(N__10230),
            .I(N__10227));
    Span4Mux_h I__2440 (
            .O(N__10227),
            .I(N__10224));
    Odrv4 I__2439 (
            .O(N__10224),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2438 (
            .O(N__10221),
            .I(N__10218));
    LocalMux I__2437 (
            .O(N__10218),
            .I(N__10215));
    Span4Mux_h I__2436 (
            .O(N__10215),
            .I(N__10212));
    Odrv4 I__2435 (
            .O(N__10212),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2434 (
            .O(N__10209),
            .I(N__10206));
    LocalMux I__2433 (
            .O(N__10206),
            .I(N__10203));
    Span4Mux_h I__2432 (
            .O(N__10203),
            .I(N__10200));
    Odrv4 I__2431 (
            .O(N__10200),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__2430 (
            .O(N__10197),
            .I(N__10191));
    InMux I__2429 (
            .O(N__10196),
            .I(N__10188));
    InMux I__2428 (
            .O(N__10195),
            .I(N__10185));
    InMux I__2427 (
            .O(N__10194),
            .I(N__10182));
    LocalMux I__2426 (
            .O(N__10191),
            .I(N__10173));
    LocalMux I__2425 (
            .O(N__10188),
            .I(N__10173));
    LocalMux I__2424 (
            .O(N__10185),
            .I(N__10173));
    LocalMux I__2423 (
            .O(N__10182),
            .I(N__10173));
    Span12Mux_h I__2422 (
            .O(N__10173),
            .I(N__10170));
    Odrv12 I__2421 (
            .O(N__10170),
            .I(DRA_c_7));
    InMux I__2420 (
            .O(N__10167),
            .I(N__10161));
    InMux I__2419 (
            .O(N__10166),
            .I(N__10158));
    InMux I__2418 (
            .O(N__10165),
            .I(N__10155));
    InMux I__2417 (
            .O(N__10164),
            .I(N__10152));
    LocalMux I__2416 (
            .O(N__10161),
            .I(N__10149));
    LocalMux I__2415 (
            .O(N__10158),
            .I(N__10142));
    LocalMux I__2414 (
            .O(N__10155),
            .I(N__10142));
    LocalMux I__2413 (
            .O(N__10152),
            .I(N__10142));
    Span4Mux_v I__2412 (
            .O(N__10149),
            .I(N__10137));
    Span4Mux_v I__2411 (
            .O(N__10142),
            .I(N__10137));
    Sp12to4 I__2410 (
            .O(N__10137),
            .I(N__10134));
    Odrv12 I__2409 (
            .O(N__10134),
            .I(DRA_c_8));
    CascadeMux I__2408 (
            .O(N__10131),
            .I(N__10128));
    InMux I__2407 (
            .O(N__10128),
            .I(N__10125));
    LocalMux I__2406 (
            .O(N__10125),
            .I(N__10122));
    Odrv12 I__2405 (
            .O(N__10122),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2404 (
            .O(N__10119),
            .I(N__10115));
    CascadeMux I__2403 (
            .O(N__10118),
            .I(N__10111));
    LocalMux I__2402 (
            .O(N__10115),
            .I(N__10108));
    InMux I__2401 (
            .O(N__10114),
            .I(N__10105));
    InMux I__2400 (
            .O(N__10111),
            .I(N__10102));
    Span4Mux_h I__2399 (
            .O(N__10108),
            .I(N__10097));
    LocalMux I__2398 (
            .O(N__10105),
            .I(N__10097));
    LocalMux I__2397 (
            .O(N__10102),
            .I(N__10094));
    Span4Mux_v I__2396 (
            .O(N__10097),
            .I(N__10090));
    Span4Mux_v I__2395 (
            .O(N__10094),
            .I(N__10087));
    InMux I__2394 (
            .O(N__10093),
            .I(N__10084));
    Sp12to4 I__2393 (
            .O(N__10090),
            .I(N__10079));
    Sp12to4 I__2392 (
            .O(N__10087),
            .I(N__10079));
    LocalMux I__2391 (
            .O(N__10084),
            .I(N__10076));
    Span12Mux_h I__2390 (
            .O(N__10079),
            .I(N__10073));
    Span12Mux_v I__2389 (
            .O(N__10076),
            .I(N__10070));
    Span12Mux_v I__2388 (
            .O(N__10073),
            .I(N__10067));
    Span12Mux_v I__2387 (
            .O(N__10070),
            .I(N__10064));
    Odrv12 I__2386 (
            .O(N__10067),
            .I(DRA_c_9));
    Odrv12 I__2385 (
            .O(N__10064),
            .I(DRA_c_9));
    InMux I__2384 (
            .O(N__10059),
            .I(N__10056));
    LocalMux I__2383 (
            .O(N__10056),
            .I(N__10053));
    Odrv12 I__2382 (
            .O(N__10053),
            .I(RAS0n_c));
    InMux I__2381 (
            .O(N__10050),
            .I(N__10045));
    CascadeMux I__2380 (
            .O(N__10049),
            .I(N__10036));
    CascadeMux I__2379 (
            .O(N__10048),
            .I(N__10028));
    LocalMux I__2378 (
            .O(N__10045),
            .I(N__10023));
    InMux I__2377 (
            .O(N__10044),
            .I(N__10018));
    InMux I__2376 (
            .O(N__10043),
            .I(N__10018));
    InMux I__2375 (
            .O(N__10042),
            .I(N__10015));
    InMux I__2374 (
            .O(N__10041),
            .I(N__10012));
    InMux I__2373 (
            .O(N__10040),
            .I(N__10008));
    InMux I__2372 (
            .O(N__10039),
            .I(N__10001));
    InMux I__2371 (
            .O(N__10036),
            .I(N__10001));
    InMux I__2370 (
            .O(N__10035),
            .I(N__10001));
    InMux I__2369 (
            .O(N__10034),
            .I(N__9994));
    InMux I__2368 (
            .O(N__10033),
            .I(N__9994));
    InMux I__2367 (
            .O(N__10032),
            .I(N__9994));
    InMux I__2366 (
            .O(N__10031),
            .I(N__9989));
    InMux I__2365 (
            .O(N__10028),
            .I(N__9984));
    InMux I__2364 (
            .O(N__10027),
            .I(N__9984));
    InMux I__2363 (
            .O(N__10026),
            .I(N__9981));
    Span4Mux_v I__2362 (
            .O(N__10023),
            .I(N__9974));
    LocalMux I__2361 (
            .O(N__10018),
            .I(N__9974));
    LocalMux I__2360 (
            .O(N__10015),
            .I(N__9974));
    LocalMux I__2359 (
            .O(N__10012),
            .I(N__9971));
    InMux I__2358 (
            .O(N__10011),
            .I(N__9968));
    LocalMux I__2357 (
            .O(N__10008),
            .I(N__9964));
    LocalMux I__2356 (
            .O(N__10001),
            .I(N__9959));
    LocalMux I__2355 (
            .O(N__9994),
            .I(N__9959));
    InMux I__2354 (
            .O(N__9993),
            .I(N__9956));
    InMux I__2353 (
            .O(N__9992),
            .I(N__9953));
    LocalMux I__2352 (
            .O(N__9989),
            .I(N__9950));
    LocalMux I__2351 (
            .O(N__9984),
            .I(N__9945));
    LocalMux I__2350 (
            .O(N__9981),
            .I(N__9945));
    Span4Mux_h I__2349 (
            .O(N__9974),
            .I(N__9939));
    Span4Mux_v I__2348 (
            .O(N__9971),
            .I(N__9939));
    LocalMux I__2347 (
            .O(N__9968),
            .I(N__9936));
    InMux I__2346 (
            .O(N__9967),
            .I(N__9933));
    Span4Mux_v I__2345 (
            .O(N__9964),
            .I(N__9930));
    Span4Mux_v I__2344 (
            .O(N__9959),
            .I(N__9923));
    LocalMux I__2343 (
            .O(N__9956),
            .I(N__9923));
    LocalMux I__2342 (
            .O(N__9953),
            .I(N__9923));
    Span4Mux_v I__2341 (
            .O(N__9950),
            .I(N__9918));
    Span4Mux_v I__2340 (
            .O(N__9945),
            .I(N__9918));
    InMux I__2339 (
            .O(N__9944),
            .I(N__9915));
    Span4Mux_h I__2338 (
            .O(N__9939),
            .I(N__9910));
    Span4Mux_v I__2337 (
            .O(N__9936),
            .I(N__9910));
    LocalMux I__2336 (
            .O(N__9933),
            .I(N__9907));
    Span4Mux_h I__2335 (
            .O(N__9930),
            .I(N__9902));
    Span4Mux_v I__2334 (
            .O(N__9923),
            .I(N__9902));
    Sp12to4 I__2333 (
            .O(N__9918),
            .I(N__9897));
    LocalMux I__2332 (
            .O(N__9915),
            .I(N__9897));
    Span4Mux_h I__2331 (
            .O(N__9910),
            .I(N__9894));
    Span12Mux_v I__2330 (
            .O(N__9907),
            .I(N__9891));
    Sp12to4 I__2329 (
            .O(N__9902),
            .I(N__9888));
    Span12Mux_h I__2328 (
            .O(N__9897),
            .I(N__9883));
    Sp12to4 I__2327 (
            .O(N__9894),
            .I(N__9883));
    Span12Mux_h I__2326 (
            .O(N__9891),
            .I(N__9880));
    Span12Mux_h I__2325 (
            .O(N__9888),
            .I(N__9877));
    Span12Mux_v I__2324 (
            .O(N__9883),
            .I(N__9874));
    Odrv12 I__2323 (
            .O(N__9880),
            .I(AGNUS_REV_c));
    Odrv12 I__2322 (
            .O(N__9877),
            .I(AGNUS_REV_c));
    Odrv12 I__2321 (
            .O(N__9874),
            .I(AGNUS_REV_c));
    InMux I__2320 (
            .O(N__9867),
            .I(N__9864));
    LocalMux I__2319 (
            .O(N__9864),
            .I(N__9861));
    Odrv12 I__2318 (
            .O(N__9861),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    ClkMux I__2317 (
            .O(N__9858),
            .I(N__9834));
    ClkMux I__2316 (
            .O(N__9857),
            .I(N__9834));
    ClkMux I__2315 (
            .O(N__9856),
            .I(N__9834));
    ClkMux I__2314 (
            .O(N__9855),
            .I(N__9834));
    ClkMux I__2313 (
            .O(N__9854),
            .I(N__9834));
    ClkMux I__2312 (
            .O(N__9853),
            .I(N__9834));
    ClkMux I__2311 (
            .O(N__9852),
            .I(N__9834));
    ClkMux I__2310 (
            .O(N__9851),
            .I(N__9834));
    GlobalMux I__2309 (
            .O(N__9834),
            .I(N__9831));
    gio2CtrlBuf I__2308 (
            .O(N__9831),
            .I(C3_c_g));
    CEMux I__2307 (
            .O(N__9828),
            .I(N__9789));
    CEMux I__2306 (
            .O(N__9827),
            .I(N__9789));
    CEMux I__2305 (
            .O(N__9826),
            .I(N__9789));
    CEMux I__2304 (
            .O(N__9825),
            .I(N__9789));
    CEMux I__2303 (
            .O(N__9824),
            .I(N__9789));
    CEMux I__2302 (
            .O(N__9823),
            .I(N__9789));
    CEMux I__2301 (
            .O(N__9822),
            .I(N__9789));
    CEMux I__2300 (
            .O(N__9821),
            .I(N__9789));
    CEMux I__2299 (
            .O(N__9820),
            .I(N__9789));
    CEMux I__2298 (
            .O(N__9819),
            .I(N__9789));
    CEMux I__2297 (
            .O(N__9818),
            .I(N__9789));
    CEMux I__2296 (
            .O(N__9817),
            .I(N__9789));
    CEMux I__2295 (
            .O(N__9816),
            .I(N__9789));
    GlobalMux I__2294 (
            .O(N__9789),
            .I(N__9786));
    gio2CtrlBuf I__2293 (
            .O(N__9786),
            .I(DBRn_c_i_0_g));
    IoInMux I__2292 (
            .O(N__9783),
            .I(N__9780));
    LocalMux I__2291 (
            .O(N__9780),
            .I(N__9777));
    Span4Mux_s2_v I__2290 (
            .O(N__9777),
            .I(N__9774));
    Span4Mux_h I__2289 (
            .O(N__9774),
            .I(N__9771));
    Span4Mux_v I__2288 (
            .O(N__9771),
            .I(N__9768));
    Odrv4 I__2287 (
            .O(N__9768),
            .I(N_216_i));
    InMux I__2286 (
            .O(N__9765),
            .I(N__9761));
    CascadeMux I__2285 (
            .O(N__9764),
            .I(N__9758));
    LocalMux I__2284 (
            .O(N__9761),
            .I(N__9755));
    InMux I__2283 (
            .O(N__9758),
            .I(N__9752));
    Span4Mux_v I__2282 (
            .O(N__9755),
            .I(N__9744));
    LocalMux I__2281 (
            .O(N__9752),
            .I(N__9744));
    InMux I__2280 (
            .O(N__9751),
            .I(N__9741));
    InMux I__2279 (
            .O(N__9750),
            .I(N__9738));
    InMux I__2278 (
            .O(N__9749),
            .I(N__9735));
    Span4Mux_h I__2277 (
            .O(N__9744),
            .I(N__9730));
    LocalMux I__2276 (
            .O(N__9741),
            .I(N__9727));
    LocalMux I__2275 (
            .O(N__9738),
            .I(N__9722));
    LocalMux I__2274 (
            .O(N__9735),
            .I(N__9722));
    InMux I__2273 (
            .O(N__9734),
            .I(N__9719));
    CascadeMux I__2272 (
            .O(N__9733),
            .I(N__9716));
    Span4Mux_v I__2271 (
            .O(N__9730),
            .I(N__9713));
    Span4Mux_v I__2270 (
            .O(N__9727),
            .I(N__9710));
    Span4Mux_h I__2269 (
            .O(N__9722),
            .I(N__9705));
    LocalMux I__2268 (
            .O(N__9719),
            .I(N__9705));
    InMux I__2267 (
            .O(N__9716),
            .I(N__9702));
    Span4Mux_h I__2266 (
            .O(N__9713),
            .I(N__9699));
    Span4Mux_h I__2265 (
            .O(N__9710),
            .I(N__9696));
    Span4Mux_h I__2264 (
            .O(N__9705),
            .I(N__9693));
    LocalMux I__2263 (
            .O(N__9702),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2262 (
            .O(N__9699),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2261 (
            .O(N__9696),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2260 (
            .O(N__9693),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__2259 (
            .O(N__9684),
            .I(N__9681));
    LocalMux I__2258 (
            .O(N__9681),
            .I(N__9678));
    IoSpan4Mux I__2257 (
            .O(N__9678),
            .I(N__9675));
    Span4Mux_s2_v I__2256 (
            .O(N__9675),
            .I(N__9672));
    Span4Mux_v I__2255 (
            .O(N__9672),
            .I(N__9669));
    Span4Mux_v I__2254 (
            .O(N__9669),
            .I(N__9666));
    Odrv4 I__2253 (
            .O(N__9666),
            .I(RASn_c));
    InMux I__2252 (
            .O(N__9663),
            .I(N__9660));
    LocalMux I__2251 (
            .O(N__9660),
            .I(N__9626));
    ClkMux I__2250 (
            .O(N__9659),
            .I(N__9531));
    ClkMux I__2249 (
            .O(N__9658),
            .I(N__9531));
    ClkMux I__2248 (
            .O(N__9657),
            .I(N__9531));
    ClkMux I__2247 (
            .O(N__9656),
            .I(N__9531));
    ClkMux I__2246 (
            .O(N__9655),
            .I(N__9531));
    ClkMux I__2245 (
            .O(N__9654),
            .I(N__9531));
    ClkMux I__2244 (
            .O(N__9653),
            .I(N__9531));
    ClkMux I__2243 (
            .O(N__9652),
            .I(N__9531));
    ClkMux I__2242 (
            .O(N__9651),
            .I(N__9531));
    ClkMux I__2241 (
            .O(N__9650),
            .I(N__9531));
    ClkMux I__2240 (
            .O(N__9649),
            .I(N__9531));
    ClkMux I__2239 (
            .O(N__9648),
            .I(N__9531));
    ClkMux I__2238 (
            .O(N__9647),
            .I(N__9531));
    ClkMux I__2237 (
            .O(N__9646),
            .I(N__9531));
    ClkMux I__2236 (
            .O(N__9645),
            .I(N__9531));
    ClkMux I__2235 (
            .O(N__9644),
            .I(N__9531));
    ClkMux I__2234 (
            .O(N__9643),
            .I(N__9531));
    ClkMux I__2233 (
            .O(N__9642),
            .I(N__9531));
    ClkMux I__2232 (
            .O(N__9641),
            .I(N__9531));
    ClkMux I__2231 (
            .O(N__9640),
            .I(N__9531));
    ClkMux I__2230 (
            .O(N__9639),
            .I(N__9531));
    ClkMux I__2229 (
            .O(N__9638),
            .I(N__9531));
    ClkMux I__2228 (
            .O(N__9637),
            .I(N__9531));
    ClkMux I__2227 (
            .O(N__9636),
            .I(N__9531));
    ClkMux I__2226 (
            .O(N__9635),
            .I(N__9531));
    ClkMux I__2225 (
            .O(N__9634),
            .I(N__9531));
    ClkMux I__2224 (
            .O(N__9633),
            .I(N__9531));
    ClkMux I__2223 (
            .O(N__9632),
            .I(N__9531));
    ClkMux I__2222 (
            .O(N__9631),
            .I(N__9531));
    ClkMux I__2221 (
            .O(N__9630),
            .I(N__9531));
    ClkMux I__2220 (
            .O(N__9629),
            .I(N__9531));
    Glb2LocalMux I__2219 (
            .O(N__9626),
            .I(N__9531));
    ClkMux I__2218 (
            .O(N__9625),
            .I(N__9531));
    ClkMux I__2217 (
            .O(N__9624),
            .I(N__9531));
    ClkMux I__2216 (
            .O(N__9623),
            .I(N__9531));
    ClkMux I__2215 (
            .O(N__9622),
            .I(N__9531));
    ClkMux I__2214 (
            .O(N__9621),
            .I(N__9531));
    ClkMux I__2213 (
            .O(N__9620),
            .I(N__9531));
    ClkMux I__2212 (
            .O(N__9619),
            .I(N__9531));
    ClkMux I__2211 (
            .O(N__9618),
            .I(N__9531));
    ClkMux I__2210 (
            .O(N__9617),
            .I(N__9531));
    ClkMux I__2209 (
            .O(N__9616),
            .I(N__9531));
    GlobalMux I__2208 (
            .O(N__9531),
            .I(CLK80_PLL));
    InMux I__2207 (
            .O(N__9528),
            .I(N__9522));
    InMux I__2206 (
            .O(N__9527),
            .I(N__9522));
    LocalMux I__2205 (
            .O(N__9522),
            .I(N__9519));
    Odrv12 I__2204 (
            .O(N__9519),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__2203 (
            .O(N__9516),
            .I(N__9513));
    LocalMux I__2202 (
            .O(N__9513),
            .I(N__9510));
    Odrv4 I__2201 (
            .O(N__9510),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    CascadeMux I__2200 (
            .O(N__9507),
            .I(N__9504));
    InMux I__2199 (
            .O(N__9504),
            .I(N__9501));
    LocalMux I__2198 (
            .O(N__9501),
            .I(N__9498));
    Span4Mux_h I__2197 (
            .O(N__9498),
            .I(N__9495));
    Odrv4 I__2196 (
            .O(N__9495),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2195 (
            .O(N__9492),
            .I(N__9489));
    LocalMux I__2194 (
            .O(N__9489),
            .I(N__9486));
    Odrv4 I__2193 (
            .O(N__9486),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2192 (
            .O(N__9483),
            .I(N__9480));
    LocalMux I__2191 (
            .O(N__9480),
            .I(N__9477));
    Span4Mux_h I__2190 (
            .O(N__9477),
            .I(N__9474));
    Odrv4 I__2189 (
            .O(N__9474),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__2188 (
            .O(N__9471),
            .I(N__9468));
    LocalMux I__2187 (
            .O(N__9468),
            .I(N__9465));
    Span4Mux_h I__2186 (
            .O(N__9465),
            .I(N__9462));
    Odrv4 I__2185 (
            .O(N__9462),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__2184 (
            .O(N__9459),
            .I(N__9454));
    InMux I__2183 (
            .O(N__9458),
            .I(N__9451));
    InMux I__2182 (
            .O(N__9457),
            .I(N__9448));
    LocalMux I__2181 (
            .O(N__9454),
            .I(N__9445));
    LocalMux I__2180 (
            .O(N__9451),
            .I(N__9439));
    LocalMux I__2179 (
            .O(N__9448),
            .I(N__9439));
    Span4Mux_v I__2178 (
            .O(N__9445),
            .I(N__9436));
    InMux I__2177 (
            .O(N__9444),
            .I(N__9433));
    Span4Mux_h I__2176 (
            .O(N__9439),
            .I(N__9430));
    Span4Mux_v I__2175 (
            .O(N__9436),
            .I(N__9427));
    LocalMux I__2174 (
            .O(N__9433),
            .I(N__9424));
    Sp12to4 I__2173 (
            .O(N__9430),
            .I(N__9421));
    Sp12to4 I__2172 (
            .O(N__9427),
            .I(N__9416));
    Span12Mux_v I__2171 (
            .O(N__9424),
            .I(N__9416));
    Span12Mux_v I__2170 (
            .O(N__9421),
            .I(N__9413));
    Span12Mux_h I__2169 (
            .O(N__9416),
            .I(N__9410));
    Odrv12 I__2168 (
            .O(N__9413),
            .I(DRA_c_2));
    Odrv12 I__2167 (
            .O(N__9410),
            .I(DRA_c_2));
    InMux I__2166 (
            .O(N__9405),
            .I(N__9402));
    LocalMux I__2165 (
            .O(N__9402),
            .I(N__9399));
    Span4Mux_h I__2164 (
            .O(N__9399),
            .I(N__9396));
    Odrv4 I__2163 (
            .O(N__9396),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    CascadeMux I__2162 (
            .O(N__9393),
            .I(N__9384));
    InMux I__2161 (
            .O(N__9392),
            .I(N__9380));
    CascadeMux I__2160 (
            .O(N__9391),
            .I(N__9375));
    InMux I__2159 (
            .O(N__9390),
            .I(N__9372));
    CascadeMux I__2158 (
            .O(N__9389),
            .I(N__9366));
    InMux I__2157 (
            .O(N__9388),
            .I(N__9360));
    InMux I__2156 (
            .O(N__9387),
            .I(N__9360));
    InMux I__2155 (
            .O(N__9384),
            .I(N__9356));
    InMux I__2154 (
            .O(N__9383),
            .I(N__9353));
    LocalMux I__2153 (
            .O(N__9380),
            .I(N__9350));
    InMux I__2152 (
            .O(N__9379),
            .I(N__9347));
    InMux I__2151 (
            .O(N__9378),
            .I(N__9341));
    InMux I__2150 (
            .O(N__9375),
            .I(N__9341));
    LocalMux I__2149 (
            .O(N__9372),
            .I(N__9337));
    InMux I__2148 (
            .O(N__9371),
            .I(N__9332));
    InMux I__2147 (
            .O(N__9370),
            .I(N__9332));
    InMux I__2146 (
            .O(N__9369),
            .I(N__9329));
    InMux I__2145 (
            .O(N__9366),
            .I(N__9325));
    InMux I__2144 (
            .O(N__9365),
            .I(N__9322));
    LocalMux I__2143 (
            .O(N__9360),
            .I(N__9318));
    InMux I__2142 (
            .O(N__9359),
            .I(N__9315));
    LocalMux I__2141 (
            .O(N__9356),
            .I(N__9311));
    LocalMux I__2140 (
            .O(N__9353),
            .I(N__9308));
    Span4Mux_v I__2139 (
            .O(N__9350),
            .I(N__9301));
    LocalMux I__2138 (
            .O(N__9347),
            .I(N__9301));
    InMux I__2137 (
            .O(N__9346),
            .I(N__9298));
    LocalMux I__2136 (
            .O(N__9341),
            .I(N__9295));
    InMux I__2135 (
            .O(N__9340),
            .I(N__9290));
    Span4Mux_v I__2134 (
            .O(N__9337),
            .I(N__9285));
    LocalMux I__2133 (
            .O(N__9332),
            .I(N__9285));
    LocalMux I__2132 (
            .O(N__9329),
            .I(N__9282));
    InMux I__2131 (
            .O(N__9328),
            .I(N__9279));
    LocalMux I__2130 (
            .O(N__9325),
            .I(N__9274));
    LocalMux I__2129 (
            .O(N__9322),
            .I(N__9274));
    InMux I__2128 (
            .O(N__9321),
            .I(N__9271));
    Span4Mux_v I__2127 (
            .O(N__9318),
            .I(N__9266));
    LocalMux I__2126 (
            .O(N__9315),
            .I(N__9266));
    InMux I__2125 (
            .O(N__9314),
            .I(N__9263));
    Span4Mux_h I__2124 (
            .O(N__9311),
            .I(N__9258));
    Span4Mux_h I__2123 (
            .O(N__9308),
            .I(N__9258));
    InMux I__2122 (
            .O(N__9307),
            .I(N__9253));
    InMux I__2121 (
            .O(N__9306),
            .I(N__9253));
    Span4Mux_v I__2120 (
            .O(N__9301),
            .I(N__9246));
    LocalMux I__2119 (
            .O(N__9298),
            .I(N__9246));
    Span4Mux_v I__2118 (
            .O(N__9295),
            .I(N__9246));
    InMux I__2117 (
            .O(N__9294),
            .I(N__9241));
    InMux I__2116 (
            .O(N__9293),
            .I(N__9241));
    LocalMux I__2115 (
            .O(N__9290),
            .I(N__9236));
    Span4Mux_h I__2114 (
            .O(N__9285),
            .I(N__9236));
    Span12Mux_h I__2113 (
            .O(N__9282),
            .I(N__9227));
    LocalMux I__2112 (
            .O(N__9279),
            .I(N__9227));
    Span12Mux_h I__2111 (
            .O(N__9274),
            .I(N__9227));
    LocalMux I__2110 (
            .O(N__9271),
            .I(N__9227));
    Odrv4 I__2109 (
            .O(N__9266),
            .I(CPU_CYCLEm));
    LocalMux I__2108 (
            .O(N__9263),
            .I(CPU_CYCLEm));
    Odrv4 I__2107 (
            .O(N__9258),
            .I(CPU_CYCLEm));
    LocalMux I__2106 (
            .O(N__9253),
            .I(CPU_CYCLEm));
    Odrv4 I__2105 (
            .O(N__9246),
            .I(CPU_CYCLEm));
    LocalMux I__2104 (
            .O(N__9241),
            .I(CPU_CYCLEm));
    Odrv4 I__2103 (
            .O(N__9236),
            .I(CPU_CYCLEm));
    Odrv12 I__2102 (
            .O(N__9227),
            .I(CPU_CYCLEm));
    InMux I__2101 (
            .O(N__9210),
            .I(N__9207));
    LocalMux I__2100 (
            .O(N__9207),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    InMux I__2099 (
            .O(N__9204),
            .I(N__9196));
    InMux I__2098 (
            .O(N__9203),
            .I(N__9191));
    CascadeMux I__2097 (
            .O(N__9202),
            .I(N__9188));
    CascadeMux I__2096 (
            .O(N__9201),
            .I(N__9185));
    CascadeMux I__2095 (
            .O(N__9200),
            .I(N__9182));
    CascadeMux I__2094 (
            .O(N__9199),
            .I(N__9177));
    LocalMux I__2093 (
            .O(N__9196),
            .I(N__9170));
    InMux I__2092 (
            .O(N__9195),
            .I(N__9167));
    InMux I__2091 (
            .O(N__9194),
            .I(N__9164));
    LocalMux I__2090 (
            .O(N__9191),
            .I(N__9161));
    InMux I__2089 (
            .O(N__9188),
            .I(N__9158));
    InMux I__2088 (
            .O(N__9185),
            .I(N__9155));
    InMux I__2087 (
            .O(N__9182),
            .I(N__9150));
    InMux I__2086 (
            .O(N__9181),
            .I(N__9144));
    InMux I__2085 (
            .O(N__9180),
            .I(N__9144));
    InMux I__2084 (
            .O(N__9177),
            .I(N__9137));
    InMux I__2083 (
            .O(N__9176),
            .I(N__9137));
    InMux I__2082 (
            .O(N__9175),
            .I(N__9137));
    InMux I__2081 (
            .O(N__9174),
            .I(N__9130));
    InMux I__2080 (
            .O(N__9173),
            .I(N__9130));
    Span4Mux_h I__2079 (
            .O(N__9170),
            .I(N__9122));
    LocalMux I__2078 (
            .O(N__9167),
            .I(N__9122));
    LocalMux I__2077 (
            .O(N__9164),
            .I(N__9113));
    Span4Mux_v I__2076 (
            .O(N__9161),
            .I(N__9113));
    LocalMux I__2075 (
            .O(N__9158),
            .I(N__9113));
    LocalMux I__2074 (
            .O(N__9155),
            .I(N__9113));
    InMux I__2073 (
            .O(N__9154),
            .I(N__9108));
    InMux I__2072 (
            .O(N__9153),
            .I(N__9108));
    LocalMux I__2071 (
            .O(N__9150),
            .I(N__9105));
    InMux I__2070 (
            .O(N__9149),
            .I(N__9101));
    LocalMux I__2069 (
            .O(N__9144),
            .I(N__9098));
    LocalMux I__2068 (
            .O(N__9137),
            .I(N__9095));
    InMux I__2067 (
            .O(N__9136),
            .I(N__9090));
    InMux I__2066 (
            .O(N__9135),
            .I(N__9090));
    LocalMux I__2065 (
            .O(N__9130),
            .I(N__9087));
    InMux I__2064 (
            .O(N__9129),
            .I(N__9082));
    InMux I__2063 (
            .O(N__9128),
            .I(N__9082));
    InMux I__2062 (
            .O(N__9127),
            .I(N__9079));
    Span4Mux_h I__2061 (
            .O(N__9122),
            .I(N__9075));
    Span4Mux_v I__2060 (
            .O(N__9113),
            .I(N__9072));
    LocalMux I__2059 (
            .O(N__9108),
            .I(N__9069));
    Span4Mux_h I__2058 (
            .O(N__9105),
            .I(N__9066));
    InMux I__2057 (
            .O(N__9104),
            .I(N__9063));
    LocalMux I__2056 (
            .O(N__9101),
            .I(N__9048));
    Span4Mux_v I__2055 (
            .O(N__9098),
            .I(N__9048));
    Span4Mux_v I__2054 (
            .O(N__9095),
            .I(N__9048));
    LocalMux I__2053 (
            .O(N__9090),
            .I(N__9048));
    Span4Mux_h I__2052 (
            .O(N__9087),
            .I(N__9048));
    LocalMux I__2051 (
            .O(N__9082),
            .I(N__9048));
    LocalMux I__2050 (
            .O(N__9079),
            .I(N__9048));
    InMux I__2049 (
            .O(N__9078),
            .I(N__9045));
    Span4Mux_v I__2048 (
            .O(N__9075),
            .I(N__9042));
    Span4Mux_h I__2047 (
            .O(N__9072),
            .I(N__9037));
    Span4Mux_v I__2046 (
            .O(N__9069),
            .I(N__9037));
    Sp12to4 I__2045 (
            .O(N__9066),
            .I(N__9032));
    LocalMux I__2044 (
            .O(N__9063),
            .I(N__9032));
    Span4Mux_h I__2043 (
            .O(N__9048),
            .I(N__9029));
    LocalMux I__2042 (
            .O(N__9045),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2041 (
            .O(N__9042),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2040 (
            .O(N__9037),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__2039 (
            .O(N__9032),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2038 (
            .O(N__9029),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    InMux I__2037 (
            .O(N__9018),
            .I(N__9015));
    LocalMux I__2036 (
            .O(N__9015),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    InMux I__2035 (
            .O(N__9012),
            .I(N__9009));
    LocalMux I__2034 (
            .O(N__9009),
            .I(N__9006));
    Odrv4 I__2033 (
            .O(N__9006),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2032 (
            .O(N__9003),
            .I(N__9000));
    LocalMux I__2031 (
            .O(N__9000),
            .I(N__8997));
    Span4Mux_h I__2030 (
            .O(N__8997),
            .I(N__8994));
    Odrv4 I__2029 (
            .O(N__8994),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__2028 (
            .O(N__8991),
            .I(N__8987));
    InMux I__2027 (
            .O(N__8990),
            .I(N__8984));
    LocalMux I__2026 (
            .O(N__8987),
            .I(N__8981));
    LocalMux I__2025 (
            .O(N__8984),
            .I(N__8978));
    Span4Mux_h I__2024 (
            .O(N__8981),
            .I(N__8975));
    Span4Mux_v I__2023 (
            .O(N__8978),
            .I(N__8972));
    Sp12to4 I__2022 (
            .O(N__8975),
            .I(N__8969));
    Sp12to4 I__2021 (
            .O(N__8972),
            .I(N__8966));
    Span12Mux_v I__2020 (
            .O(N__8969),
            .I(N__8963));
    Span12Mux_h I__2019 (
            .O(N__8966),
            .I(N__8960));
    Span12Mux_h I__2018 (
            .O(N__8963),
            .I(N__8955));
    Span12Mux_v I__2017 (
            .O(N__8960),
            .I(N__8955));
    Odrv12 I__2016 (
            .O(N__8955),
            .I(DRA_c_0));
    InMux I__2015 (
            .O(N__8952),
            .I(N__8949));
    LocalMux I__2014 (
            .O(N__8949),
            .I(N__8946));
    Odrv12 I__2013 (
            .O(N__8946),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__2012 (
            .O(N__8943),
            .I(N__8940));
    LocalMux I__2011 (
            .O(N__8940),
            .I(N__8934));
    InMux I__2010 (
            .O(N__8939),
            .I(N__8929));
    InMux I__2009 (
            .O(N__8938),
            .I(N__8929));
    InMux I__2008 (
            .O(N__8937),
            .I(N__8926));
    Sp12to4 I__2007 (
            .O(N__8934),
            .I(N__8919));
    LocalMux I__2006 (
            .O(N__8929),
            .I(N__8919));
    LocalMux I__2005 (
            .O(N__8926),
            .I(N__8919));
    Span12Mux_v I__2004 (
            .O(N__8919),
            .I(N__8916));
    Span12Mux_h I__2003 (
            .O(N__8916),
            .I(N__8913));
    Odrv12 I__2002 (
            .O(N__8913),
            .I(DRA_c_1));
    InMux I__2001 (
            .O(N__8910),
            .I(N__8904));
    InMux I__2000 (
            .O(N__8909),
            .I(N__8904));
    LocalMux I__1999 (
            .O(N__8904),
            .I(N__8901));
    Span4Mux_v I__1998 (
            .O(N__8901),
            .I(N__8898));
    Odrv4 I__1997 (
            .O(N__8898),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    IoInMux I__1996 (
            .O(N__8895),
            .I(N__8892));
    LocalMux I__1995 (
            .O(N__8892),
            .I(N__8889));
    Span4Mux_s0_v I__1994 (
            .O(N__8889),
            .I(N__8886));
    Span4Mux_v I__1993 (
            .O(N__8886),
            .I(N__8883));
    Odrv4 I__1992 (
            .O(N__8883),
            .I(U712_BYTE_ENABLE_UUBE_i));
    IoInMux I__1991 (
            .O(N__8880),
            .I(N__8877));
    LocalMux I__1990 (
            .O(N__8877),
            .I(N__8874));
    Span4Mux_s2_v I__1989 (
            .O(N__8874),
            .I(N__8871));
    Span4Mux_v I__1988 (
            .O(N__8871),
            .I(N__8868));
    Odrv4 I__1987 (
            .O(N__8868),
            .I(N_215_i));
    IoInMux I__1986 (
            .O(N__8865),
            .I(N__8862));
    LocalMux I__1985 (
            .O(N__8862),
            .I(N__8859));
    IoSpan4Mux I__1984 (
            .O(N__8859),
            .I(N__8856));
    Span4Mux_s3_v I__1983 (
            .O(N__8856),
            .I(N__8853));
    Odrv4 I__1982 (
            .O(N__8853),
            .I(N_217_i));
    InMux I__1981 (
            .O(N__8850),
            .I(N__8844));
    InMux I__1980 (
            .O(N__8849),
            .I(N__8835));
    InMux I__1979 (
            .O(N__8848),
            .I(N__8835));
    InMux I__1978 (
            .O(N__8847),
            .I(N__8835));
    LocalMux I__1977 (
            .O(N__8844),
            .I(N__8832));
    InMux I__1976 (
            .O(N__8843),
            .I(N__8829));
    InMux I__1975 (
            .O(N__8842),
            .I(N__8826));
    LocalMux I__1974 (
            .O(N__8835),
            .I(N__8823));
    Span4Mux_h I__1973 (
            .O(N__8832),
            .I(N__8817));
    LocalMux I__1972 (
            .O(N__8829),
            .I(N__8817));
    LocalMux I__1971 (
            .O(N__8826),
            .I(N__8813));
    Span4Mux_v I__1970 (
            .O(N__8823),
            .I(N__8810));
    InMux I__1969 (
            .O(N__8822),
            .I(N__8807));
    Span4Mux_h I__1968 (
            .O(N__8817),
            .I(N__8804));
    InMux I__1967 (
            .O(N__8816),
            .I(N__8801));
    Span12Mux_v I__1966 (
            .O(N__8813),
            .I(N__8798));
    Sp12to4 I__1965 (
            .O(N__8810),
            .I(N__8793));
    LocalMux I__1964 (
            .O(N__8807),
            .I(N__8793));
    Span4Mux_v I__1963 (
            .O(N__8804),
            .I(N__8790));
    LocalMux I__1962 (
            .O(N__8801),
            .I(N__8787));
    Span12Mux_h I__1961 (
            .O(N__8798),
            .I(N__8784));
    Span12Mux_h I__1960 (
            .O(N__8793),
            .I(N__8777));
    Sp12to4 I__1959 (
            .O(N__8790),
            .I(N__8777));
    Span12Mux_v I__1958 (
            .O(N__8787),
            .I(N__8777));
    Odrv12 I__1957 (
            .O(N__8784),
            .I(A_c_1));
    Odrv12 I__1956 (
            .O(N__8777),
            .I(A_c_1));
    InMux I__1955 (
            .O(N__8772),
            .I(N__8759));
    InMux I__1954 (
            .O(N__8771),
            .I(N__8759));
    InMux I__1953 (
            .O(N__8770),
            .I(N__8759));
    InMux I__1952 (
            .O(N__8769),
            .I(N__8756));
    InMux I__1951 (
            .O(N__8768),
            .I(N__8753));
    InMux I__1950 (
            .O(N__8767),
            .I(N__8750));
    InMux I__1949 (
            .O(N__8766),
            .I(N__8747));
    LocalMux I__1948 (
            .O(N__8759),
            .I(N__8741));
    LocalMux I__1947 (
            .O(N__8756),
            .I(N__8741));
    LocalMux I__1946 (
            .O(N__8753),
            .I(N__8736));
    LocalMux I__1945 (
            .O(N__8750),
            .I(N__8736));
    LocalMux I__1944 (
            .O(N__8747),
            .I(N__8733));
    InMux I__1943 (
            .O(N__8746),
            .I(N__8729));
    Span4Mux_v I__1942 (
            .O(N__8741),
            .I(N__8725));
    Span4Mux_v I__1941 (
            .O(N__8736),
            .I(N__8720));
    Span4Mux_v I__1940 (
            .O(N__8733),
            .I(N__8720));
    InMux I__1939 (
            .O(N__8732),
            .I(N__8717));
    LocalMux I__1938 (
            .O(N__8729),
            .I(N__8714));
    InMux I__1937 (
            .O(N__8728),
            .I(N__8711));
    Sp12to4 I__1936 (
            .O(N__8725),
            .I(N__8704));
    Sp12to4 I__1935 (
            .O(N__8720),
            .I(N__8704));
    LocalMux I__1934 (
            .O(N__8717),
            .I(N__8704));
    Span4Mux_v I__1933 (
            .O(N__8714),
            .I(N__8701));
    LocalMux I__1932 (
            .O(N__8711),
            .I(N__8698));
    Span12Mux_h I__1931 (
            .O(N__8704),
            .I(N__8695));
    Sp12to4 I__1930 (
            .O(N__8701),
            .I(N__8690));
    Span12Mux_v I__1929 (
            .O(N__8698),
            .I(N__8690));
    Odrv12 I__1928 (
            .O(N__8695),
            .I(A_c_0));
    Odrv12 I__1927 (
            .O(N__8690),
            .I(A_c_0));
    CascadeMux I__1926 (
            .O(N__8685),
            .I(N__8679));
    CascadeMux I__1925 (
            .O(N__8684),
            .I(N__8675));
    CascadeMux I__1924 (
            .O(N__8683),
            .I(N__8672));
    CascadeMux I__1923 (
            .O(N__8682),
            .I(N__8669));
    InMux I__1922 (
            .O(N__8679),
            .I(N__8665));
    InMux I__1921 (
            .O(N__8678),
            .I(N__8662));
    InMux I__1920 (
            .O(N__8675),
            .I(N__8655));
    InMux I__1919 (
            .O(N__8672),
            .I(N__8655));
    InMux I__1918 (
            .O(N__8669),
            .I(N__8655));
    CascadeMux I__1917 (
            .O(N__8668),
            .I(N__8652));
    LocalMux I__1916 (
            .O(N__8665),
            .I(N__8649));
    LocalMux I__1915 (
            .O(N__8662),
            .I(N__8646));
    LocalMux I__1914 (
            .O(N__8655),
            .I(N__8643));
    InMux I__1913 (
            .O(N__8652),
            .I(N__8640));
    Span4Mux_h I__1912 (
            .O(N__8649),
            .I(N__8634));
    Span4Mux_v I__1911 (
            .O(N__8646),
            .I(N__8634));
    Span4Mux_h I__1910 (
            .O(N__8643),
            .I(N__8629));
    LocalMux I__1909 (
            .O(N__8640),
            .I(N__8629));
    InMux I__1908 (
            .O(N__8639),
            .I(N__8626));
    Span4Mux_v I__1907 (
            .O(N__8634),
            .I(N__8621));
    Span4Mux_h I__1906 (
            .O(N__8629),
            .I(N__8621));
    LocalMux I__1905 (
            .O(N__8626),
            .I(N__8618));
    Span4Mux_v I__1904 (
            .O(N__8621),
            .I(N__8615));
    Span12Mux_v I__1903 (
            .O(N__8618),
            .I(N__8610));
    Sp12to4 I__1902 (
            .O(N__8615),
            .I(N__8610));
    Odrv12 I__1901 (
            .O(N__8610),
            .I(SIZ_c_0));
    CascadeMux I__1900 (
            .O(N__8607),
            .I(N__8602));
    CascadeMux I__1899 (
            .O(N__8606),
            .I(N__8599));
    InMux I__1898 (
            .O(N__8605),
            .I(N__8593));
    InMux I__1897 (
            .O(N__8602),
            .I(N__8590));
    InMux I__1896 (
            .O(N__8599),
            .I(N__8587));
    InMux I__1895 (
            .O(N__8598),
            .I(N__8580));
    InMux I__1894 (
            .O(N__8597),
            .I(N__8580));
    InMux I__1893 (
            .O(N__8596),
            .I(N__8580));
    LocalMux I__1892 (
            .O(N__8593),
            .I(N__8576));
    LocalMux I__1891 (
            .O(N__8590),
            .I(N__8573));
    LocalMux I__1890 (
            .O(N__8587),
            .I(N__8570));
    LocalMux I__1889 (
            .O(N__8580),
            .I(N__8567));
    InMux I__1888 (
            .O(N__8579),
            .I(N__8564));
    Span4Mux_h I__1887 (
            .O(N__8576),
            .I(N__8557));
    Span4Mux_v I__1886 (
            .O(N__8573),
            .I(N__8557));
    Span4Mux_v I__1885 (
            .O(N__8570),
            .I(N__8557));
    Span4Mux_h I__1884 (
            .O(N__8567),
            .I(N__8552));
    LocalMux I__1883 (
            .O(N__8564),
            .I(N__8552));
    Span4Mux_v I__1882 (
            .O(N__8557),
            .I(N__8547));
    Span4Mux_h I__1881 (
            .O(N__8552),
            .I(N__8547));
    Span4Mux_v I__1880 (
            .O(N__8547),
            .I(N__8544));
    Span4Mux_h I__1879 (
            .O(N__8544),
            .I(N__8541));
    Sp12to4 I__1878 (
            .O(N__8541),
            .I(N__8538));
    Odrv12 I__1877 (
            .O(N__8538),
            .I(SIZ_c_1));
    IoInMux I__1876 (
            .O(N__8535),
            .I(N__8532));
    LocalMux I__1875 (
            .O(N__8532),
            .I(N__8529));
    Span4Mux_s3_h I__1874 (
            .O(N__8529),
            .I(N__8526));
    Span4Mux_v I__1873 (
            .O(N__8526),
            .I(N__8523));
    Sp12to4 I__1872 (
            .O(N__8523),
            .I(N__8520));
    Span12Mux_h I__1871 (
            .O(N__8520),
            .I(N__8517));
    Odrv12 I__1870 (
            .O(N__8517),
            .I(WEn_c));
    IoInMux I__1869 (
            .O(N__8514),
            .I(N__8511));
    LocalMux I__1868 (
            .O(N__8511),
            .I(N__8508));
    Span4Mux_s0_v I__1867 (
            .O(N__8508),
            .I(N__8505));
    Sp12to4 I__1866 (
            .O(N__8505),
            .I(N__8502));
    Span12Mux_h I__1865 (
            .O(N__8502),
            .I(N__8499));
    Odrv12 I__1864 (
            .O(N__8499),
            .I(CASn_c));
    IoInMux I__1863 (
            .O(N__8496),
            .I(N__8493));
    LocalMux I__1862 (
            .O(N__8493),
            .I(N__8490));
    IoSpan4Mux I__1861 (
            .O(N__8490),
            .I(N__8487));
    Span4Mux_s2_v I__1860 (
            .O(N__8487),
            .I(N__8484));
    Span4Mux_v I__1859 (
            .O(N__8484),
            .I(N__8481));
    Span4Mux_v I__1858 (
            .O(N__8481),
            .I(N__8478));
    Odrv4 I__1857 (
            .O(N__8478),
            .I(CRCSn_c));
    InMux I__1856 (
            .O(N__8475),
            .I(N__8472));
    LocalMux I__1855 (
            .O(N__8472),
            .I(N__8469));
    Odrv12 I__1854 (
            .O(N__8469),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    InMux I__1853 (
            .O(N__8466),
            .I(N__8461));
    CascadeMux I__1852 (
            .O(N__8465),
            .I(N__8458));
    InMux I__1851 (
            .O(N__8464),
            .I(N__8454));
    LocalMux I__1850 (
            .O(N__8461),
            .I(N__8451));
    InMux I__1849 (
            .O(N__8458),
            .I(N__8448));
    CascadeMux I__1848 (
            .O(N__8457),
            .I(N__8445));
    LocalMux I__1847 (
            .O(N__8454),
            .I(N__8442));
    Span4Mux_h I__1846 (
            .O(N__8451),
            .I(N__8439));
    LocalMux I__1845 (
            .O(N__8448),
            .I(N__8436));
    InMux I__1844 (
            .O(N__8445),
            .I(N__8433));
    Sp12to4 I__1843 (
            .O(N__8442),
            .I(N__8429));
    Span4Mux_v I__1842 (
            .O(N__8439),
            .I(N__8422));
    Span4Mux_h I__1841 (
            .O(N__8436),
            .I(N__8422));
    LocalMux I__1840 (
            .O(N__8433),
            .I(N__8422));
    InMux I__1839 (
            .O(N__8432),
            .I(N__8419));
    Span12Mux_v I__1838 (
            .O(N__8429),
            .I(N__8416));
    Span4Mux_h I__1837 (
            .O(N__8422),
            .I(N__8413));
    LocalMux I__1836 (
            .O(N__8419),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv12 I__1835 (
            .O(N__8416),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1834 (
            .O(N__8413),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    InMux I__1833 (
            .O(N__8406),
            .I(N__8400));
    InMux I__1832 (
            .O(N__8405),
            .I(N__8397));
    InMux I__1831 (
            .O(N__8404),
            .I(N__8394));
    InMux I__1830 (
            .O(N__8403),
            .I(N__8391));
    LocalMux I__1829 (
            .O(N__8400),
            .I(N__8386));
    LocalMux I__1828 (
            .O(N__8397),
            .I(N__8383));
    LocalMux I__1827 (
            .O(N__8394),
            .I(N__8380));
    LocalMux I__1826 (
            .O(N__8391),
            .I(N__8377));
    InMux I__1825 (
            .O(N__8390),
            .I(N__8374));
    CascadeMux I__1824 (
            .O(N__8389),
            .I(N__8370));
    Span4Mux_v I__1823 (
            .O(N__8386),
            .I(N__8367));
    Span12Mux_h I__1822 (
            .O(N__8383),
            .I(N__8364));
    Span4Mux_v I__1821 (
            .O(N__8380),
            .I(N__8357));
    Span4Mux_h I__1820 (
            .O(N__8377),
            .I(N__8357));
    LocalMux I__1819 (
            .O(N__8374),
            .I(N__8357));
    InMux I__1818 (
            .O(N__8373),
            .I(N__8354));
    InMux I__1817 (
            .O(N__8370),
            .I(N__8351));
    Span4Mux_h I__1816 (
            .O(N__8367),
            .I(N__8348));
    Span12Mux_v I__1815 (
            .O(N__8364),
            .I(N__8345));
    Span4Mux_h I__1814 (
            .O(N__8357),
            .I(N__8342));
    LocalMux I__1813 (
            .O(N__8354),
            .I(N__8339));
    LocalMux I__1812 (
            .O(N__8351),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1811 (
            .O(N__8348),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv12 I__1810 (
            .O(N__8345),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1809 (
            .O(N__8342),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv12 I__1808 (
            .O(N__8339),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1807 (
            .O(N__8328),
            .I(N__8325));
    LocalMux I__1806 (
            .O(N__8325),
            .I(N__8322));
    Span4Mux_s3_v I__1805 (
            .O(N__8322),
            .I(N__8319));
    Sp12to4 I__1804 (
            .O(N__8319),
            .I(N__8316));
    Span12Mux_h I__1803 (
            .O(N__8316),
            .I(N__8313));
    Odrv12 I__1802 (
            .O(N__8313),
            .I(CMA_c_10));
    InMux I__1801 (
            .O(N__8310),
            .I(N__8307));
    LocalMux I__1800 (
            .O(N__8307),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    IoInMux I__1799 (
            .O(N__8304),
            .I(N__8301));
    LocalMux I__1798 (
            .O(N__8301),
            .I(N__8298));
    Span4Mux_s3_h I__1797 (
            .O(N__8298),
            .I(N__8295));
    Span4Mux_v I__1796 (
            .O(N__8295),
            .I(N__8292));
    Sp12to4 I__1795 (
            .O(N__8292),
            .I(N__8289));
    Span12Mux_h I__1794 (
            .O(N__8289),
            .I(N__8286));
    Odrv12 I__1793 (
            .O(N__8286),
            .I(CMA_c_4));
    InMux I__1792 (
            .O(N__8283),
            .I(N__8279));
    InMux I__1791 (
            .O(N__8282),
            .I(N__8276));
    LocalMux I__1790 (
            .O(N__8279),
            .I(N__8273));
    LocalMux I__1789 (
            .O(N__8276),
            .I(N__8270));
    Span4Mux_v I__1788 (
            .O(N__8273),
            .I(N__8263));
    Span4Mux_h I__1787 (
            .O(N__8270),
            .I(N__8260));
    InMux I__1786 (
            .O(N__8269),
            .I(N__8255));
    InMux I__1785 (
            .O(N__8268),
            .I(N__8255));
    InMux I__1784 (
            .O(N__8267),
            .I(N__8250));
    InMux I__1783 (
            .O(N__8266),
            .I(N__8250));
    Odrv4 I__1782 (
            .O(N__8263),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    Odrv4 I__1781 (
            .O(N__8260),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    LocalMux I__1780 (
            .O(N__8255),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    LocalMux I__1779 (
            .O(N__8250),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    CascadeMux I__1778 (
            .O(N__8241),
            .I(N__8238));
    InMux I__1777 (
            .O(N__8238),
            .I(N__8231));
    CascadeMux I__1776 (
            .O(N__8237),
            .I(N__8227));
    CascadeMux I__1775 (
            .O(N__8236),
            .I(N__8223));
    CascadeMux I__1774 (
            .O(N__8235),
            .I(N__8220));
    InMux I__1773 (
            .O(N__8234),
            .I(N__8216));
    LocalMux I__1772 (
            .O(N__8231),
            .I(N__8213));
    CascadeMux I__1771 (
            .O(N__8230),
            .I(N__8210));
    InMux I__1770 (
            .O(N__8227),
            .I(N__8207));
    InMux I__1769 (
            .O(N__8226),
            .I(N__8204));
    InMux I__1768 (
            .O(N__8223),
            .I(N__8201));
    InMux I__1767 (
            .O(N__8220),
            .I(N__8198));
    InMux I__1766 (
            .O(N__8219),
            .I(N__8195));
    LocalMux I__1765 (
            .O(N__8216),
            .I(N__8192));
    Span4Mux_v I__1764 (
            .O(N__8213),
            .I(N__8189));
    InMux I__1763 (
            .O(N__8210),
            .I(N__8186));
    LocalMux I__1762 (
            .O(N__8207),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1761 (
            .O(N__8204),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1760 (
            .O(N__8201),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1759 (
            .O(N__8198),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1758 (
            .O(N__8195),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv12 I__1757 (
            .O(N__8192),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__1756 (
            .O(N__8189),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1755 (
            .O(N__8186),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    IoInMux I__1754 (
            .O(N__8169),
            .I(N__8166));
    LocalMux I__1753 (
            .O(N__8166),
            .I(N__8163));
    Span4Mux_s2_h I__1752 (
            .O(N__8163),
            .I(N__8160));
    Sp12to4 I__1751 (
            .O(N__8160),
            .I(N__8157));
    Span12Mux_s9_v I__1750 (
            .O(N__8157),
            .I(N__8154));
    Span12Mux_h I__1749 (
            .O(N__8154),
            .I(N__8151));
    Odrv12 I__1748 (
            .O(N__8151),
            .I(CMA_c_6));
    InMux I__1747 (
            .O(N__8148),
            .I(N__8145));
    LocalMux I__1746 (
            .O(N__8145),
            .I(N__8140));
    InMux I__1745 (
            .O(N__8144),
            .I(N__8137));
    InMux I__1744 (
            .O(N__8143),
            .I(N__8134));
    Odrv4 I__1743 (
            .O(N__8140),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1742 (
            .O(N__8137),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1741 (
            .O(N__8134),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    InMux I__1740 (
            .O(N__8127),
            .I(N__8124));
    LocalMux I__1739 (
            .O(N__8124),
            .I(N__8121));
    Span4Mux_h I__1738 (
            .O(N__8121),
            .I(N__8118));
    Sp12to4 I__1737 (
            .O(N__8118),
            .I(N__8115));
    Span12Mux_v I__1736 (
            .O(N__8115),
            .I(N__8112));
    Span12Mux_h I__1735 (
            .O(N__8112),
            .I(N__8109));
    Odrv12 I__1734 (
            .O(N__8109),
            .I(A_c_19));
    IoInMux I__1733 (
            .O(N__8106),
            .I(N__8103));
    LocalMux I__1732 (
            .O(N__8103),
            .I(N__8100));
    IoSpan4Mux I__1731 (
            .O(N__8100),
            .I(N__8097));
    Span4Mux_s0_h I__1730 (
            .O(N__8097),
            .I(N__8094));
    Sp12to4 I__1729 (
            .O(N__8094),
            .I(N__8091));
    Span12Mux_h I__1728 (
            .O(N__8091),
            .I(N__8088));
    Odrv12 I__1727 (
            .O(N__8088),
            .I(CMA_c_9));
    CEMux I__1726 (
            .O(N__8085),
            .I(N__8077));
    CEMux I__1725 (
            .O(N__8084),
            .I(N__8074));
    CEMux I__1724 (
            .O(N__8083),
            .I(N__8070));
    CEMux I__1723 (
            .O(N__8082),
            .I(N__8067));
    CEMux I__1722 (
            .O(N__8081),
            .I(N__8064));
    CEMux I__1721 (
            .O(N__8080),
            .I(N__8061));
    LocalMux I__1720 (
            .O(N__8077),
            .I(N__8056));
    LocalMux I__1719 (
            .O(N__8074),
            .I(N__8056));
    CEMux I__1718 (
            .O(N__8073),
            .I(N__8053));
    LocalMux I__1717 (
            .O(N__8070),
            .I(N__8050));
    LocalMux I__1716 (
            .O(N__8067),
            .I(N__8047));
    LocalMux I__1715 (
            .O(N__8064),
            .I(N__8044));
    LocalMux I__1714 (
            .O(N__8061),
            .I(N__8041));
    Span4Mux_v I__1713 (
            .O(N__8056),
            .I(N__8036));
    LocalMux I__1712 (
            .O(N__8053),
            .I(N__8036));
    Span4Mux_v I__1711 (
            .O(N__8050),
            .I(N__8031));
    Span4Mux_h I__1710 (
            .O(N__8047),
            .I(N__8031));
    Span4Mux_h I__1709 (
            .O(N__8044),
            .I(N__8026));
    Span4Mux_h I__1708 (
            .O(N__8041),
            .I(N__8026));
    Span4Mux_v I__1707 (
            .O(N__8036),
            .I(N__8023));
    Odrv4 I__1706 (
            .O(N__8031),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__1705 (
            .O(N__8026),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__1704 (
            .O(N__8023),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    InMux I__1703 (
            .O(N__8016),
            .I(N__8010));
    InMux I__1702 (
            .O(N__8015),
            .I(N__8010));
    LocalMux I__1701 (
            .O(N__8010),
            .I(N__8007));
    Sp12to4 I__1700 (
            .O(N__8007),
            .I(N__8004));
    Span12Mux_v I__1699 (
            .O(N__8004),
            .I(N__8001));
    Span12Mux_h I__1698 (
            .O(N__8001),
            .I(N__7998));
    Odrv12 I__1697 (
            .O(N__7998),
            .I(A_c_14));
    CascadeMux I__1696 (
            .O(N__7995),
            .I(\U712_CHIP_RAM.CMA_5_0_8_cascade_ ));
    InMux I__1695 (
            .O(N__7992),
            .I(N__7989));
    LocalMux I__1694 (
            .O(N__7989),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    InMux I__1693 (
            .O(N__7986),
            .I(N__7983));
    LocalMux I__1692 (
            .O(N__7983),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i ));
    InMux I__1691 (
            .O(N__7980),
            .I(N__7977));
    LocalMux I__1690 (
            .O(N__7977),
            .I(N__7974));
    Span4Mux_v I__1689 (
            .O(N__7974),
            .I(N__7971));
    Sp12to4 I__1688 (
            .O(N__7971),
            .I(N__7968));
    Span12Mux_h I__1687 (
            .O(N__7968),
            .I(N__7965));
    Span12Mux_v I__1686 (
            .O(N__7965),
            .I(N__7962));
    Odrv12 I__1685 (
            .O(N__7962),
            .I(A_c_15));
    InMux I__1684 (
            .O(N__7959),
            .I(N__7956));
    LocalMux I__1683 (
            .O(N__7956),
            .I(N__7953));
    Span4Mux_v I__1682 (
            .O(N__7953),
            .I(N__7950));
    Sp12to4 I__1681 (
            .O(N__7950),
            .I(N__7947));
    Span12Mux_h I__1680 (
            .O(N__7947),
            .I(N__7944));
    Odrv12 I__1679 (
            .O(N__7944),
            .I(A_c_8));
    InMux I__1678 (
            .O(N__7941),
            .I(N__7938));
    LocalMux I__1677 (
            .O(N__7938),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__1676 (
            .O(N__7935),
            .I(N__7932));
    LocalMux I__1675 (
            .O(N__7932),
            .I(N__7929));
    Span12Mux_s3_v I__1674 (
            .O(N__7929),
            .I(N__7926));
    Span12Mux_v I__1673 (
            .O(N__7926),
            .I(N__7923));
    Odrv12 I__1672 (
            .O(N__7923),
            .I(CMA_c_0));
    InMux I__1671 (
            .O(N__7920),
            .I(N__7917));
    LocalMux I__1670 (
            .O(N__7917),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__1669 (
            .O(N__7914),
            .I(N__7911));
    LocalMux I__1668 (
            .O(N__7911),
            .I(N__7908));
    IoSpan4Mux I__1667 (
            .O(N__7908),
            .I(N__7905));
    Span4Mux_s2_h I__1666 (
            .O(N__7905),
            .I(N__7902));
    Sp12to4 I__1665 (
            .O(N__7902),
            .I(N__7899));
    Span12Mux_h I__1664 (
            .O(N__7899),
            .I(N__7896));
    Odrv12 I__1663 (
            .O(N__7896),
            .I(CMA_c_7));
    InMux I__1662 (
            .O(N__7893),
            .I(N__7890));
    LocalMux I__1661 (
            .O(N__7890),
            .I(\U712_CHIP_RAM.CLK_EN_6_0_a5_2 ));
    InMux I__1660 (
            .O(N__7887),
            .I(N__7884));
    LocalMux I__1659 (
            .O(N__7884),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_0 ));
    IoInMux I__1658 (
            .O(N__7881),
            .I(N__7878));
    LocalMux I__1657 (
            .O(N__7878),
            .I(N__7875));
    IoSpan4Mux I__1656 (
            .O(N__7875),
            .I(N__7872));
    IoSpan4Mux I__1655 (
            .O(N__7872),
            .I(N__7869));
    Span4Mux_s2_h I__1654 (
            .O(N__7869),
            .I(N__7866));
    Sp12to4 I__1653 (
            .O(N__7866),
            .I(N__7863));
    Span12Mux_h I__1652 (
            .O(N__7863),
            .I(N__7859));
    InMux I__1651 (
            .O(N__7862),
            .I(N__7856));
    Odrv12 I__1650 (
            .O(N__7859),
            .I(CLK_EN_c));
    LocalMux I__1649 (
            .O(N__7856),
            .I(CLK_EN_c));
    InMux I__1648 (
            .O(N__7851),
            .I(N__7848));
    LocalMux I__1647 (
            .O(N__7848),
            .I(N__7845));
    Odrv4 I__1646 (
            .O(N__7845),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__1645 (
            .O(N__7842),
            .I(N__7839));
    LocalMux I__1644 (
            .O(N__7839),
            .I(N__7835));
    InMux I__1643 (
            .O(N__7838),
            .I(N__7832));
    Span4Mux_v I__1642 (
            .O(N__7835),
            .I(N__7829));
    LocalMux I__1641 (
            .O(N__7832),
            .I(N__7826));
    Span4Mux_h I__1640 (
            .O(N__7829),
            .I(N__7823));
    Span4Mux_v I__1639 (
            .O(N__7826),
            .I(N__7820));
    Span4Mux_v I__1638 (
            .O(N__7823),
            .I(N__7816));
    Span4Mux_h I__1637 (
            .O(N__7820),
            .I(N__7813));
    InMux I__1636 (
            .O(N__7819),
            .I(N__7810));
    Odrv4 I__1635 (
            .O(N__7816),
            .I(DS_ENm));
    Odrv4 I__1634 (
            .O(N__7813),
            .I(DS_ENm));
    LocalMux I__1633 (
            .O(N__7810),
            .I(DS_ENm));
    IoInMux I__1632 (
            .O(N__7803),
            .I(N__7800));
    LocalMux I__1631 (
            .O(N__7800),
            .I(N__7797));
    Span4Mux_s2_v I__1630 (
            .O(N__7797),
            .I(N__7794));
    Span4Mux_h I__1629 (
            .O(N__7794),
            .I(N__7791));
    Span4Mux_h I__1628 (
            .O(N__7791),
            .I(N__7788));
    Span4Mux_v I__1627 (
            .O(N__7788),
            .I(N__7785));
    Odrv4 I__1626 (
            .O(N__7785),
            .I(U712_BYTE_ENABLE_un1_UDSn_i));
    InMux I__1625 (
            .O(N__7782),
            .I(N__7774));
    InMux I__1624 (
            .O(N__7781),
            .I(N__7771));
    InMux I__1623 (
            .O(N__7780),
            .I(N__7768));
    InMux I__1622 (
            .O(N__7779),
            .I(N__7765));
    InMux I__1621 (
            .O(N__7778),
            .I(N__7762));
    InMux I__1620 (
            .O(N__7777),
            .I(N__7759));
    LocalMux I__1619 (
            .O(N__7774),
            .I(N__7736));
    LocalMux I__1618 (
            .O(N__7771),
            .I(N__7736));
    LocalMux I__1617 (
            .O(N__7768),
            .I(N__7729));
    LocalMux I__1616 (
            .O(N__7765),
            .I(N__7729));
    LocalMux I__1615 (
            .O(N__7762),
            .I(N__7729));
    LocalMux I__1614 (
            .O(N__7759),
            .I(N__7726));
    InMux I__1613 (
            .O(N__7758),
            .I(N__7721));
    InMux I__1612 (
            .O(N__7757),
            .I(N__7721));
    InMux I__1611 (
            .O(N__7756),
            .I(N__7718));
    InMux I__1610 (
            .O(N__7755),
            .I(N__7715));
    InMux I__1609 (
            .O(N__7754),
            .I(N__7712));
    InMux I__1608 (
            .O(N__7753),
            .I(N__7709));
    InMux I__1607 (
            .O(N__7752),
            .I(N__7706));
    InMux I__1606 (
            .O(N__7751),
            .I(N__7699));
    InMux I__1605 (
            .O(N__7750),
            .I(N__7699));
    InMux I__1604 (
            .O(N__7749),
            .I(N__7699));
    InMux I__1603 (
            .O(N__7748),
            .I(N__7696));
    InMux I__1602 (
            .O(N__7747),
            .I(N__7693));
    InMux I__1601 (
            .O(N__7746),
            .I(N__7684));
    InMux I__1600 (
            .O(N__7745),
            .I(N__7684));
    InMux I__1599 (
            .O(N__7744),
            .I(N__7684));
    InMux I__1598 (
            .O(N__7743),
            .I(N__7684));
    InMux I__1597 (
            .O(N__7742),
            .I(N__7681));
    InMux I__1596 (
            .O(N__7741),
            .I(N__7678));
    Span4Mux_v I__1595 (
            .O(N__7736),
            .I(N__7673));
    Span4Mux_v I__1594 (
            .O(N__7729),
            .I(N__7673));
    Span4Mux_v I__1593 (
            .O(N__7726),
            .I(N__7660));
    LocalMux I__1592 (
            .O(N__7721),
            .I(N__7660));
    LocalMux I__1591 (
            .O(N__7718),
            .I(N__7660));
    LocalMux I__1590 (
            .O(N__7715),
            .I(N__7660));
    LocalMux I__1589 (
            .O(N__7712),
            .I(N__7660));
    LocalMux I__1588 (
            .O(N__7709),
            .I(N__7660));
    LocalMux I__1587 (
            .O(N__7706),
            .I(N__7657));
    LocalMux I__1586 (
            .O(N__7699),
            .I(N__7654));
    LocalMux I__1585 (
            .O(N__7696),
            .I(N__7647));
    LocalMux I__1584 (
            .O(N__7693),
            .I(N__7647));
    LocalMux I__1583 (
            .O(N__7684),
            .I(N__7647));
    LocalMux I__1582 (
            .O(N__7681),
            .I(N__7641));
    LocalMux I__1581 (
            .O(N__7678),
            .I(N__7638));
    Span4Mux_h I__1580 (
            .O(N__7673),
            .I(N__7631));
    Span4Mux_v I__1579 (
            .O(N__7660),
            .I(N__7631));
    Span4Mux_v I__1578 (
            .O(N__7657),
            .I(N__7631));
    Span4Mux_v I__1577 (
            .O(N__7654),
            .I(N__7626));
    Span4Mux_v I__1576 (
            .O(N__7647),
            .I(N__7626));
    InMux I__1575 (
            .O(N__7646),
            .I(N__7623));
    InMux I__1574 (
            .O(N__7645),
            .I(N__7620));
    InMux I__1573 (
            .O(N__7644),
            .I(N__7617));
    Span12Mux_v I__1572 (
            .O(N__7641),
            .I(N__7610));
    Span12Mux_h I__1571 (
            .O(N__7638),
            .I(N__7610));
    Sp12to4 I__1570 (
            .O(N__7631),
            .I(N__7610));
    Sp12to4 I__1569 (
            .O(N__7626),
            .I(N__7601));
    LocalMux I__1568 (
            .O(N__7623),
            .I(N__7601));
    LocalMux I__1567 (
            .O(N__7620),
            .I(N__7601));
    LocalMux I__1566 (
            .O(N__7617),
            .I(N__7601));
    Span12Mux_h I__1565 (
            .O(N__7610),
            .I(N__7598));
    Span12Mux_h I__1564 (
            .O(N__7601),
            .I(N__7595));
    Odrv12 I__1563 (
            .O(N__7598),
            .I(RESETn_c));
    Odrv12 I__1562 (
            .O(N__7595),
            .I(RESETn_c));
    IoInMux I__1561 (
            .O(N__7590),
            .I(N__7587));
    LocalMux I__1560 (
            .O(N__7587),
            .I(N__7584));
    Span12Mux_s2_v I__1559 (
            .O(N__7584),
            .I(N__7581));
    Odrv12 I__1558 (
            .O(N__7581),
            .I(RESETn_c_i));
    IoInMux I__1557 (
            .O(N__7578),
            .I(N__7575));
    LocalMux I__1556 (
            .O(N__7575),
            .I(N__7572));
    Span12Mux_s11_v I__1555 (
            .O(N__7572),
            .I(N__7569));
    Span12Mux_h I__1554 (
            .O(N__7569),
            .I(N__7566));
    Odrv12 I__1553 (
            .O(N__7566),
            .I(N_163));
    InMux I__1552 (
            .O(N__7563),
            .I(N__7560));
    LocalMux I__1551 (
            .O(N__7560),
            .I(N__7557));
    Span4Mux_v I__1550 (
            .O(N__7557),
            .I(N__7554));
    Span4Mux_v I__1549 (
            .O(N__7554),
            .I(N__7551));
    Sp12to4 I__1548 (
            .O(N__7551),
            .I(N__7548));
    Span12Mux_h I__1547 (
            .O(N__7548),
            .I(N__7545));
    Odrv12 I__1546 (
            .O(N__7545),
            .I(A_c_17));
    IoInMux I__1545 (
            .O(N__7542),
            .I(N__7539));
    LocalMux I__1544 (
            .O(N__7539),
            .I(N__7536));
    Span12Mux_s3_h I__1543 (
            .O(N__7536),
            .I(N__7533));
    Span12Mux_h I__1542 (
            .O(N__7533),
            .I(N__7530));
    Odrv12 I__1541 (
            .O(N__7530),
            .I(CMA_c_8));
    CascadeMux I__1540 (
            .O(N__7527),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ));
    InMux I__1539 (
            .O(N__7524),
            .I(N__7521));
    LocalMux I__1538 (
            .O(N__7521),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    InMux I__1537 (
            .O(N__7518),
            .I(N__7515));
    LocalMux I__1536 (
            .O(N__7515),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    InMux I__1535 (
            .O(N__7512),
            .I(N__7509));
    LocalMux I__1534 (
            .O(N__7509),
            .I(N__7506));
    Odrv4 I__1533 (
            .O(N__7506),
            .I(\U712_CHIP_RAM.N_146 ));
    CascadeMux I__1532 (
            .O(N__7503),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5_cascade_ ));
    IoInMux I__1531 (
            .O(N__7500),
            .I(N__7497));
    LocalMux I__1530 (
            .O(N__7497),
            .I(N__7494));
    Span4Mux_s3_h I__1529 (
            .O(N__7494),
            .I(N__7491));
    Sp12to4 I__1528 (
            .O(N__7491),
            .I(N__7488));
    Span12Mux_s8_v I__1527 (
            .O(N__7488),
            .I(N__7485));
    Span12Mux_h I__1526 (
            .O(N__7485),
            .I(N__7482));
    Odrv12 I__1525 (
            .O(N__7482),
            .I(CMA_c_5));
    InMux I__1524 (
            .O(N__7479),
            .I(N__7476));
    LocalMux I__1523 (
            .O(N__7476),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    CascadeMux I__1522 (
            .O(N__7473),
            .I(N__7468));
    InMux I__1521 (
            .O(N__7472),
            .I(N__7465));
    InMux I__1520 (
            .O(N__7471),
            .I(N__7462));
    InMux I__1519 (
            .O(N__7468),
            .I(N__7459));
    LocalMux I__1518 (
            .O(N__7465),
            .I(N__7454));
    LocalMux I__1517 (
            .O(N__7462),
            .I(N__7454));
    LocalMux I__1516 (
            .O(N__7459),
            .I(REG_TACK));
    Odrv12 I__1515 (
            .O(N__7454),
            .I(REG_TACK));
    InMux I__1514 (
            .O(N__7449),
            .I(N__7445));
    InMux I__1513 (
            .O(N__7448),
            .I(N__7441));
    LocalMux I__1512 (
            .O(N__7445),
            .I(N__7438));
    InMux I__1511 (
            .O(N__7444),
            .I(N__7435));
    LocalMux I__1510 (
            .O(N__7441),
            .I(N__7432));
    Span4Mux_h I__1509 (
            .O(N__7438),
            .I(N__7427));
    LocalMux I__1508 (
            .O(N__7435),
            .I(N__7427));
    Odrv12 I__1507 (
            .O(N__7432),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    Odrv4 I__1506 (
            .O(N__7427),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    InMux I__1505 (
            .O(N__7422),
            .I(N__7416));
    InMux I__1504 (
            .O(N__7421),
            .I(N__7413));
    InMux I__1503 (
            .O(N__7420),
            .I(N__7409));
    InMux I__1502 (
            .O(N__7419),
            .I(N__7406));
    LocalMux I__1501 (
            .O(N__7416),
            .I(N__7399));
    LocalMux I__1500 (
            .O(N__7413),
            .I(N__7399));
    InMux I__1499 (
            .O(N__7412),
            .I(N__7396));
    LocalMux I__1498 (
            .O(N__7409),
            .I(N__7393));
    LocalMux I__1497 (
            .O(N__7406),
            .I(N__7389));
    InMux I__1496 (
            .O(N__7405),
            .I(N__7384));
    InMux I__1495 (
            .O(N__7404),
            .I(N__7384));
    Span4Mux_v I__1494 (
            .O(N__7399),
            .I(N__7379));
    LocalMux I__1493 (
            .O(N__7396),
            .I(N__7379));
    Span4Mux_h I__1492 (
            .O(N__7393),
            .I(N__7376));
    InMux I__1491 (
            .O(N__7392),
            .I(N__7373));
    Odrv12 I__1490 (
            .O(N__7389),
            .I(WRITE_CYCLEm));
    LocalMux I__1489 (
            .O(N__7384),
            .I(WRITE_CYCLEm));
    Odrv4 I__1488 (
            .O(N__7379),
            .I(WRITE_CYCLEm));
    Odrv4 I__1487 (
            .O(N__7376),
            .I(WRITE_CYCLEm));
    LocalMux I__1486 (
            .O(N__7373),
            .I(WRITE_CYCLEm));
    CascadeMux I__1485 (
            .O(N__7362),
            .I(N__7359));
    InMux I__1484 (
            .O(N__7359),
            .I(N__7356));
    LocalMux I__1483 (
            .O(N__7356),
            .I(N__7353));
    Span4Mux_h I__1482 (
            .O(N__7353),
            .I(N__7349));
    InMux I__1481 (
            .O(N__7352),
            .I(N__7346));
    Odrv4 I__1480 (
            .O(N__7349),
            .I(CPU_TACKm));
    LocalMux I__1479 (
            .O(N__7346),
            .I(CPU_TACKm));
    CEMux I__1478 (
            .O(N__7341),
            .I(N__7338));
    LocalMux I__1477 (
            .O(N__7338),
            .I(N__7335));
    Odrv4 I__1476 (
            .O(N__7335),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0 ));
    IoInMux I__1475 (
            .O(N__7332),
            .I(N__7329));
    LocalMux I__1474 (
            .O(N__7329),
            .I(N__7326));
    IoSpan4Mux I__1473 (
            .O(N__7326),
            .I(N__7323));
    Span4Mux_s3_h I__1472 (
            .O(N__7323),
            .I(N__7320));
    Sp12to4 I__1471 (
            .O(N__7320),
            .I(N__7317));
    Span12Mux_s8_h I__1470 (
            .O(N__7317),
            .I(N__7314));
    Span12Mux_v I__1469 (
            .O(N__7314),
            .I(N__7311));
    Odrv12 I__1468 (
            .O(N__7311),
            .I(N_118_i));
    IoInMux I__1467 (
            .O(N__7308),
            .I(N__7305));
    LocalMux I__1466 (
            .O(N__7305),
            .I(N__7302));
    Span4Mux_s0_h I__1465 (
            .O(N__7302),
            .I(N__7299));
    Sp12to4 I__1464 (
            .O(N__7299),
            .I(N__7296));
    Span12Mux_s6_v I__1463 (
            .O(N__7296),
            .I(N__7293));
    Span12Mux_h I__1462 (
            .O(N__7293),
            .I(N__7290));
    Span12Mux_v I__1461 (
            .O(N__7290),
            .I(N__7287));
    Odrv12 I__1460 (
            .O(N__7287),
            .I(N_119_i));
    InMux I__1459 (
            .O(N__7284),
            .I(N__7281));
    LocalMux I__1458 (
            .O(N__7281),
            .I(N__7277));
    InMux I__1457 (
            .O(N__7280),
            .I(N__7274));
    Span4Mux_h I__1456 (
            .O(N__7277),
            .I(N__7268));
    LocalMux I__1455 (
            .O(N__7274),
            .I(N__7265));
    InMux I__1454 (
            .O(N__7273),
            .I(N__7262));
    InMux I__1453 (
            .O(N__7272),
            .I(N__7257));
    InMux I__1452 (
            .O(N__7271),
            .I(N__7257));
    Odrv4 I__1451 (
            .O(N__7268),
            .I(\U712_CHIP_RAM.N_323 ));
    Odrv4 I__1450 (
            .O(N__7265),
            .I(\U712_CHIP_RAM.N_323 ));
    LocalMux I__1449 (
            .O(N__7262),
            .I(\U712_CHIP_RAM.N_323 ));
    LocalMux I__1448 (
            .O(N__7257),
            .I(\U712_CHIP_RAM.N_323 ));
    InMux I__1447 (
            .O(N__7248),
            .I(N__7242));
    CascadeMux I__1446 (
            .O(N__7247),
            .I(N__7238));
    InMux I__1445 (
            .O(N__7246),
            .I(N__7230));
    InMux I__1444 (
            .O(N__7245),
            .I(N__7230));
    LocalMux I__1443 (
            .O(N__7242),
            .I(N__7226));
    InMux I__1442 (
            .O(N__7241),
            .I(N__7218));
    InMux I__1441 (
            .O(N__7238),
            .I(N__7218));
    CascadeMux I__1440 (
            .O(N__7237),
            .I(N__7213));
    InMux I__1439 (
            .O(N__7236),
            .I(N__7210));
    InMux I__1438 (
            .O(N__7235),
            .I(N__7207));
    LocalMux I__1437 (
            .O(N__7230),
            .I(N__7204));
    InMux I__1436 (
            .O(N__7229),
            .I(N__7201));
    Span4Mux_h I__1435 (
            .O(N__7226),
            .I(N__7198));
    InMux I__1434 (
            .O(N__7225),
            .I(N__7191));
    InMux I__1433 (
            .O(N__7224),
            .I(N__7191));
    InMux I__1432 (
            .O(N__7223),
            .I(N__7191));
    LocalMux I__1431 (
            .O(N__7218),
            .I(N__7188));
    InMux I__1430 (
            .O(N__7217),
            .I(N__7183));
    InMux I__1429 (
            .O(N__7216),
            .I(N__7183));
    InMux I__1428 (
            .O(N__7213),
            .I(N__7180));
    LocalMux I__1427 (
            .O(N__7210),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1426 (
            .O(N__7207),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1425 (
            .O(N__7204),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1424 (
            .O(N__7201),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1423 (
            .O(N__7198),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1422 (
            .O(N__7191),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1421 (
            .O(N__7188),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1420 (
            .O(N__7183),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1419 (
            .O(N__7180),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__1418 (
            .O(N__7161),
            .I(N__7156));
    InMux I__1417 (
            .O(N__7160),
            .I(N__7152));
    InMux I__1416 (
            .O(N__7159),
            .I(N__7149));
    InMux I__1415 (
            .O(N__7156),
            .I(N__7142));
    CascadeMux I__1414 (
            .O(N__7155),
            .I(N__7138));
    LocalMux I__1413 (
            .O(N__7152),
            .I(N__7135));
    LocalMux I__1412 (
            .O(N__7149),
            .I(N__7132));
    InMux I__1411 (
            .O(N__7148),
            .I(N__7127));
    InMux I__1410 (
            .O(N__7147),
            .I(N__7127));
    CascadeMux I__1409 (
            .O(N__7146),
            .I(N__7124));
    InMux I__1408 (
            .O(N__7145),
            .I(N__7118));
    LocalMux I__1407 (
            .O(N__7142),
            .I(N__7115));
    InMux I__1406 (
            .O(N__7141),
            .I(N__7112));
    InMux I__1405 (
            .O(N__7138),
            .I(N__7109));
    Span4Mux_v I__1404 (
            .O(N__7135),
            .I(N__7102));
    Span4Mux_v I__1403 (
            .O(N__7132),
            .I(N__7102));
    LocalMux I__1402 (
            .O(N__7127),
            .I(N__7102));
    InMux I__1401 (
            .O(N__7124),
            .I(N__7097));
    InMux I__1400 (
            .O(N__7123),
            .I(N__7097));
    InMux I__1399 (
            .O(N__7122),
            .I(N__7094));
    InMux I__1398 (
            .O(N__7121),
            .I(N__7091));
    LocalMux I__1397 (
            .O(N__7118),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1396 (
            .O(N__7115),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1395 (
            .O(N__7112),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1394 (
            .O(N__7109),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1393 (
            .O(N__7102),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1392 (
            .O(N__7097),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1391 (
            .O(N__7094),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1390 (
            .O(N__7091),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1389 (
            .O(N__7074),
            .I(N__7071));
    LocalMux I__1388 (
            .O(N__7071),
            .I(\U712_CHIP_RAM.CPU_TACK_7_iv_i_a5_0_1_0 ));
    CascadeMux I__1387 (
            .O(N__7068),
            .I(N__7065));
    InMux I__1386 (
            .O(N__7065),
            .I(N__7062));
    LocalMux I__1385 (
            .O(N__7062),
            .I(\U712_CHIP_RAM.N_287 ));
    InMux I__1384 (
            .O(N__7059),
            .I(N__7053));
    InMux I__1383 (
            .O(N__7058),
            .I(N__7050));
    InMux I__1382 (
            .O(N__7057),
            .I(N__7047));
    InMux I__1381 (
            .O(N__7056),
            .I(N__7044));
    LocalMux I__1380 (
            .O(N__7053),
            .I(N__7041));
    LocalMux I__1379 (
            .O(N__7050),
            .I(N__7038));
    LocalMux I__1378 (
            .O(N__7047),
            .I(N__7033));
    LocalMux I__1377 (
            .O(N__7044),
            .I(N__7030));
    Span4Mux_v I__1376 (
            .O(N__7041),
            .I(N__7024));
    Span4Mux_v I__1375 (
            .O(N__7038),
            .I(N__7024));
    InMux I__1374 (
            .O(N__7037),
            .I(N__7019));
    InMux I__1373 (
            .O(N__7036),
            .I(N__7019));
    Span4Mux_v I__1372 (
            .O(N__7033),
            .I(N__7014));
    Span4Mux_v I__1371 (
            .O(N__7030),
            .I(N__7014));
    InMux I__1370 (
            .O(N__7029),
            .I(N__7011));
    Odrv4 I__1369 (
            .O(N__7024),
            .I(DMA_CYCLEm));
    LocalMux I__1368 (
            .O(N__7019),
            .I(DMA_CYCLEm));
    Odrv4 I__1367 (
            .O(N__7014),
            .I(DMA_CYCLEm));
    LocalMux I__1366 (
            .O(N__7011),
            .I(DMA_CYCLEm));
    IoInMux I__1365 (
            .O(N__7002),
            .I(N__6999));
    LocalMux I__1364 (
            .O(N__6999),
            .I(N__6995));
    InMux I__1363 (
            .O(N__6998),
            .I(N__6992));
    Span12Mux_s4_v I__1362 (
            .O(N__6995),
            .I(N__6989));
    LocalMux I__1361 (
            .O(N__6992),
            .I(N__6986));
    Span12Mux_v I__1360 (
            .O(N__6989),
            .I(N__6981));
    Span4Mux_v I__1359 (
            .O(N__6986),
            .I(N__6978));
    InMux I__1358 (
            .O(N__6985),
            .I(N__6975));
    InMux I__1357 (
            .O(N__6984),
            .I(N__6972));
    Odrv12 I__1356 (
            .O(N__6981),
            .I(DBENn_c));
    Odrv4 I__1355 (
            .O(N__6978),
            .I(DBENn_c));
    LocalMux I__1354 (
            .O(N__6975),
            .I(DBENn_c));
    LocalMux I__1353 (
            .O(N__6972),
            .I(DBENn_c));
    InMux I__1352 (
            .O(N__6963),
            .I(N__6957));
    InMux I__1351 (
            .O(N__6962),
            .I(N__6957));
    LocalMux I__1350 (
            .O(N__6957),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a5_0Z0Z_0 ));
    CascadeMux I__1349 (
            .O(N__6954),
            .I(N__6951));
    InMux I__1348 (
            .O(N__6951),
            .I(N__6948));
    LocalMux I__1347 (
            .O(N__6948),
            .I(N__6945));
    Odrv4 I__1346 (
            .O(N__6945),
            .I(\U712_BYTE_ENABLE.UUBE ));
    InMux I__1345 (
            .O(N__6942),
            .I(N__6939));
    LocalMux I__1344 (
            .O(N__6939),
            .I(N__6936));
    Odrv4 I__1343 (
            .O(N__6936),
            .I(\U712_BYTE_ENABLE.N_216 ));
    CascadeMux I__1342 (
            .O(N__6933),
            .I(N__6930));
    InMux I__1341 (
            .O(N__6930),
            .I(N__6927));
    LocalMux I__1340 (
            .O(N__6927),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    InMux I__1339 (
            .O(N__6924),
            .I(N__6921));
    LocalMux I__1338 (
            .O(N__6921),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    InMux I__1337 (
            .O(N__6918),
            .I(N__6915));
    LocalMux I__1336 (
            .O(N__6915),
            .I(N__6912));
    Span12Mux_h I__1335 (
            .O(N__6912),
            .I(N__6909));
    Odrv12 I__1334 (
            .O(N__6909),
            .I(A_c_9));
    InMux I__1333 (
            .O(N__6906),
            .I(N__6903));
    LocalMux I__1332 (
            .O(N__6903),
            .I(N__6900));
    Span12Mux_v I__1331 (
            .O(N__6900),
            .I(N__6897));
    Span12Mux_h I__1330 (
            .O(N__6897),
            .I(N__6894));
    Odrv12 I__1329 (
            .O(N__6894),
            .I(A_c_2));
    CascadeMux I__1328 (
            .O(N__6891),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ));
    InMux I__1327 (
            .O(N__6888),
            .I(N__6885));
    LocalMux I__1326 (
            .O(N__6885),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__1325 (
            .O(N__6882),
            .I(N__6879));
    LocalMux I__1324 (
            .O(N__6879),
            .I(N__6876));
    Span12Mux_v I__1323 (
            .O(N__6876),
            .I(N__6873));
    Span12Mux_h I__1322 (
            .O(N__6873),
            .I(N__6870));
    Odrv12 I__1321 (
            .O(N__6870),
            .I(A_c_7));
    InMux I__1320 (
            .O(N__6867),
            .I(N__6862));
    CascadeMux I__1319 (
            .O(N__6866),
            .I(N__6859));
    InMux I__1318 (
            .O(N__6865),
            .I(N__6856));
    LocalMux I__1317 (
            .O(N__6862),
            .I(N__6853));
    InMux I__1316 (
            .O(N__6859),
            .I(N__6850));
    LocalMux I__1315 (
            .O(N__6856),
            .I(N__6846));
    Span4Mux_h I__1314 (
            .O(N__6853),
            .I(N__6841));
    LocalMux I__1313 (
            .O(N__6850),
            .I(N__6841));
    InMux I__1312 (
            .O(N__6849),
            .I(N__6838));
    Span4Mux_v I__1311 (
            .O(N__6846),
            .I(N__6833));
    Span4Mux_h I__1310 (
            .O(N__6841),
            .I(N__6833));
    LocalMux I__1309 (
            .O(N__6838),
            .I(N__6830));
    Span4Mux_v I__1308 (
            .O(N__6833),
            .I(N__6827));
    Span12Mux_h I__1307 (
            .O(N__6830),
            .I(N__6824));
    Span4Mux_v I__1306 (
            .O(N__6827),
            .I(N__6821));
    Span12Mux_v I__1305 (
            .O(N__6824),
            .I(N__6818));
    Span4Mux_v I__1304 (
            .O(N__6821),
            .I(N__6815));
    Odrv12 I__1303 (
            .O(N__6818),
            .I(CLK40_PLL_i));
    Odrv4 I__1302 (
            .O(N__6815),
            .I(CLK40_PLL_i));
    IoInMux I__1301 (
            .O(N__6810),
            .I(N__6807));
    LocalMux I__1300 (
            .O(N__6807),
            .I(N__6802));
    IoInMux I__1299 (
            .O(N__6806),
            .I(N__6799));
    IoInMux I__1298 (
            .O(N__6805),
            .I(N__6796));
    Span4Mux_s1_v I__1297 (
            .O(N__6802),
            .I(N__6793));
    LocalMux I__1296 (
            .O(N__6799),
            .I(N__6790));
    LocalMux I__1295 (
            .O(N__6796),
            .I(N__6787));
    Span4Mux_h I__1294 (
            .O(N__6793),
            .I(N__6784));
    Span4Mux_s1_v I__1293 (
            .O(N__6790),
            .I(N__6781));
    Span4Mux_s3_h I__1292 (
            .O(N__6787),
            .I(N__6778));
    Sp12to4 I__1291 (
            .O(N__6784),
            .I(N__6773));
    Sp12to4 I__1290 (
            .O(N__6781),
            .I(N__6773));
    Span4Mux_h I__1289 (
            .O(N__6778),
            .I(N__6770));
    Span12Mux_h I__1288 (
            .O(N__6773),
            .I(N__6767));
    Span4Mux_h I__1287 (
            .O(N__6770),
            .I(N__6764));
    Span12Mux_v I__1286 (
            .O(N__6767),
            .I(N__6761));
    Span4Mux_h I__1285 (
            .O(N__6764),
            .I(N__6758));
    Odrv12 I__1284 (
            .O(N__6761),
            .I(CLK40_PLL_i_i));
    Odrv4 I__1283 (
            .O(N__6758),
            .I(CLK40_PLL_i_i));
    InMux I__1282 (
            .O(N__6753),
            .I(N__6750));
    LocalMux I__1281 (
            .O(N__6750),
            .I(N__6744));
    InMux I__1280 (
            .O(N__6749),
            .I(N__6741));
    InMux I__1279 (
            .O(N__6748),
            .I(N__6734));
    InMux I__1278 (
            .O(N__6747),
            .I(N__6731));
    Span4Mux_h I__1277 (
            .O(N__6744),
            .I(N__6726));
    LocalMux I__1276 (
            .O(N__6741),
            .I(N__6726));
    InMux I__1275 (
            .O(N__6740),
            .I(N__6723));
    InMux I__1274 (
            .O(N__6739),
            .I(N__6720));
    InMux I__1273 (
            .O(N__6738),
            .I(N__6715));
    InMux I__1272 (
            .O(N__6737),
            .I(N__6715));
    LocalMux I__1271 (
            .O(N__6734),
            .I(\U712_CHIP_RAM.N_327 ));
    LocalMux I__1270 (
            .O(N__6731),
            .I(\U712_CHIP_RAM.N_327 ));
    Odrv4 I__1269 (
            .O(N__6726),
            .I(\U712_CHIP_RAM.N_327 ));
    LocalMux I__1268 (
            .O(N__6723),
            .I(\U712_CHIP_RAM.N_327 ));
    LocalMux I__1267 (
            .O(N__6720),
            .I(\U712_CHIP_RAM.N_327 ));
    LocalMux I__1266 (
            .O(N__6715),
            .I(\U712_CHIP_RAM.N_327 ));
    InMux I__1265 (
            .O(N__6702),
            .I(N__6697));
    InMux I__1264 (
            .O(N__6701),
            .I(N__6694));
    InMux I__1263 (
            .O(N__6700),
            .I(N__6691));
    LocalMux I__1262 (
            .O(N__6697),
            .I(\U712_CHIP_RAM.N_339 ));
    LocalMux I__1261 (
            .O(N__6694),
            .I(\U712_CHIP_RAM.N_339 ));
    LocalMux I__1260 (
            .O(N__6691),
            .I(\U712_CHIP_RAM.N_339 ));
    CascadeMux I__1259 (
            .O(N__6684),
            .I(N__6680));
    CascadeMux I__1258 (
            .O(N__6683),
            .I(N__6677));
    InMux I__1257 (
            .O(N__6680),
            .I(N__6669));
    InMux I__1256 (
            .O(N__6677),
            .I(N__6669));
    InMux I__1255 (
            .O(N__6676),
            .I(N__6664));
    InMux I__1254 (
            .O(N__6675),
            .I(N__6664));
    CascadeMux I__1253 (
            .O(N__6674),
            .I(N__6658));
    LocalMux I__1252 (
            .O(N__6669),
            .I(N__6651));
    LocalMux I__1251 (
            .O(N__6664),
            .I(N__6651));
    InMux I__1250 (
            .O(N__6663),
            .I(N__6646));
    CascadeMux I__1249 (
            .O(N__6662),
            .I(N__6642));
    InMux I__1248 (
            .O(N__6661),
            .I(N__6636));
    InMux I__1247 (
            .O(N__6658),
            .I(N__6636));
    InMux I__1246 (
            .O(N__6657),
            .I(N__6630));
    InMux I__1245 (
            .O(N__6656),
            .I(N__6627));
    Span4Mux_v I__1244 (
            .O(N__6651),
            .I(N__6624));
    InMux I__1243 (
            .O(N__6650),
            .I(N__6619));
    InMux I__1242 (
            .O(N__6649),
            .I(N__6619));
    LocalMux I__1241 (
            .O(N__6646),
            .I(N__6616));
    InMux I__1240 (
            .O(N__6645),
            .I(N__6613));
    InMux I__1239 (
            .O(N__6642),
            .I(N__6608));
    InMux I__1238 (
            .O(N__6641),
            .I(N__6608));
    LocalMux I__1237 (
            .O(N__6636),
            .I(N__6605));
    InMux I__1236 (
            .O(N__6635),
            .I(N__6600));
    InMux I__1235 (
            .O(N__6634),
            .I(N__6600));
    InMux I__1234 (
            .O(N__6633),
            .I(N__6597));
    LocalMux I__1233 (
            .O(N__6630),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1232 (
            .O(N__6627),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1231 (
            .O(N__6624),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1230 (
            .O(N__6619),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1229 (
            .O(N__6616),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1228 (
            .O(N__6613),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1227 (
            .O(N__6608),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv12 I__1226 (
            .O(N__6605),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1225 (
            .O(N__6600),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1224 (
            .O(N__6597),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    CascadeMux I__1223 (
            .O(N__6576),
            .I(N__6568));
    CascadeMux I__1222 (
            .O(N__6575),
            .I(N__6565));
    CascadeMux I__1221 (
            .O(N__6574),
            .I(N__6558));
    CascadeMux I__1220 (
            .O(N__6573),
            .I(N__6555));
    InMux I__1219 (
            .O(N__6572),
            .I(N__6551));
    InMux I__1218 (
            .O(N__6571),
            .I(N__6542));
    InMux I__1217 (
            .O(N__6568),
            .I(N__6542));
    InMux I__1216 (
            .O(N__6565),
            .I(N__6542));
    InMux I__1215 (
            .O(N__6564),
            .I(N__6539));
    InMux I__1214 (
            .O(N__6563),
            .I(N__6535));
    InMux I__1213 (
            .O(N__6562),
            .I(N__6530));
    InMux I__1212 (
            .O(N__6561),
            .I(N__6530));
    InMux I__1211 (
            .O(N__6558),
            .I(N__6527));
    InMux I__1210 (
            .O(N__6555),
            .I(N__6524));
    InMux I__1209 (
            .O(N__6554),
            .I(N__6521));
    LocalMux I__1208 (
            .O(N__6551),
            .I(N__6518));
    InMux I__1207 (
            .O(N__6550),
            .I(N__6513));
    InMux I__1206 (
            .O(N__6549),
            .I(N__6513));
    LocalMux I__1205 (
            .O(N__6542),
            .I(N__6510));
    LocalMux I__1204 (
            .O(N__6539),
            .I(N__6507));
    InMux I__1203 (
            .O(N__6538),
            .I(N__6504));
    LocalMux I__1202 (
            .O(N__6535),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1201 (
            .O(N__6530),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1200 (
            .O(N__6527),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1199 (
            .O(N__6524),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1198 (
            .O(N__6521),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1197 (
            .O(N__6518),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1196 (
            .O(N__6513),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1195 (
            .O(N__6510),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1194 (
            .O(N__6507),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1193 (
            .O(N__6504),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    CascadeMux I__1192 (
            .O(N__6483),
            .I(N__6480));
    InMux I__1191 (
            .O(N__6480),
            .I(N__6477));
    LocalMux I__1190 (
            .O(N__6477),
            .I(\U712_CHIP_RAM.un3_DMA_CYCLE_START ));
    InMux I__1189 (
            .O(N__6474),
            .I(N__6471));
    LocalMux I__1188 (
            .O(N__6471),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__1187 (
            .O(N__6468),
            .I(N__6462));
    InMux I__1186 (
            .O(N__6467),
            .I(N__6462));
    LocalMux I__1185 (
            .O(N__6462),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    IoInMux I__1184 (
            .O(N__6459),
            .I(N__6456));
    LocalMux I__1183 (
            .O(N__6456),
            .I(N__6453));
    IoSpan4Mux I__1182 (
            .O(N__6453),
            .I(N__6450));
    Span4Mux_s3_v I__1181 (
            .O(N__6450),
            .I(N__6447));
    Span4Mux_v I__1180 (
            .O(N__6447),
            .I(N__6444));
    Odrv4 I__1179 (
            .O(N__6444),
            .I(CONSTANT_ONE_NET));
    InMux I__1178 (
            .O(N__6441),
            .I(N__6438));
    LocalMux I__1177 (
            .O(N__6438),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    IoInMux I__1176 (
            .O(N__6435),
            .I(N__6432));
    LocalMux I__1175 (
            .O(N__6432),
            .I(N__6429));
    Span12Mux_s5_v I__1174 (
            .O(N__6429),
            .I(N__6426));
    Odrv12 I__1173 (
            .O(N__6426),
            .I(CMA_c_1));
    InMux I__1172 (
            .O(N__6423),
            .I(N__6420));
    LocalMux I__1171 (
            .O(N__6420),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__1170 (
            .O(N__6417),
            .I(N__6414));
    LocalMux I__1169 (
            .O(N__6414),
            .I(N__6411));
    IoSpan4Mux I__1168 (
            .O(N__6411),
            .I(N__6408));
    Span4Mux_s3_v I__1167 (
            .O(N__6408),
            .I(N__6405));
    Sp12to4 I__1166 (
            .O(N__6405),
            .I(N__6402));
    Odrv12 I__1165 (
            .O(N__6402),
            .I(CMA_c_2));
    IoInMux I__1164 (
            .O(N__6399),
            .I(N__6396));
    LocalMux I__1163 (
            .O(N__6396),
            .I(N__6393));
    Span12Mux_s6_h I__1162 (
            .O(N__6393),
            .I(N__6390));
    Span12Mux_v I__1161 (
            .O(N__6390),
            .I(N__6387));
    Odrv12 I__1160 (
            .O(N__6387),
            .I(CMA_c_3));
    InMux I__1159 (
            .O(N__6384),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    CEMux I__1158 (
            .O(N__6381),
            .I(N__6378));
    LocalMux I__1157 (
            .O(N__6378),
            .I(N__6375));
    Span4Mux_v I__1156 (
            .O(N__6375),
            .I(N__6371));
    CEMux I__1155 (
            .O(N__6374),
            .I(N__6368));
    Span4Mux_h I__1154 (
            .O(N__6371),
            .I(N__6365));
    LocalMux I__1153 (
            .O(N__6368),
            .I(N__6362));
    Odrv4 I__1152 (
            .O(N__6365),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv4 I__1151 (
            .O(N__6362),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__1150 (
            .O(N__6357),
            .I(N__6354));
    LocalMux I__1149 (
            .O(N__6354),
            .I(N__6351));
    Span4Mux_v I__1148 (
            .O(N__6351),
            .I(N__6348));
    Sp12to4 I__1147 (
            .O(N__6348),
            .I(N__6345));
    Span12Mux_h I__1146 (
            .O(N__6345),
            .I(N__6342));
    Odrv12 I__1145 (
            .O(N__6342),
            .I(A_c_20));
    CascadeMux I__1144 (
            .O(N__6339),
            .I(\U712_CHIP_RAM.N_289_cascade_ ));
    InMux I__1143 (
            .O(N__6336),
            .I(N__6333));
    LocalMux I__1142 (
            .O(N__6333),
            .I(N__6330));
    Odrv4 I__1141 (
            .O(N__6330),
            .I(\U712_CHIP_RAM.N_288 ));
    IoInMux I__1140 (
            .O(N__6327),
            .I(N__6324));
    LocalMux I__1139 (
            .O(N__6324),
            .I(N__6321));
    IoSpan4Mux I__1138 (
            .O(N__6321),
            .I(N__6318));
    Sp12to4 I__1137 (
            .O(N__6318),
            .I(N__6315));
    Span12Mux_s7_v I__1136 (
            .O(N__6315),
            .I(N__6311));
    InMux I__1135 (
            .O(N__6314),
            .I(N__6308));
    Odrv12 I__1134 (
            .O(N__6311),
            .I(BANK0_c));
    LocalMux I__1133 (
            .O(N__6308),
            .I(BANK0_c));
    InMux I__1132 (
            .O(N__6303),
            .I(N__6299));
    InMux I__1131 (
            .O(N__6302),
            .I(N__6296));
    LocalMux I__1130 (
            .O(N__6299),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a5_0 ));
    LocalMux I__1129 (
            .O(N__6296),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a5_0 ));
    InMux I__1128 (
            .O(N__6291),
            .I(N__6287));
    CascadeMux I__1127 (
            .O(N__6290),
            .I(N__6283));
    LocalMux I__1126 (
            .O(N__6287),
            .I(N__6280));
    InMux I__1125 (
            .O(N__6286),
            .I(N__6277));
    InMux I__1124 (
            .O(N__6283),
            .I(N__6274));
    Odrv4 I__1123 (
            .O(N__6280),
            .I(\U712_CHIP_RAM.N_186 ));
    LocalMux I__1122 (
            .O(N__6277),
            .I(\U712_CHIP_RAM.N_186 ));
    LocalMux I__1121 (
            .O(N__6274),
            .I(\U712_CHIP_RAM.N_186 ));
    InMux I__1120 (
            .O(N__6267),
            .I(N__6264));
    LocalMux I__1119 (
            .O(N__6264),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0 ));
    InMux I__1118 (
            .O(N__6261),
            .I(N__6257));
    InMux I__1117 (
            .O(N__6260),
            .I(N__6254));
    LocalMux I__1116 (
            .O(N__6257),
            .I(N__6251));
    LocalMux I__1115 (
            .O(N__6254),
            .I(N__6247));
    Span4Mux_v I__1114 (
            .O(N__6251),
            .I(N__6244));
    InMux I__1113 (
            .O(N__6250),
            .I(N__6241));
    Span4Mux_h I__1112 (
            .O(N__6247),
            .I(N__6238));
    Odrv4 I__1111 (
            .O(N__6244),
            .I(\U712_CHIP_RAM.N_341 ));
    LocalMux I__1110 (
            .O(N__6241),
            .I(\U712_CHIP_RAM.N_341 ));
    Odrv4 I__1109 (
            .O(N__6238),
            .I(\U712_CHIP_RAM.N_341 ));
    InMux I__1108 (
            .O(N__6231),
            .I(N__6228));
    LocalMux I__1107 (
            .O(N__6228),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ));
    InMux I__1106 (
            .O(N__6225),
            .I(N__6222));
    LocalMux I__1105 (
            .O(N__6222),
            .I(\U712_CHIP_RAM.N_331 ));
    InMux I__1104 (
            .O(N__6219),
            .I(N__6214));
    InMux I__1103 (
            .O(N__6218),
            .I(N__6211));
    InMux I__1102 (
            .O(N__6217),
            .I(N__6208));
    LocalMux I__1101 (
            .O(N__6214),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__1100 (
            .O(N__6211),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__1099 (
            .O(N__6208),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__1098 (
            .O(N__6201),
            .I(N__6196));
    InMux I__1097 (
            .O(N__6200),
            .I(N__6193));
    InMux I__1096 (
            .O(N__6199),
            .I(N__6190));
    LocalMux I__1095 (
            .O(N__6196),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__1094 (
            .O(N__6193),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__1093 (
            .O(N__6190),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    CascadeMux I__1092 (
            .O(N__6183),
            .I(\U712_CHIP_RAM.N_331_cascade_ ));
    InMux I__1091 (
            .O(N__6180),
            .I(N__6175));
    InMux I__1090 (
            .O(N__6179),
            .I(N__6172));
    InMux I__1089 (
            .O(N__6178),
            .I(N__6169));
    LocalMux I__1088 (
            .O(N__6175),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__1087 (
            .O(N__6172),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__1086 (
            .O(N__6169),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__1085 (
            .O(N__6162),
            .I(N__6158));
    InMux I__1084 (
            .O(N__6161),
            .I(N__6153));
    InMux I__1083 (
            .O(N__6158),
            .I(N__6150));
    InMux I__1082 (
            .O(N__6157),
            .I(N__6147));
    InMux I__1081 (
            .O(N__6156),
            .I(N__6143));
    LocalMux I__1080 (
            .O(N__6153),
            .I(N__6138));
    LocalMux I__1079 (
            .O(N__6150),
            .I(N__6138));
    LocalMux I__1078 (
            .O(N__6147),
            .I(N__6135));
    InMux I__1077 (
            .O(N__6146),
            .I(N__6130));
    LocalMux I__1076 (
            .O(N__6143),
            .I(N__6125));
    Span4Mux_v I__1075 (
            .O(N__6138),
            .I(N__6120));
    Span4Mux_v I__1074 (
            .O(N__6135),
            .I(N__6120));
    InMux I__1073 (
            .O(N__6134),
            .I(N__6117));
    InMux I__1072 (
            .O(N__6133),
            .I(N__6114));
    LocalMux I__1071 (
            .O(N__6130),
            .I(N__6111));
    InMux I__1070 (
            .O(N__6129),
            .I(N__6106));
    InMux I__1069 (
            .O(N__6128),
            .I(N__6106));
    Odrv4 I__1068 (
            .O(N__6125),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__1067 (
            .O(N__6120),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__1066 (
            .O(N__6117),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__1065 (
            .O(N__6114),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__1064 (
            .O(N__6111),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__1063 (
            .O(N__6106),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    CascadeMux I__1062 (
            .O(N__6093),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ));
    InMux I__1061 (
            .O(N__6090),
            .I(N__6087));
    LocalMux I__1060 (
            .O(N__6087),
            .I(N__6082));
    InMux I__1059 (
            .O(N__6086),
            .I(N__6075));
    InMux I__1058 (
            .O(N__6085),
            .I(N__6075));
    Span4Mux_h I__1057 (
            .O(N__6082),
            .I(N__6072));
    InMux I__1056 (
            .O(N__6081),
            .I(N__6067));
    InMux I__1055 (
            .O(N__6080),
            .I(N__6067));
    LocalMux I__1054 (
            .O(N__6075),
            .I(\U712_CHIP_RAM.N_337 ));
    Odrv4 I__1053 (
            .O(N__6072),
            .I(\U712_CHIP_RAM.N_337 ));
    LocalMux I__1052 (
            .O(N__6067),
            .I(\U712_CHIP_RAM.N_337 ));
    InMux I__1051 (
            .O(N__6060),
            .I(N__6055));
    InMux I__1050 (
            .O(N__6059),
            .I(N__6052));
    InMux I__1049 (
            .O(N__6058),
            .I(N__6045));
    LocalMux I__1048 (
            .O(N__6055),
            .I(N__6040));
    LocalMux I__1047 (
            .O(N__6052),
            .I(N__6040));
    InMux I__1046 (
            .O(N__6051),
            .I(N__6037));
    InMux I__1045 (
            .O(N__6050),
            .I(N__6032));
    InMux I__1044 (
            .O(N__6049),
            .I(N__6029));
    InMux I__1043 (
            .O(N__6048),
            .I(N__6025));
    LocalMux I__1042 (
            .O(N__6045),
            .I(N__6022));
    Span4Mux_v I__1041 (
            .O(N__6040),
            .I(N__6017));
    LocalMux I__1040 (
            .O(N__6037),
            .I(N__6017));
    InMux I__1039 (
            .O(N__6036),
            .I(N__6014));
    InMux I__1038 (
            .O(N__6035),
            .I(N__6011));
    LocalMux I__1037 (
            .O(N__6032),
            .I(N__6006));
    LocalMux I__1036 (
            .O(N__6029),
            .I(N__6006));
    InMux I__1035 (
            .O(N__6028),
            .I(N__6003));
    LocalMux I__1034 (
            .O(N__6025),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv12 I__1033 (
            .O(N__6022),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1032 (
            .O(N__6017),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1031 (
            .O(N__6014),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1030 (
            .O(N__6011),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1029 (
            .O(N__6006),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1028 (
            .O(N__6003),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    CascadeMux I__1027 (
            .O(N__5988),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_ ));
    InMux I__1026 (
            .O(N__5985),
            .I(N__5982));
    LocalMux I__1025 (
            .O(N__5982),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    InMux I__1024 (
            .O(N__5979),
            .I(bfn_11_12_0_));
    InMux I__1023 (
            .O(N__5976),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__1022 (
            .O(N__5973),
            .I(N__5970));
    LocalMux I__1021 (
            .O(N__5970),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__1020 (
            .O(N__5967),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__1019 (
            .O(N__5964),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    CascadeMux I__1018 (
            .O(N__5961),
            .I(N__5956));
    InMux I__1017 (
            .O(N__5960),
            .I(N__5953));
    InMux I__1016 (
            .O(N__5959),
            .I(N__5950));
    InMux I__1015 (
            .O(N__5956),
            .I(N__5947));
    LocalMux I__1014 (
            .O(N__5953),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1013 (
            .O(N__5950),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1012 (
            .O(N__5947),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__1011 (
            .O(N__5940),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__1010 (
            .O(N__5937),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__1009 (
            .O(N__5934),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__1008 (
            .O(N__5931),
            .I(N__5915));
    InMux I__1007 (
            .O(N__5930),
            .I(N__5915));
    InMux I__1006 (
            .O(N__5929),
            .I(N__5915));
    InMux I__1005 (
            .O(N__5928),
            .I(N__5915));
    InMux I__1004 (
            .O(N__5927),
            .I(N__5910));
    InMux I__1003 (
            .O(N__5926),
            .I(N__5910));
    InMux I__1002 (
            .O(N__5925),
            .I(N__5905));
    InMux I__1001 (
            .O(N__5924),
            .I(N__5905));
    LocalMux I__1000 (
            .O(N__5915),
            .I(\U712_CHIP_RAM.N_181 ));
    LocalMux I__999 (
            .O(N__5910),
            .I(\U712_CHIP_RAM.N_181 ));
    LocalMux I__998 (
            .O(N__5905),
            .I(\U712_CHIP_RAM.N_181 ));
    InMux I__997 (
            .O(N__5898),
            .I(N__5895));
    LocalMux I__996 (
            .O(N__5895),
            .I(N__5892));
    Sp12to4 I__995 (
            .O(N__5892),
            .I(N__5889));
    Span12Mux_v I__994 (
            .O(N__5889),
            .I(N__5886));
    Span12Mux_h I__993 (
            .O(N__5886),
            .I(N__5883));
    Odrv12 I__992 (
            .O(N__5883),
            .I(A_c_5));
    InMux I__991 (
            .O(N__5880),
            .I(N__5877));
    LocalMux I__990 (
            .O(N__5877),
            .I(N__5874));
    Span4Mux_v I__989 (
            .O(N__5874),
            .I(N__5871));
    Sp12to4 I__988 (
            .O(N__5871),
            .I(N__5868));
    Span12Mux_h I__987 (
            .O(N__5868),
            .I(N__5865));
    Odrv12 I__986 (
            .O(N__5865),
            .I(A_c_12));
    InMux I__985 (
            .O(N__5862),
            .I(N__5859));
    LocalMux I__984 (
            .O(N__5859),
            .I(N__5856));
    Span4Mux_h I__983 (
            .O(N__5856),
            .I(N__5853));
    Span4Mux_h I__982 (
            .O(N__5853),
            .I(N__5850));
    Sp12to4 I__981 (
            .O(N__5850),
            .I(N__5847));
    Span12Mux_v I__980 (
            .O(N__5847),
            .I(N__5844));
    Odrv12 I__979 (
            .O(N__5844),
            .I(A_c_16));
    InMux I__978 (
            .O(N__5841),
            .I(N__5838));
    LocalMux I__977 (
            .O(N__5838),
            .I(N__5835));
    Span4Mux_v I__976 (
            .O(N__5835),
            .I(N__5832));
    Sp12to4 I__975 (
            .O(N__5832),
            .I(N__5829));
    Span12Mux_h I__974 (
            .O(N__5829),
            .I(N__5826));
    Span12Mux_v I__973 (
            .O(N__5826),
            .I(N__5823));
    Odrv12 I__972 (
            .O(N__5823),
            .I(A_c_18));
    CascadeMux I__971 (
            .O(N__5820),
            .I(N__5817));
    InMux I__970 (
            .O(N__5817),
            .I(N__5811));
    InMux I__969 (
            .O(N__5816),
            .I(N__5808));
    InMux I__968 (
            .O(N__5815),
            .I(N__5805));
    InMux I__967 (
            .O(N__5814),
            .I(N__5802));
    LocalMux I__966 (
            .O(N__5811),
            .I(N__5797));
    LocalMux I__965 (
            .O(N__5808),
            .I(N__5797));
    LocalMux I__964 (
            .O(N__5805),
            .I(N__5794));
    LocalMux I__963 (
            .O(N__5802),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    Odrv4 I__962 (
            .O(N__5797),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    Odrv12 I__961 (
            .O(N__5794),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__960 (
            .O(N__5787),
            .I(N__5784));
    InMux I__959 (
            .O(N__5784),
            .I(N__5781));
    LocalMux I__958 (
            .O(N__5781),
            .I(N__5778));
    Span4Mux_v I__957 (
            .O(N__5778),
            .I(N__5774));
    InMux I__956 (
            .O(N__5777),
            .I(N__5771));
    Span4Mux_h I__955 (
            .O(N__5774),
            .I(N__5768));
    LocalMux I__954 (
            .O(N__5771),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    Odrv4 I__953 (
            .O(N__5768),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__952 (
            .O(N__5763),
            .I(\U712_CYCLE_TERM.N_211_i_0_en_cascade_ ));
    CEMux I__951 (
            .O(N__5760),
            .I(N__5757));
    LocalMux I__950 (
            .O(N__5757),
            .I(N__5754));
    Odrv12 I__949 (
            .O(N__5754),
            .I(\U712_CYCLE_TERM.N_211_i_0_en_0 ));
    InMux I__948 (
            .O(N__5751),
            .I(N__5748));
    LocalMux I__947 (
            .O(N__5748),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0 ));
    CEMux I__946 (
            .O(N__5745),
            .I(N__5742));
    LocalMux I__945 (
            .O(N__5742),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0 ));
    CascadeMux I__944 (
            .O(N__5739),
            .I(\U712_CHIP_RAM.N_339_cascade_ ));
    InMux I__943 (
            .O(N__5736),
            .I(N__5732));
    InMux I__942 (
            .O(N__5735),
            .I(N__5727));
    LocalMux I__941 (
            .O(N__5732),
            .I(N__5724));
    InMux I__940 (
            .O(N__5731),
            .I(N__5720));
    InMux I__939 (
            .O(N__5730),
            .I(N__5717));
    LocalMux I__938 (
            .O(N__5727),
            .I(N__5712));
    Span4Mux_h I__937 (
            .O(N__5724),
            .I(N__5712));
    InMux I__936 (
            .O(N__5723),
            .I(N__5709));
    LocalMux I__935 (
            .O(N__5720),
            .I(\U712_CHIP_RAM.N_335 ));
    LocalMux I__934 (
            .O(N__5717),
            .I(\U712_CHIP_RAM.N_335 ));
    Odrv4 I__933 (
            .O(N__5712),
            .I(\U712_CHIP_RAM.N_335 ));
    LocalMux I__932 (
            .O(N__5709),
            .I(\U712_CHIP_RAM.N_335 ));
    CascadeMux I__931 (
            .O(N__5700),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_1_cascade_ ));
    InMux I__930 (
            .O(N__5697),
            .I(N__5693));
    InMux I__929 (
            .O(N__5696),
            .I(N__5690));
    LocalMux I__928 (
            .O(N__5693),
            .I(\U712_CHIP_RAM.N_296 ));
    LocalMux I__927 (
            .O(N__5690),
            .I(\U712_CHIP_RAM.N_296 ));
    CascadeMux I__926 (
            .O(N__5685),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_i_a5_0_1_cascade_ ));
    CascadeMux I__925 (
            .O(N__5682),
            .I(\U712_CHIP_RAM.N_257_cascade_ ));
    InMux I__924 (
            .O(N__5679),
            .I(N__5676));
    LocalMux I__923 (
            .O(N__5676),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_i_0 ));
    CascadeMux I__922 (
            .O(N__5673),
            .I(\U712_CHIP_RAM.N_338_cascade_ ));
    CascadeMux I__921 (
            .O(N__5670),
            .I(N__5658));
    InMux I__920 (
            .O(N__5669),
            .I(N__5655));
    InMux I__919 (
            .O(N__5668),
            .I(N__5648));
    InMux I__918 (
            .O(N__5667),
            .I(N__5648));
    InMux I__917 (
            .O(N__5666),
            .I(N__5648));
    InMux I__916 (
            .O(N__5665),
            .I(N__5642));
    InMux I__915 (
            .O(N__5664),
            .I(N__5637));
    InMux I__914 (
            .O(N__5663),
            .I(N__5637));
    InMux I__913 (
            .O(N__5662),
            .I(N__5632));
    InMux I__912 (
            .O(N__5661),
            .I(N__5632));
    InMux I__911 (
            .O(N__5658),
            .I(N__5629));
    LocalMux I__910 (
            .O(N__5655),
            .I(N__5624));
    LocalMux I__909 (
            .O(N__5648),
            .I(N__5624));
    InMux I__908 (
            .O(N__5647),
            .I(N__5617));
    InMux I__907 (
            .O(N__5646),
            .I(N__5617));
    InMux I__906 (
            .O(N__5645),
            .I(N__5617));
    LocalMux I__905 (
            .O(N__5642),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__904 (
            .O(N__5637),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__903 (
            .O(N__5632),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__902 (
            .O(N__5629),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__901 (
            .O(N__5624),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__900 (
            .O(N__5617),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__899 (
            .O(N__5604),
            .I(N__5601));
    LocalMux I__898 (
            .O(N__5601),
            .I(\U712_CHIP_RAM.N_284_2 ));
    InMux I__897 (
            .O(N__5598),
            .I(N__5594));
    InMux I__896 (
            .O(N__5597),
            .I(N__5591));
    LocalMux I__895 (
            .O(N__5594),
            .I(N__5588));
    LocalMux I__894 (
            .O(N__5591),
            .I(N__5585));
    Odrv4 I__893 (
            .O(N__5588),
            .I(\U712_CHIP_RAM.N_253 ));
    Odrv4 I__892 (
            .O(N__5585),
            .I(\U712_CHIP_RAM.N_253 ));
    InMux I__891 (
            .O(N__5580),
            .I(N__5577));
    LocalMux I__890 (
            .O(N__5577),
            .I(N__5571));
    InMux I__889 (
            .O(N__5576),
            .I(N__5566));
    InMux I__888 (
            .O(N__5575),
            .I(N__5566));
    InMux I__887 (
            .O(N__5574),
            .I(N__5563));
    Span4Mux_v I__886 (
            .O(N__5571),
            .I(N__5556));
    LocalMux I__885 (
            .O(N__5566),
            .I(N__5556));
    LocalMux I__884 (
            .O(N__5563),
            .I(N__5556));
    Odrv4 I__883 (
            .O(N__5556),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    CascadeMux I__882 (
            .O(N__5553),
            .I(\U712_CHIP_RAM.N_284_2_cascade_ ));
    InMux I__881 (
            .O(N__5550),
            .I(N__5547));
    LocalMux I__880 (
            .O(N__5547),
            .I(\U712_CHIP_RAM.N_254 ));
    InMux I__879 (
            .O(N__5544),
            .I(N__5541));
    LocalMux I__878 (
            .O(N__5541),
            .I(\U712_CHIP_RAM.N_322 ));
    InMux I__877 (
            .O(N__5538),
            .I(N__5535));
    LocalMux I__876 (
            .O(N__5535),
            .I(N__5532));
    Odrv4 I__875 (
            .O(N__5532),
            .I(\U712_CHIP_RAM.N_206 ));
    InMux I__874 (
            .O(N__5529),
            .I(N__5525));
    InMux I__873 (
            .O(N__5528),
            .I(N__5520));
    LocalMux I__872 (
            .O(N__5525),
            .I(N__5517));
    InMux I__871 (
            .O(N__5524),
            .I(N__5512));
    InMux I__870 (
            .O(N__5523),
            .I(N__5512));
    LocalMux I__869 (
            .O(N__5520),
            .I(\U712_CHIP_RAM.N_338 ));
    Odrv4 I__868 (
            .O(N__5517),
            .I(\U712_CHIP_RAM.N_338 ));
    LocalMux I__867 (
            .O(N__5512),
            .I(\U712_CHIP_RAM.N_338 ));
    InMux I__866 (
            .O(N__5505),
            .I(N__5502));
    LocalMux I__865 (
            .O(N__5502),
            .I(\U712_CHIP_RAM.N_256 ));
    InMux I__864 (
            .O(N__5499),
            .I(N__5496));
    LocalMux I__863 (
            .O(N__5496),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ));
    CascadeMux I__862 (
            .O(N__5493),
            .I(N__5490));
    InMux I__861 (
            .O(N__5490),
            .I(N__5487));
    LocalMux I__860 (
            .O(N__5487),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    InMux I__859 (
            .O(N__5484),
            .I(N__5481));
    LocalMux I__858 (
            .O(N__5481),
            .I(\U712_CHIP_RAM.N_284 ));
    CascadeMux I__857 (
            .O(N__5478),
            .I(\U712_CHIP_RAM.N_284_cascade_ ));
    InMux I__856 (
            .O(N__5475),
            .I(N__5467));
    InMux I__855 (
            .O(N__5474),
            .I(N__5467));
    InMux I__854 (
            .O(N__5473),
            .I(N__5462));
    InMux I__853 (
            .O(N__5472),
            .I(N__5462));
    LocalMux I__852 (
            .O(N__5467),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__851 (
            .O(N__5462),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__850 (
            .O(N__5457),
            .I(N__5453));
    CascadeMux I__849 (
            .O(N__5456),
            .I(N__5450));
    InMux I__848 (
            .O(N__5453),
            .I(N__5445));
    InMux I__847 (
            .O(N__5450),
            .I(N__5445));
    LocalMux I__846 (
            .O(N__5445),
            .I(N__5440));
    InMux I__845 (
            .O(N__5444),
            .I(N__5437));
    InMux I__844 (
            .O(N__5443),
            .I(N__5434));
    Span4Mux_v I__843 (
            .O(N__5440),
            .I(N__5429));
    LocalMux I__842 (
            .O(N__5437),
            .I(N__5429));
    LocalMux I__841 (
            .O(N__5434),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__840 (
            .O(N__5429),
            .I(DBR_SYNCZ0Z_1));
    InMux I__839 (
            .O(N__5424),
            .I(N__5421));
    LocalMux I__838 (
            .O(N__5421),
            .I(\U712_CHIP_RAM.N_218 ));
    CascadeMux I__837 (
            .O(N__5418),
            .I(\U712_CHIP_RAM.N_218_cascade_ ));
    CascadeMux I__836 (
            .O(N__5415),
            .I(N__5412));
    InMux I__835 (
            .O(N__5412),
            .I(N__5409));
    LocalMux I__834 (
            .O(N__5409),
            .I(N__5405));
    InMux I__833 (
            .O(N__5408),
            .I(N__5402));
    Odrv4 I__832 (
            .O(N__5405),
            .I(\U712_CHIP_RAM.N_259 ));
    LocalMux I__831 (
            .O(N__5402),
            .I(\U712_CHIP_RAM.N_259 ));
    CascadeMux I__830 (
            .O(N__5397),
            .I(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a2_0_a5_0_cascade_ ));
    CascadeMux I__829 (
            .O(N__5394),
            .I(\U712_CHIP_RAM.N_206_cascade_ ));
    InMux I__828 (
            .O(N__5391),
            .I(N__5388));
    LocalMux I__827 (
            .O(N__5388),
            .I(\U712_CHIP_RAM.N_329 ));
    InMux I__826 (
            .O(N__5385),
            .I(N__5382));
    LocalMux I__825 (
            .O(N__5382),
            .I(N__5377));
    InMux I__824 (
            .O(N__5381),
            .I(N__5374));
    InMux I__823 (
            .O(N__5380),
            .I(N__5371));
    Odrv4 I__822 (
            .O(N__5377),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    LocalMux I__821 (
            .O(N__5374),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    LocalMux I__820 (
            .O(N__5371),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    CascadeMux I__819 (
            .O(N__5364),
            .I(\U712_CHIP_RAM.N_323_cascade_ ));
    InMux I__818 (
            .O(N__5361),
            .I(N__5358));
    LocalMux I__817 (
            .O(N__5358),
            .I(\U712_CHIP_RAM.N_374 ));
    InMux I__816 (
            .O(N__5355),
            .I(N__5350));
    InMux I__815 (
            .O(N__5354),
            .I(N__5345));
    InMux I__814 (
            .O(N__5353),
            .I(N__5345));
    LocalMux I__813 (
            .O(N__5350),
            .I(\U712_CHIP_RAM.N_378 ));
    LocalMux I__812 (
            .O(N__5345),
            .I(\U712_CHIP_RAM.N_378 ));
    InMux I__811 (
            .O(N__5340),
            .I(N__5334));
    InMux I__810 (
            .O(N__5339),
            .I(N__5334));
    LocalMux I__809 (
            .O(N__5334),
            .I(\U712_CHIP_RAM.N_184 ));
    CascadeMux I__808 (
            .O(N__5331),
            .I(\U712_CHIP_RAM.N_335_cascade_ ));
    CascadeMux I__807 (
            .O(N__5328),
            .I(N__5324));
    CascadeMux I__806 (
            .O(N__5327),
            .I(N__5321));
    InMux I__805 (
            .O(N__5324),
            .I(N__5318));
    InMux I__804 (
            .O(N__5321),
            .I(N__5315));
    LocalMux I__803 (
            .O(N__5318),
            .I(\U712_CHIP_RAM.N_280 ));
    LocalMux I__802 (
            .O(N__5315),
            .I(\U712_CHIP_RAM.N_280 ));
    SRMux I__801 (
            .O(N__5310),
            .I(N__5307));
    LocalMux I__800 (
            .O(N__5307),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__799 (
            .O(N__5304),
            .I(N__5300));
    InMux I__798 (
            .O(N__5303),
            .I(N__5297));
    LocalMux I__797 (
            .O(N__5300),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    LocalMux I__796 (
            .O(N__5297),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__795 (
            .O(N__5292),
            .I(N__5288));
    InMux I__794 (
            .O(N__5291),
            .I(N__5285));
    LocalMux I__793 (
            .O(N__5288),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    LocalMux I__792 (
            .O(N__5285),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    CascadeMux I__791 (
            .O(N__5280),
            .I(N__5276));
    InMux I__790 (
            .O(N__5279),
            .I(N__5273));
    InMux I__789 (
            .O(N__5276),
            .I(N__5270));
    LocalMux I__788 (
            .O(N__5273),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__787 (
            .O(N__5270),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__786 (
            .O(N__5265),
            .I(N__5261));
    InMux I__785 (
            .O(N__5264),
            .I(N__5258));
    LocalMux I__784 (
            .O(N__5261),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    LocalMux I__783 (
            .O(N__5258),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    InMux I__782 (
            .O(N__5253),
            .I(N__5249));
    InMux I__781 (
            .O(N__5252),
            .I(N__5246));
    LocalMux I__780 (
            .O(N__5249),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__779 (
            .O(N__5246),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__778 (
            .O(N__5241),
            .I(N__5237));
    InMux I__777 (
            .O(N__5240),
            .I(N__5234));
    LocalMux I__776 (
            .O(N__5237),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__775 (
            .O(N__5234),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__774 (
            .O(N__5229),
            .I(N__5225));
    InMux I__773 (
            .O(N__5228),
            .I(N__5222));
    LocalMux I__772 (
            .O(N__5225),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__771 (
            .O(N__5222),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__770 (
            .O(N__5217),
            .I(N__5213));
    InMux I__769 (
            .O(N__5216),
            .I(N__5210));
    LocalMux I__768 (
            .O(N__5213),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__767 (
            .O(N__5210),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    CascadeMux I__766 (
            .O(N__5205),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_ ));
    InMux I__765 (
            .O(N__5202),
            .I(N__5199));
    LocalMux I__764 (
            .O(N__5199),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    InMux I__763 (
            .O(N__5196),
            .I(N__5193));
    LocalMux I__762 (
            .O(N__5193),
            .I(\U712_CHIP_RAM.N_340 ));
    CascadeMux I__761 (
            .O(N__5190),
            .I(\U712_CHIP_RAM.N_340_cascade_ ));
    CascadeMux I__760 (
            .O(N__5187),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_ ));
    InMux I__759 (
            .O(N__5184),
            .I(N__5181));
    LocalMux I__758 (
            .O(N__5181),
            .I(\U712_CHIP_RAM.N_97 ));
    IoInMux I__757 (
            .O(N__5178),
            .I(N__5175));
    LocalMux I__756 (
            .O(N__5175),
            .I(N__5172));
    Span12Mux_s3_v I__755 (
            .O(N__5172),
            .I(N__5169));
    Span12Mux_v I__754 (
            .O(N__5169),
            .I(N__5165));
    InMux I__753 (
            .O(N__5168),
            .I(N__5162));
    Odrv12 I__752 (
            .O(N__5165),
            .I(LATCH_CLK_c));
    LocalMux I__751 (
            .O(N__5162),
            .I(LATCH_CLK_c));
    InMux I__750 (
            .O(N__5157),
            .I(N__5152));
    InMux I__749 (
            .O(N__5156),
            .I(N__5148));
    InMux I__748 (
            .O(N__5155),
            .I(N__5145));
    LocalMux I__747 (
            .O(N__5152),
            .I(N__5142));
    InMux I__746 (
            .O(N__5151),
            .I(N__5139));
    LocalMux I__745 (
            .O(N__5148),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__744 (
            .O(N__5145),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    Odrv4 I__743 (
            .O(N__5142),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__742 (
            .O(N__5139),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__741 (
            .O(N__5130),
            .I(N__5127));
    LocalMux I__740 (
            .O(N__5127),
            .I(\U712_CYCLE_TERM.N_312 ));
    InMux I__739 (
            .O(N__5124),
            .I(N__5121));
    LocalMux I__738 (
            .O(N__5121),
            .I(N__5118));
    Span12Mux_h I__737 (
            .O(N__5118),
            .I(N__5115));
    Span12Mux_v I__736 (
            .O(N__5115),
            .I(N__5112));
    Odrv12 I__735 (
            .O(N__5112),
            .I(A_c_3));
    InMux I__734 (
            .O(N__5109),
            .I(N__5106));
    LocalMux I__733 (
            .O(N__5106),
            .I(N__5103));
    Span12Mux_v I__732 (
            .O(N__5103),
            .I(N__5100));
    Span12Mux_h I__731 (
            .O(N__5100),
            .I(N__5097));
    Odrv12 I__730 (
            .O(N__5097),
            .I(A_c_10));
    InMux I__729 (
            .O(N__5094),
            .I(bfn_10_9_0_));
    InMux I__728 (
            .O(N__5091),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__727 (
            .O(N__5088),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__726 (
            .O(N__5085),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__725 (
            .O(N__5082),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__724 (
            .O(N__5079),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__723 (
            .O(N__5076),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__722 (
            .O(N__5073),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__721 (
            .O(N__5070),
            .I(N__5049));
    ClkMux I__720 (
            .O(N__5069),
            .I(N__5049));
    ClkMux I__719 (
            .O(N__5068),
            .I(N__5049));
    ClkMux I__718 (
            .O(N__5067),
            .I(N__5049));
    ClkMux I__717 (
            .O(N__5066),
            .I(N__5049));
    ClkMux I__716 (
            .O(N__5065),
            .I(N__5049));
    ClkMux I__715 (
            .O(N__5064),
            .I(N__5049));
    GlobalMux I__714 (
            .O(N__5049),
            .I(N__5046));
    gio2CtrlBuf I__713 (
            .O(N__5046),
            .I(C1_c_g));
    InMux I__712 (
            .O(N__5043),
            .I(N__5040));
    LocalMux I__711 (
            .O(N__5040),
            .I(\U712_CHIP_RAM.N_258 ));
    CascadeMux I__710 (
            .O(N__5037),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_ ));
    IoInMux I__709 (
            .O(N__5034),
            .I(N__5031));
    LocalMux I__708 (
            .O(N__5031),
            .I(N__5028));
    Span4Mux_s0_h I__707 (
            .O(N__5028),
            .I(N__5025));
    Span4Mux_h I__706 (
            .O(N__5025),
            .I(N__5022));
    Span4Mux_h I__705 (
            .O(N__5022),
            .I(N__5019));
    Sp12to4 I__704 (
            .O(N__5019),
            .I(N__5016));
    Span12Mux_v I__703 (
            .O(N__5016),
            .I(N__5013));
    Odrv12 I__702 (
            .O(N__5013),
            .I(N_235));
    InMux I__701 (
            .O(N__5010),
            .I(N__5005));
    InMux I__700 (
            .O(N__5009),
            .I(N__4999));
    InMux I__699 (
            .O(N__5008),
            .I(N__4999));
    LocalMux I__698 (
            .O(N__5005),
            .I(N__4996));
    InMux I__697 (
            .O(N__5004),
            .I(N__4993));
    LocalMux I__696 (
            .O(N__4999),
            .I(N__4990));
    Span4Mux_v I__695 (
            .O(N__4996),
            .I(N__4985));
    LocalMux I__694 (
            .O(N__4993),
            .I(N__4985));
    Span4Mux_v I__693 (
            .O(N__4990),
            .I(N__4982));
    Span4Mux_v I__692 (
            .O(N__4985),
            .I(N__4979));
    Sp12to4 I__691 (
            .O(N__4982),
            .I(N__4974));
    Sp12to4 I__690 (
            .O(N__4979),
            .I(N__4974));
    Span12Mux_h I__689 (
            .O(N__4974),
            .I(N__4971));
    Odrv12 I__688 (
            .O(N__4971),
            .I(RnW_c));
    InMux I__687 (
            .O(N__4968),
            .I(N__4965));
    LocalMux I__686 (
            .O(N__4965),
            .I(N__4961));
    InMux I__685 (
            .O(N__4964),
            .I(N__4958));
    Span4Mux_v I__684 (
            .O(N__4961),
            .I(N__4953));
    LocalMux I__683 (
            .O(N__4958),
            .I(N__4953));
    Span4Mux_v I__682 (
            .O(N__4953),
            .I(N__4950));
    Sp12to4 I__681 (
            .O(N__4950),
            .I(N__4947));
    Span12Mux_h I__680 (
            .O(N__4947),
            .I(N__4944));
    Odrv12 I__679 (
            .O(N__4944),
            .I(AWEn_c));
    InMux I__678 (
            .O(N__4941),
            .I(N__4938));
    LocalMux I__677 (
            .O(N__4938),
            .I(\U712_CHIP_RAM.N_222 ));
    InMux I__676 (
            .O(N__4935),
            .I(N__4932));
    LocalMux I__675 (
            .O(N__4932),
            .I(N__4929));
    Span4Mux_v I__674 (
            .O(N__4929),
            .I(N__4926));
    Odrv4 I__673 (
            .O(N__4926),
            .I(\U712_BYTE_ENABLE.N_217 ));
    IoInMux I__672 (
            .O(N__4923),
            .I(N__4920));
    LocalMux I__671 (
            .O(N__4920),
            .I(N__4917));
    Span4Mux_s3_v I__670 (
            .O(N__4917),
            .I(N__4914));
    Span4Mux_h I__669 (
            .O(N__4914),
            .I(N__4911));
    Span4Mux_v I__668 (
            .O(N__4911),
            .I(N__4908));
    Odrv4 I__667 (
            .O(N__4908),
            .I(DMA_LATCH_EN_c));
    InMux I__666 (
            .O(N__4905),
            .I(N__4902));
    LocalMux I__665 (
            .O(N__4902),
            .I(N__4899));
    Span4Mux_v I__664 (
            .O(N__4899),
            .I(N__4896));
    Sp12to4 I__663 (
            .O(N__4896),
            .I(N__4893));
    Span12Mux_h I__662 (
            .O(N__4893),
            .I(N__4890));
    Odrv12 I__661 (
            .O(N__4890),
            .I(A_c_11));
    InMux I__660 (
            .O(N__4887),
            .I(N__4884));
    LocalMux I__659 (
            .O(N__4884),
            .I(N__4881));
    Span12Mux_v I__658 (
            .O(N__4881),
            .I(N__4878));
    Span12Mux_h I__657 (
            .O(N__4878),
            .I(N__4875));
    Odrv12 I__656 (
            .O(N__4875),
            .I(A_c_4));
    CascadeMux I__655 (
            .O(N__4872),
            .I(\U712_CHIP_RAM.N_187_cascade_ ));
    CascadeMux I__654 (
            .O(N__4869),
            .I(\U712_CHIP_RAM.N_316_cascade_ ));
    InMux I__653 (
            .O(N__4866),
            .I(N__4863));
    LocalMux I__652 (
            .O(N__4863),
            .I(\U712_CHIP_RAM.N_316 ));
    InMux I__651 (
            .O(N__4860),
            .I(N__4857));
    LocalMux I__650 (
            .O(N__4857),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a5_1 ));
    CascadeMux I__649 (
            .O(N__4854),
            .I(\U712_CHIP_RAM.N_283_cascade_ ));
    CascadeMux I__648 (
            .O(N__4851),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ));
    InMux I__647 (
            .O(N__4848),
            .I(N__4843));
    InMux I__646 (
            .O(N__4847),
            .I(N__4838));
    InMux I__645 (
            .O(N__4846),
            .I(N__4838));
    LocalMux I__644 (
            .O(N__4843),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    LocalMux I__643 (
            .O(N__4838),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    InMux I__642 (
            .O(N__4833),
            .I(N__4830));
    LocalMux I__641 (
            .O(N__4830),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0 ));
    CascadeMux I__640 (
            .O(N__4827),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_ ));
    CEMux I__639 (
            .O(N__4824),
            .I(N__4821));
    LocalMux I__638 (
            .O(N__4821),
            .I(N__4818));
    Span4Mux_v I__637 (
            .O(N__4818),
            .I(N__4815));
    Span4Mux_h I__636 (
            .O(N__4815),
            .I(N__4812));
    Odrv4 I__635 (
            .O(N__4812),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0 ));
    InMux I__634 (
            .O(N__4809),
            .I(N__4806));
    LocalMux I__633 (
            .O(N__4806),
            .I(N__4803));
    Span4Mux_h I__632 (
            .O(N__4803),
            .I(N__4800));
    Span4Mux_v I__631 (
            .O(N__4800),
            .I(N__4797));
    Span4Mux_v I__630 (
            .O(N__4797),
            .I(N__4794));
    Span4Mux_v I__629 (
            .O(N__4794),
            .I(N__4791));
    Odrv4 I__628 (
            .O(N__4791),
            .I(RAMSPACEn_c));
    InMux I__627 (
            .O(N__4788),
            .I(N__4785));
    LocalMux I__626 (
            .O(N__4785),
            .I(N__4782));
    Span4Mux_v I__625 (
            .O(N__4782),
            .I(N__4778));
    InMux I__624 (
            .O(N__4781),
            .I(N__4775));
    Span4Mux_v I__623 (
            .O(N__4778),
            .I(N__4772));
    LocalMux I__622 (
            .O(N__4775),
            .I(N__4769));
    Sp12to4 I__621 (
            .O(N__4772),
            .I(N__4766));
    Span12Mux_h I__620 (
            .O(N__4769),
            .I(N__4763));
    Span12Mux_h I__619 (
            .O(N__4766),
            .I(N__4760));
    Span12Mux_v I__618 (
            .O(N__4763),
            .I(N__4757));
    Odrv12 I__617 (
            .O(N__4760),
            .I(TSn_c));
    Odrv12 I__616 (
            .O(N__4757),
            .I(TSn_c));
    CascadeMux I__615 (
            .O(N__4752),
            .I(\U712_CHIP_RAM.N_279_cascade_ ));
    CascadeMux I__614 (
            .O(N__4749),
            .I(\U712_BYTE_ENABLE.N_215_cascade_ ));
    IoInMux I__613 (
            .O(N__4746),
            .I(N__4743));
    LocalMux I__612 (
            .O(N__4743),
            .I(N__4740));
    Span12Mux_s11_v I__611 (
            .O(N__4740),
            .I(N__4737));
    Odrv12 I__610 (
            .O(N__4737),
            .I(N_167_i));
    InMux I__609 (
            .O(N__4734),
            .I(N__4728));
    CascadeMux I__608 (
            .O(N__4733),
            .I(N__4718));
    CascadeMux I__607 (
            .O(N__4732),
            .I(N__4715));
    InMux I__606 (
            .O(N__4731),
            .I(N__4712));
    LocalMux I__605 (
            .O(N__4728),
            .I(N__4709));
    InMux I__604 (
            .O(N__4727),
            .I(N__4706));
    InMux I__603 (
            .O(N__4726),
            .I(N__4697));
    InMux I__602 (
            .O(N__4725),
            .I(N__4697));
    InMux I__601 (
            .O(N__4724),
            .I(N__4697));
    InMux I__600 (
            .O(N__4723),
            .I(N__4697));
    InMux I__599 (
            .O(N__4722),
            .I(N__4688));
    InMux I__598 (
            .O(N__4721),
            .I(N__4688));
    InMux I__597 (
            .O(N__4718),
            .I(N__4688));
    InMux I__596 (
            .O(N__4715),
            .I(N__4688));
    LocalMux I__595 (
            .O(N__4712),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__594 (
            .O(N__4709),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__593 (
            .O(N__4706),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__592 (
            .O(N__4697),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__591 (
            .O(N__4688),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    IoInMux I__590 (
            .O(N__4677),
            .I(N__4674));
    LocalMux I__589 (
            .O(N__4674),
            .I(N__4670));
    IoInMux I__588 (
            .O(N__4673),
            .I(N__4667));
    Span4Mux_s2_v I__587 (
            .O(N__4670),
            .I(N__4664));
    LocalMux I__586 (
            .O(N__4667),
            .I(N__4661));
    Span4Mux_h I__585 (
            .O(N__4664),
            .I(N__4658));
    IoSpan4Mux I__584 (
            .O(N__4661),
            .I(N__4655));
    Span4Mux_v I__583 (
            .O(N__4658),
            .I(N__4652));
    Span4Mux_s3_v I__582 (
            .O(N__4655),
            .I(N__4649));
    Span4Mux_v I__581 (
            .O(N__4652),
            .I(N__4646));
    Span4Mux_h I__580 (
            .O(N__4649),
            .I(N__4643));
    Sp12to4 I__579 (
            .O(N__4646),
            .I(N__4640));
    Span4Mux_v I__578 (
            .O(N__4643),
            .I(N__4637));
    Odrv12 I__577 (
            .O(N__4640),
            .I(ASn_c));
    Odrv4 I__576 (
            .O(N__4637),
            .I(ASn_c));
    CEMux I__575 (
            .O(N__4632),
            .I(N__4629));
    LocalMux I__574 (
            .O(N__4629),
            .I(N__4626));
    Span4Mux_h I__573 (
            .O(N__4626),
            .I(N__4623));
    Odrv4 I__572 (
            .O(N__4623),
            .I(\U712_REG_SM.N_219_0_0 ));
    InMux I__571 (
            .O(N__4620),
            .I(N__4617));
    LocalMux I__570 (
            .O(N__4617),
            .I(N__4614));
    Sp12to4 I__569 (
            .O(N__4614),
            .I(N__4611));
    Span12Mux_v I__568 (
            .O(N__4611),
            .I(N__4608));
    Span12Mux_h I__567 (
            .O(N__4608),
            .I(N__4605));
    Odrv12 I__566 (
            .O(N__4605),
            .I(A_c_6));
    InMux I__565 (
            .O(N__4602),
            .I(N__4599));
    LocalMux I__564 (
            .O(N__4599),
            .I(N__4596));
    Span4Mux_v I__563 (
            .O(N__4596),
            .I(N__4593));
    Sp12to4 I__562 (
            .O(N__4593),
            .I(N__4590));
    Odrv12 I__561 (
            .O(N__4590),
            .I(A_c_13));
    IoInMux I__560 (
            .O(N__4587),
            .I(N__4584));
    LocalMux I__559 (
            .O(N__4584),
            .I(N__4581));
    Span4Mux_s3_v I__558 (
            .O(N__4581),
            .I(N__4578));
    Span4Mux_v I__557 (
            .O(N__4578),
            .I(N__4575));
    Span4Mux_v I__556 (
            .O(N__4575),
            .I(N__4572));
    Span4Mux_v I__555 (
            .O(N__4572),
            .I(N__4568));
    InMux I__554 (
            .O(N__4571),
            .I(N__4565));
    Odrv4 I__553 (
            .O(N__4568),
            .I(DBDIR_c));
    LocalMux I__552 (
            .O(N__4565),
            .I(DBDIR_c));
    InMux I__551 (
            .O(N__4560),
            .I(N__4555));
    InMux I__550 (
            .O(N__4559),
            .I(N__4550));
    InMux I__549 (
            .O(N__4558),
            .I(N__4550));
    LocalMux I__548 (
            .O(N__4555),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__547 (
            .O(N__4550),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    IoInMux I__546 (
            .O(N__4545),
            .I(N__4542));
    LocalMux I__545 (
            .O(N__4542),
            .I(N__4539));
    Span4Mux_s1_h I__544 (
            .O(N__4539),
            .I(N__4536));
    Sp12to4 I__543 (
            .O(N__4536),
            .I(N__4533));
    Span12Mux_v I__542 (
            .O(N__4533),
            .I(N__4529));
    InMux I__541 (
            .O(N__4532),
            .I(N__4526));
    Odrv12 I__540 (
            .O(N__4529),
            .I(TACK_OUTn));
    LocalMux I__539 (
            .O(N__4526),
            .I(TACK_OUTn));
    IoInMux I__538 (
            .O(N__4521),
            .I(N__4518));
    LocalMux I__537 (
            .O(N__4518),
            .I(N__4515));
    IoSpan4Mux I__536 (
            .O(N__4515),
            .I(N__4512));
    Sp12to4 I__535 (
            .O(N__4512),
            .I(N__4509));
    Span12Mux_s7_h I__534 (
            .O(N__4509),
            .I(N__4506));
    Span12Mux_h I__533 (
            .O(N__4506),
            .I(N__4503));
    Odrv12 I__532 (
            .O(N__4503),
            .I(N_165_i));
    InMux I__531 (
            .O(N__4500),
            .I(N__4497));
    LocalMux I__530 (
            .O(N__4497),
            .I(N__4494));
    Span4Mux_v I__529 (
            .O(N__4494),
            .I(N__4490));
    InMux I__528 (
            .O(N__4493),
            .I(N__4487));
    Odrv4 I__527 (
            .O(N__4490),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_a5_0Z0Z_0 ));
    LocalMux I__526 (
            .O(N__4487),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_a5_0Z0Z_0 ));
    CascadeMux I__525 (
            .O(N__4482),
            .I(N__4479));
    InMux I__524 (
            .O(N__4479),
            .I(N__4476));
    LocalMux I__523 (
            .O(N__4476),
            .I(N__4473));
    Span4Mux_h I__522 (
            .O(N__4473),
            .I(N__4470));
    Span4Mux_h I__521 (
            .O(N__4470),
            .I(N__4467));
    Sp12to4 I__520 (
            .O(N__4467),
            .I(N__4464));
    Span12Mux_v I__519 (
            .O(N__4464),
            .I(N__4461));
    Odrv12 I__518 (
            .O(N__4461),
            .I(REGSPACEn_c));
    InMux I__517 (
            .O(N__4458),
            .I(N__4455));
    LocalMux I__516 (
            .O(N__4455),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_i_i_0 ));
    CascadeMux I__515 (
            .O(N__4452),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_i_i_0_cascade_ ));
    InMux I__514 (
            .O(N__4449),
            .I(N__4446));
    LocalMux I__513 (
            .O(N__4446),
            .I(\U712_CHIP_RAM.N_23 ));
    InMux I__512 (
            .O(N__4443),
            .I(N__4439));
    InMux I__511 (
            .O(N__4442),
            .I(N__4436));
    LocalMux I__510 (
            .O(N__4439),
            .I(\U712_REG_SM.N_219 ));
    LocalMux I__509 (
            .O(N__4436),
            .I(\U712_REG_SM.N_219 ));
    InMux I__508 (
            .O(N__4431),
            .I(N__4424));
    InMux I__507 (
            .O(N__4430),
            .I(N__4424));
    InMux I__506 (
            .O(N__4429),
            .I(N__4421));
    LocalMux I__505 (
            .O(N__4424),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__504 (
            .O(N__4421),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__503 (
            .O(N__4416),
            .I(N__4413));
    LocalMux I__502 (
            .O(N__4413),
            .I(\U712_REG_SM.N_261 ));
    InMux I__501 (
            .O(N__4410),
            .I(N__4407));
    LocalMux I__500 (
            .O(N__4407),
            .I(\U712_REG_SM.DS_EN_RNOZ0Z_0 ));
    CascadeMux I__499 (
            .O(N__4404),
            .I(N__4401));
    InMux I__498 (
            .O(N__4401),
            .I(N__4393));
    InMux I__497 (
            .O(N__4400),
            .I(N__4388));
    InMux I__496 (
            .O(N__4399),
            .I(N__4388));
    InMux I__495 (
            .O(N__4398),
            .I(N__4385));
    InMux I__494 (
            .O(N__4397),
            .I(N__4380));
    InMux I__493 (
            .O(N__4396),
            .I(N__4380));
    LocalMux I__492 (
            .O(N__4393),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__491 (
            .O(N__4388),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__490 (
            .O(N__4385),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__489 (
            .O(N__4380),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    InMux I__488 (
            .O(N__4371),
            .I(N__4367));
    InMux I__487 (
            .O(N__4370),
            .I(N__4364));
    LocalMux I__486 (
            .O(N__4367),
            .I(N__4361));
    LocalMux I__485 (
            .O(N__4364),
            .I(N__4358));
    Span4Mux_v I__484 (
            .O(N__4361),
            .I(N__4355));
    Span4Mux_v I__483 (
            .O(N__4358),
            .I(N__4352));
    Sp12to4 I__482 (
            .O(N__4355),
            .I(N__4349));
    Span4Mux_h I__481 (
            .O(N__4352),
            .I(N__4346));
    Span12Mux_h I__480 (
            .O(N__4349),
            .I(N__4341));
    Sp12to4 I__479 (
            .O(N__4346),
            .I(N__4341));
    Odrv12 I__478 (
            .O(N__4341),
            .I(DBRn_c));
    InMux I__477 (
            .O(N__4338),
            .I(N__4335));
    LocalMux I__476 (
            .O(N__4335),
            .I(N__4332));
    Odrv4 I__475 (
            .O(N__4332),
            .I(DBR_SYNCZ0Z_0));
    InMux I__474 (
            .O(N__4329),
            .I(N__4326));
    LocalMux I__473 (
            .O(N__4326),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__472 (
            .O(N__4323),
            .I(N__4319));
    InMux I__471 (
            .O(N__4322),
            .I(N__4310));
    LocalMux I__470 (
            .O(N__4319),
            .I(N__4307));
    InMux I__469 (
            .O(N__4318),
            .I(N__4304));
    InMux I__468 (
            .O(N__4317),
            .I(N__4299));
    InMux I__467 (
            .O(N__4316),
            .I(N__4299));
    InMux I__466 (
            .O(N__4315),
            .I(N__4292));
    InMux I__465 (
            .O(N__4314),
            .I(N__4292));
    InMux I__464 (
            .O(N__4313),
            .I(N__4292));
    LocalMux I__463 (
            .O(N__4310),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__462 (
            .O(N__4307),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__461 (
            .O(N__4304),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__460 (
            .O(N__4299),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__459 (
            .O(N__4292),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__458 (
            .O(N__4281),
            .I(N__4277));
    IoInMux I__457 (
            .O(N__4280),
            .I(N__4274));
    LocalMux I__456 (
            .O(N__4277),
            .I(N__4271));
    LocalMux I__455 (
            .O(N__4274),
            .I(N__4268));
    Span4Mux_v I__454 (
            .O(N__4271),
            .I(N__4265));
    IoSpan4Mux I__453 (
            .O(N__4268),
            .I(N__4262));
    Sp12to4 I__452 (
            .O(N__4265),
            .I(N__4259));
    IoSpan4Mux I__451 (
            .O(N__4262),
            .I(N__4256));
    Span12Mux_h I__450 (
            .O(N__4259),
            .I(N__4253));
    IoSpan4Mux I__449 (
            .O(N__4256),
            .I(N__4250));
    Odrv12 I__448 (
            .O(N__4253),
            .I(C1_c));
    Odrv4 I__447 (
            .O(N__4250),
            .I(C1_c));
    InMux I__446 (
            .O(N__4245),
            .I(N__4242));
    LocalMux I__445 (
            .O(N__4242),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    IoInMux I__444 (
            .O(N__4239),
            .I(N__4236));
    LocalMux I__443 (
            .O(N__4236),
            .I(N__4233));
    Span12Mux_s11_v I__442 (
            .O(N__4233),
            .I(N__4230));
    Odrv12 I__441 (
            .O(N__4230),
            .I(VBENn_c));
    InMux I__440 (
            .O(N__4227),
            .I(N__4221));
    InMux I__439 (
            .O(N__4226),
            .I(N__4221));
    LocalMux I__438 (
            .O(N__4221),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    CascadeMux I__437 (
            .O(N__4218),
            .I(N__4215));
    InMux I__436 (
            .O(N__4215),
            .I(N__4212));
    LocalMux I__435 (
            .O(N__4212),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a5_0_0_0 ));
    InMux I__434 (
            .O(N__4209),
            .I(N__4204));
    InMux I__433 (
            .O(N__4208),
            .I(N__4199));
    InMux I__432 (
            .O(N__4207),
            .I(N__4199));
    LocalMux I__431 (
            .O(N__4204),
            .I(\U712_REG_SM.N_209 ));
    LocalMux I__430 (
            .O(N__4199),
            .I(\U712_REG_SM.N_209 ));
    CascadeMux I__429 (
            .O(N__4194),
            .I(\U712_REG_SM.STATE_COUNTc_1_0_cascade_ ));
    CascadeMux I__428 (
            .O(N__4191),
            .I(\U712_REG_SM.N_272_cascade_ ));
    InMux I__427 (
            .O(N__4188),
            .I(N__4180));
    InMux I__426 (
            .O(N__4187),
            .I(N__4173));
    InMux I__425 (
            .O(N__4186),
            .I(N__4173));
    InMux I__424 (
            .O(N__4185),
            .I(N__4173));
    InMux I__423 (
            .O(N__4184),
            .I(N__4170));
    InMux I__422 (
            .O(N__4183),
            .I(N__4167));
    LocalMux I__421 (
            .O(N__4180),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__420 (
            .O(N__4173),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__419 (
            .O(N__4170),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__418 (
            .O(N__4167),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    CascadeMux I__417 (
            .O(N__4158),
            .I(N__4155));
    InMux I__416 (
            .O(N__4155),
            .I(N__4143));
    InMux I__415 (
            .O(N__4154),
            .I(N__4143));
    InMux I__414 (
            .O(N__4153),
            .I(N__4143));
    InMux I__413 (
            .O(N__4152),
            .I(N__4143));
    LocalMux I__412 (
            .O(N__4143),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    InMux I__411 (
            .O(N__4140),
            .I(N__4137));
    LocalMux I__410 (
            .O(N__4137),
            .I(\U712_REG_SM.STATE_COUNT_srsts_i_0_a5_0_0_0 ));
    InMux I__409 (
            .O(N__4134),
            .I(N__4131));
    LocalMux I__408 (
            .O(N__4131),
            .I(N__4127));
    InMux I__407 (
            .O(N__4130),
            .I(N__4124));
    Odrv4 I__406 (
            .O(N__4127),
            .I(\U712_REG_SM.N_207 ));
    LocalMux I__405 (
            .O(N__4124),
            .I(\U712_REG_SM.N_207 ));
    CascadeMux I__404 (
            .O(N__4119),
            .I(N__4114));
    CascadeMux I__403 (
            .O(N__4118),
            .I(N__4109));
    InMux I__402 (
            .O(N__4117),
            .I(N__4105));
    InMux I__401 (
            .O(N__4114),
            .I(N__4102));
    InMux I__400 (
            .O(N__4113),
            .I(N__4099));
    InMux I__399 (
            .O(N__4112),
            .I(N__4096));
    InMux I__398 (
            .O(N__4109),
            .I(N__4091));
    InMux I__397 (
            .O(N__4108),
            .I(N__4091));
    LocalMux I__396 (
            .O(N__4105),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__395 (
            .O(N__4102),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__394 (
            .O(N__4099),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__393 (
            .O(N__4096),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__392 (
            .O(N__4091),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    InMux I__391 (
            .O(N__4080),
            .I(N__4077));
    LocalMux I__390 (
            .O(N__4077),
            .I(\U712_REG_SM.N_191 ));
    InMux I__389 (
            .O(N__4074),
            .I(N__4071));
    LocalMux I__388 (
            .O(N__4071),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    CascadeMux I__387 (
            .O(N__4068),
            .I(\U712_REG_SM.N_191_cascade_ ));
    IoInMux I__386 (
            .O(N__4065),
            .I(N__4062));
    LocalMux I__385 (
            .O(N__4062),
            .I(N__4059));
    IoSpan4Mux I__384 (
            .O(N__4059),
            .I(N__4056));
    Span4Mux_s3_h I__383 (
            .O(N__4056),
            .I(N__4053));
    Span4Mux_v I__382 (
            .O(N__4053),
            .I(N__4050));
    Span4Mux_h I__381 (
            .O(N__4050),
            .I(N__4047));
    Sp12to4 I__380 (
            .O(N__4047),
            .I(N__4043));
    InMux I__379 (
            .O(N__4046),
            .I(N__4040));
    Span12Mux_h I__378 (
            .O(N__4043),
            .I(N__4035));
    LocalMux I__377 (
            .O(N__4040),
            .I(N__4035));
    Span12Mux_h I__376 (
            .O(N__4035),
            .I(N__4032));
    Odrv12 I__375 (
            .O(N__4032),
            .I(C3_c));
    InMux I__374 (
            .O(N__4029),
            .I(N__4026));
    LocalMux I__373 (
            .O(N__4026),
            .I(\U712_REG_SM.N_85 ));
    InMux I__372 (
            .O(N__4023),
            .I(N__4020));
    LocalMux I__371 (
            .O(N__4020),
            .I(N__4017));
    Odrv4 I__370 (
            .O(N__4017),
            .I(\U712_REG_SM.N_263 ));
    IoInMux I__369 (
            .O(N__4014),
            .I(N__4011));
    LocalMux I__368 (
            .O(N__4011),
            .I(N__4008));
    Span12Mux_s8_h I__367 (
            .O(N__4008),
            .I(N__4005));
    Odrv12 I__366 (
            .O(N__4005),
            .I(N_812_i));
    InMux I__365 (
            .O(N__4002),
            .I(N__3999));
    LocalMux I__364 (
            .O(N__3999),
            .I(N__3996));
    Span4Mux_v I__363 (
            .O(N__3996),
            .I(N__3993));
    Odrv4 I__362 (
            .O(N__3993),
            .I(TACK_EN_i_ess));
    IoInMux I__361 (
            .O(N__3990),
            .I(N__3987));
    LocalMux I__360 (
            .O(N__3987),
            .I(N__3984));
    IoSpan4Mux I__359 (
            .O(N__3984),
            .I(N__3981));
    Span4Mux_s3_h I__358 (
            .O(N__3981),
            .I(N__3978));
    Span4Mux_h I__357 (
            .O(N__3978),
            .I(N__3975));
    Odrv4 I__356 (
            .O(N__3975),
            .I(DBRn_c_i_0));
    CascadeMux I__355 (
            .O(N__3972),
            .I(\U712_REG_SM.N_266_cascade_ ));
    CascadeMux I__354 (
            .O(N__3969),
            .I(\U712_REG_SM.N_269_cascade_ ));
    InMux I__353 (
            .O(N__3966),
            .I(N__3962));
    InMux I__352 (
            .O(N__3965),
            .I(N__3959));
    LocalMux I__351 (
            .O(N__3962),
            .I(\U712_REG_SM.N_233 ));
    LocalMux I__350 (
            .O(N__3959),
            .I(\U712_REG_SM.N_233 ));
    IoInMux I__349 (
            .O(N__3954),
            .I(N__3951));
    LocalMux I__348 (
            .O(N__3951),
            .I(N__3948));
    Span4Mux_s2_v I__347 (
            .O(N__3948),
            .I(N__3945));
    Span4Mux_v I__346 (
            .O(N__3945),
            .I(N__3942));
    Odrv4 I__345 (
            .O(N__3942),
            .I(CLK80_PLL_i_i));
    IoInMux I__344 (
            .O(N__3939),
            .I(N__3936));
    LocalMux I__343 (
            .O(N__3936),
            .I(N__3933));
    IoSpan4Mux I__342 (
            .O(N__3933),
            .I(N__3930));
    Span4Mux_s2_v I__341 (
            .O(N__3930),
            .I(N__3927));
    Sp12to4 I__340 (
            .O(N__3927),
            .I(N__3924));
    Span12Mux_v I__339 (
            .O(N__3924),
            .I(N__3921));
    Odrv12 I__338 (
            .O(N__3921),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__5067));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .I(N__5068));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__5070));
    INV \INVU712_CHIP_RAM.DMA_A20C  (
            .O(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .I(N__5064));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__5066));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__5065));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_9_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7590),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__4280),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__3990),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__4065),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_2_1_1.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_2_1_1.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_2_1_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_2_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9663),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_obuft_RNO_LC_5_15_6.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_5_15_6.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_5_15_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 TACKn_obuft_RNO_LC_5_15_6 (
            .in0(N__4002),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_812_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_6_11_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_6_11_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_6_11_0 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_6_11_0  (
            .in0(N__7741),
            .in1(N__5814),
            .in2(_gnd_net_),
            .in3(N__7448),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9648),
            .ce(N__5760),
            .sr(N__10812));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_6_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_6_12_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_6_12_0  (
            .in0(_gnd_net_),
            .in1(N__10848),
            .in2(_gnd_net_),
            .in3(N__10460),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_6_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_6_12_1 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_6_12_1  (
            .in0(N__5010),
            .in1(N__4113),
            .in2(_gnd_net_),
            .in3(N__3965),
            .lcout(\U712_REG_SM.N_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_6_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_6_13_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_6_13_1  (
            .in0(N__4400),
            .in1(N__4208),
            .in2(_gnd_net_),
            .in3(N__4725),
            .lcout(),
            .ltout(\U712_REG_SM.N_266_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_6_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_6_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_6_13_2 .LUT_INIT=16'b1110101011100010;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_6_13_2  (
            .in0(N__10653),
            .in1(N__7780),
            .in2(N__3972),
            .in3(N__3966),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9654),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_6_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_6_13_3 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_6_13_3  (
            .in0(N__4399),
            .in1(_gnd_net_),
            .in2(N__4118),
            .in3(N__4207),
            .lcout(),
            .ltout(\U712_REG_SM.N_269_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_6_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_6_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_6_13_4 .LUT_INIT=16'b0000101100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_6_13_4  (
            .in0(N__4726),
            .in1(N__4323),
            .in2(N__3969),
            .in3(N__7781),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9654),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_6_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_6_13_5 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_6_13_5  (
            .in0(N__4108),
            .in1(N__4724),
            .in2(_gnd_net_),
            .in3(N__4317),
            .lcout(\U712_REG_SM.N_263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_6_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_6_13_7 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_6_13_7  (
            .in0(N__4184),
            .in1(N__4316),
            .in2(_gnd_net_),
            .in3(N__4723),
            .lcout(\U712_REG_SM.N_233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_6_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_6_14_0 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_6_14_0  (
            .in0(N__4185),
            .in1(N__5004),
            .in2(_gnd_net_),
            .in3(N__4398),
            .lcout(\U712_REG_SM.DS_EN_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_6_14_3.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_6_14_3.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_6_14_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_6_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4370),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_6_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_6_14_6 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_6_14_6  (
            .in0(N__4186),
            .in1(N__4318),
            .in2(_gnd_net_),
            .in3(N__4727),
            .lcout(\U712_REG_SM.N_191 ),
            .ltout(\U712_REG_SM.N_191_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_6_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_6_14_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_6_14_7 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_6_14_7  (
            .in0(N__4117),
            .in1(N__7782),
            .in2(N__4068),
            .in3(N__4187),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9656),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_0_LC_6_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_6_15_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_6_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_6_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4046),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9659),
            .ce(),
            .sr(N__10783));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_7_11_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_7_11_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_7_11_0 .LUT_INIT=16'b0011001000100010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_7_11_0  (
            .in0(N__5777),
            .in1(N__5157),
            .in2(N__4218),
            .in3(N__7449),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9644),
            .ce(),
            .sr(N__10805));
    defparam \U712_REG_SM.REG_TACK_LC_7_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_7_11_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_7_11_4  (
            .in0(N__4134),
            .in1(N__4029),
            .in2(N__7473),
            .in3(N__4023),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9644),
            .ce(),
            .sr(N__10805));
    defparam DBR_SYNC_1_LC_7_12_4.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_7_12_4.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_7_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_7_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4338),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9649),
            .ce(),
            .sr(N__10799));
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_7_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_7_13_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_7_13_0  (
            .in0(N__4153),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4396),
            .lcout(\U712_REG_SM.N_207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_7_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_7_13_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__4314),
            .in2(_gnd_net_),
            .in3(N__5443),
            .lcout(\U712_REG_SM.N_209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_7_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_7_13_2 .LUT_INIT=16'b0000000011101111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_7_13_2  (
            .in0(N__4315),
            .in1(N__4721),
            .in2(N__4158),
            .in3(N__4397),
            .lcout(),
            .ltout(\U712_REG_SM.STATE_COUNTc_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_7_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_7_13_3 .LUT_INIT=16'b0000100000001010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_7_13_3  (
            .in0(N__7779),
            .in1(N__4209),
            .in2(N__4194),
            .in3(N__4731),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9653),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_7_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_7_13_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_7_13_4  (
            .in0(N__4188),
            .in1(N__4431),
            .in2(_gnd_net_),
            .in3(N__4112),
            .lcout(\U712_REG_SM.STATE_COUNT_srsts_i_0_a5_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_13_5 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_13_5  (
            .in0(N__4430),
            .in1(N__4154),
            .in2(N__4733),
            .in3(N__4074),
            .lcout(),
            .ltout(\U712_REG_SM.N_272_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_7_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_7_13_6 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_7_13_6  (
            .in0(N__7778),
            .in1(N__4322),
            .in2(N__4191),
            .in3(N__4722),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9653),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_7_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_7_13_7 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_7_13_7  (
            .in0(N__4183),
            .in1(N__4313),
            .in2(N__4732),
            .in3(N__4152),
            .lcout(\U712_REG_SM.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_7_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_7_14_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_7_14_1 .LUT_INIT=16'b0010001000100011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_7_14_1  (
            .in0(N__4140),
            .in1(N__4130),
            .in2(N__4119),
            .in3(N__4080),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9655),
            .ce(),
            .sr(N__10784));
    defparam \U712_REG_SM.C1_SYNC_1_LC_7_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_7_14_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_7_14_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__4245),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9655),
            .ce(),
            .sr(N__10784));
    defparam \U712_REG_SM.DS_EN_LC_7_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_7_14_4 .LUT_INIT=16'b0011101000110011;
    LogicCell40 \U712_REG_SM.DS_EN_LC_7_14_4  (
            .in0(N__7819),
            .in1(N__4410),
            .in2(N__4404),
            .in3(N__4443),
            .lcout(DS_ENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9655),
            .ce(),
            .sr(N__10784));
    defparam DBR_SYNC_0_LC_7_14_6.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_7_14_6.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_7_14_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 DBR_SYNC_0_LC_7_14_6 (
            .in0(N__4371),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9655),
            .ce(),
            .sr(N__10784));
    defparam \U712_REG_SM.C3_SYNC_1_LC_7_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_7_14_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_7_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4329),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9655),
            .ce(),
            .sr(N__10784));
    defparam \U712_REG_SM.C1_SYNC_0_LC_7_15_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_7_15_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_7_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4281),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9657),
            .ce(),
            .sr(N__10773));
    defparam \U712_BUFFERS.un1_VBENn_0_a5_LC_8_6_4 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a5_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a5_LC_8_6_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a5_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__9369),
            .in2(_gnd_net_),
            .in3(N__10673),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_10_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_10_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_8_10_0  (
            .in0(N__7749),
            .in1(N__6867),
            .in2(_gnd_net_),
            .in3(N__5156),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9637),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_10_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_10_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_8_10_3  (
            .in0(N__4227),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7750),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9637),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_10_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_8_10_5  (
            .in0(N__4559),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7751),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9637),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_10_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_10_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__4558),
            .in2(_gnd_net_),
            .in3(N__4226),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a5_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_8_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_8_11_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_8_11_0 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_8_11_0  (
            .in0(N__4833),
            .in1(N__6984),
            .in2(N__6162),
            .in3(N__8952),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9640),
            .ce(),
            .sr(N__10800));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_12_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_12_0  (
            .in0(N__5665),
            .in1(N__6060),
            .in2(_gnd_net_),
            .in3(N__6161),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9645),
            .ce(N__4824),
            .sr(N__10789));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_13_0 .LUT_INIT=16'b1111000000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_13_0  (
            .in0(N__5043),
            .in1(N__4458),
            .in2(N__9733),
            .in3(N__4847),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9650),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_8_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_8_13_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_8_13_1  (
            .in0(N__4846),
            .in1(N__4449),
            .in2(_gnd_net_),
            .in3(N__8432),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9650),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_13_3 .LUT_INIT=16'b1010101000000010;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_8_13_3  (
            .in0(N__7748),
            .in1(N__4781),
            .in2(N__4482),
            .in3(N__4416),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9650),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_8_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_8_13_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_0_LC_8_13_5  (
            .in0(N__6059),
            .in1(N__6146),
            .in2(_gnd_net_),
            .in3(N__10443),
            .lcout(\U712_CHIP_RAM.N_288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIE24B8_LC_8_14_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIE24B8_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIE24B8_LC_8_14_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIE24B8_LC_8_14_1  (
            .in0(N__5597),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6090),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_i_i_0 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_i_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_8_14_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_8_14_2 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__5529),
            .in2(N__4452),
            .in3(N__5736),
            .lcout(\U712_CHIP_RAM.N_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_RNO_LC_8_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_8_14_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U712_REG_SM.ASn_ess_RNO_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__10845),
            .in2(_gnd_net_),
            .in3(N__4442),
            .lcout(\U712_REG_SM.N_219_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_8_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_8_14_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__4429),
            .in2(_gnd_net_),
            .in3(N__10666),
            .lcout(\U712_REG_SM.N_261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_i_o5_LC_8_15_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_i_o5_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_i_o5_LC_8_15_2 .LUT_INIT=16'b1110110111100101;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_i_o5_LC_8_15_2  (
            .in0(N__8639),
            .in1(N__8816),
            .in2(N__8606),
            .in3(N__8728),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_167_i_LC_8_15_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_167_i_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_167_i_LC_8_15_3 .LUT_INIT=16'b0000110111011101;
    LogicCell40 \U712_BYTE_ENABLE.N_167_i_LC_8_15_3  (
            .in0(N__4500),
            .in1(N__10544),
            .in2(N__4749),
            .in3(N__9392),
            .lcout(N_167_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_LC_8_16_4 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_LC_8_16_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_ess_LC_8_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.ASn_ess_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4734),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9658),
            .ce(N__4632),
            .sr(N__10770));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_6_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_6_1  (
            .in0(N__4620),
            .in1(N__4602),
            .in2(_gnd_net_),
            .in3(N__9104),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_9_9_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_9_9_5  (
            .in0(N__8373),
            .in1(N__9734),
            .in2(N__8457),
            .in3(N__9127),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBDIR_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_10_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_10_1 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_9_10_1  (
            .in0(N__4968),
            .in1(N__4571),
            .in2(_gnd_net_),
            .in3(N__5385),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9634),
            .ce(),
            .sr(N__10801));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_9_10_7 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_9_10_7 .LUT_INIT=16'b1110110011101110;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_9_10_7  (
            .in0(N__4532),
            .in1(N__4560),
            .in2(N__6866),
            .in3(N__5155),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9634),
            .ce(),
            .sr(N__10801));
    defparam \U712_BYTE_ENABLE.N_165_i_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_165_i_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_165_i_LC_9_11_0 .LUT_INIT=16'b0011000111110101;
    LogicCell40 \U712_BYTE_ENABLE.N_165_i_LC_9_11_0  (
            .in0(N__4493),
            .in1(N__4935),
            .in2(N__10628),
            .in3(N__9379),
            .lcout(N_165_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a5_0_0_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a5_0_0_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a5_0_0_LC_9_11_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_a5_0_0_LC_9_11_2  (
            .in0(N__7037),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6985),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_a5_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIALFTC_2_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIALFTC_2_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIALFTC_2_LC_9_11_3 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIALFTC_2_LC_9_11_3  (
            .in0(N__5196),
            .in1(N__6663),
            .in2(N__5327),
            .in3(N__5380),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_11_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4827),
            .in3(N__10846),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_11_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_11_5 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_9_11_5  (
            .in0(N__7646),
            .in1(N__6849),
            .in2(N__5820),
            .in3(N__5130),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9638),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_9_11_7 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__7036),
            .in2(_gnd_net_),
            .in3(N__7160),
            .lcout(\U712_CHIP_RAM.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_1_LC_9_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_1_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_1_LC_9_12_0 .LUT_INIT=16'b0000100010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_1_LC_9_12_0  (
            .in0(N__7241),
            .in1(N__7746),
            .in2(N__6573),
            .in3(N__7148),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_12_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__9383),
            .in2(_gnd_net_),
            .in3(N__5473),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_279_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_12_2 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_12_2  (
            .in0(N__4809),
            .in1(N__4788),
            .in2(N__4752),
            .in3(N__7743),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9641),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_9_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_9_12_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_9_12_3  (
            .in0(N__5444),
            .in1(N__5472),
            .in2(_gnd_net_),
            .in3(N__5574),
            .lcout(\U712_CHIP_RAM.N_341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_12_4 .LUT_INIT=16'b0000001001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_12_4  (
            .in0(N__6645),
            .in1(N__7147),
            .in2(N__7247),
            .in3(N__6550),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_187_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_9_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_9_12_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_9_12_5  (
            .in0(N__7745),
            .in1(N__5661),
            .in2(N__4872),
            .in3(N__7273),
            .lcout(\U712_CHIP_RAM.N_253 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_9_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_9_12_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_9_12_6  (
            .in0(N__7029),
            .in1(N__6641),
            .in2(_gnd_net_),
            .in3(N__6549),
            .lcout(\U712_CHIP_RAM.N_329 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_12_7 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_12_7  (
            .in0(N__7744),
            .in1(N__5355),
            .in2(N__6662),
            .in3(N__5662),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9641),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_1_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_1_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_1_LC_9_13_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_1_LC_9_13_0  (
            .in0(N__7248),
            .in1(N__7159),
            .in2(N__6576),
            .in3(N__6737),
            .lcout(\U712_CHIP_RAM.N_316 ),
            .ltout(\U712_CHIP_RAM.N_316_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4HBB7_2_LC_9_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4HBB7_2_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4HBB7_2_LC_9_13_1 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4HBB7_2_LC_9_13_1  (
            .in0(N__6635),
            .in1(_gnd_net_),
            .in2(N__4869),
            .in3(N__5353),
            .lcout(\U712_CHIP_RAM.N_259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_1_LC_9_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_1_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_1_LC_9_13_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_1_LC_9_13_2  (
            .in0(N__5354),
            .in1(N__5523),
            .in2(_gnd_net_),
            .in3(N__4866),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_283_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_9_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_9_13_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_9_13_3  (
            .in0(N__6738),
            .in1(N__4860),
            .in2(N__4854),
            .in3(N__5484),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_13_4 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__5544),
            .in2(N__4851),
            .in3(N__9078),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9646),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_13_5 .LUT_INIT=16'b1100000011010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_13_5  (
            .in0(N__5679),
            .in1(N__4848),
            .in2(N__8389),
            .in3(N__5505),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9646),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_9_13_6 .LUT_INIT=16'b1100111111001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__6634),
            .in2(N__6575),
            .in3(N__7392),
            .lcout(\U712_CHIP_RAM.N_184 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_13_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_13_7  (
            .in0(N__5524),
            .in1(N__6571),
            .in2(_gnd_net_),
            .in3(N__5731),
            .lcout(\U712_CHIP_RAM.N_258 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_9_14_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_9_14_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_9_14_1  (
            .in0(N__6286),
            .in1(N__5669),
            .in2(_gnd_net_),
            .in3(N__6157),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_14_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_14_2 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_9_14_2  (
            .in0(N__7404),
            .in1(N__4941),
            .in2(N__5037),
            .in3(N__7747),
            .lcout(WRITE_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9651),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_9_14_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_9_14_5 .LUT_INIT=16'b0101001100110011;
    LogicCell40 \U712_BUFFERS.DRDDIR_0_m2_LC_9_14_5  (
            .in0(N__5008),
            .in1(N__7405),
            .in2(N__10620),
            .in3(N__10543),
            .lcout(N_235),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_14_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_14_7 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_14_7  (
            .in0(N__5009),
            .in1(N__4964),
            .in2(_gnd_net_),
            .in3(N__6051),
            .lcout(\U712_CHIP_RAM.N_222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LMBE_i_o5_LC_9_15_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LMBE_i_o5_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LMBE_i_o5_LC_9_15_3 .LUT_INIT=16'b1111010001001111;
    LogicCell40 \U712_BYTE_ENABLE.LMBE_i_o5_LC_9_15_3  (
            .in0(N__8746),
            .in1(N__8843),
            .in2(N__8607),
            .in3(N__8678),
            .lcout(\U712_BYTE_ENABLE.N_217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a5_LC_9_19_7 .C_ON=1'b0;
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a5_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a5_LC_9_19_7 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \U712_BUFFERS.DMA_LATCH_EN_0_a5_LC_9_19_7  (
            .in0(N__10596),
            .in1(N__10518),
            .in2(_gnd_net_),
            .in3(N__7419),
            .lcout(DMA_LATCH_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_1  (
            .in0(N__9154),
            .in1(N__4905),
            .in2(_gnd_net_),
            .in3(N__4887),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_7_6  (
            .in0(N__5124),
            .in1(N__5109),
            .in2(_gnd_net_),
            .in3(N__9153),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_9_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_9_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__5304),
            .in2(_gnd_net_),
            .in3(N__5094),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__5069),
            .ce(),
            .sr(N__5310));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_9_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_9_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__5292),
            .in2(_gnd_net_),
            .in3(N__5091),
            .lcout(\U712_CHIP_RAM.REFRESH5lto1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__5069),
            .ce(),
            .sr(N__5310));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_9_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_9_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__5265),
            .in2(_gnd_net_),
            .in3(N__5088),
            .lcout(\U712_CHIP_RAM.REFRESH5lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__5069),
            .ce(),
            .sr(N__5310));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_9_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_9_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__5217),
            .in2(_gnd_net_),
            .in3(N__5085),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__5069),
            .ce(),
            .sr(N__5310));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_9_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_9_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__5279),
            .in2(_gnd_net_),
            .in3(N__5082),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__5069),
            .ce(),
            .sr(N__5310));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_9_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_9_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__5229),
            .in2(_gnd_net_),
            .in3(N__5079),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__5069),
            .ce(),
            .sr(N__5310));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_9_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_9_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__5241),
            .in2(_gnd_net_),
            .in3(N__5076),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__5069),
            .ce(),
            .sr(N__5310));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_9_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__5253),
            .in2(_gnd_net_),
            .in3(N__5073),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5069),
            .ce(),
            .sr(N__5310));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_10_0 .LUT_INIT=16'b0000111101111111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_10_0  (
            .in0(N__5303),
            .in1(N__5291),
            .in2(N__5280),
            .in3(N__5264),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_10_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_10_1  (
            .in0(N__5252),
            .in1(N__5240),
            .in2(_gnd_net_),
            .in3(N__5228),
            .lcout(),
            .ltout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_10_2 .LUT_INIT=16'b0000101010001010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_10_10_2  (
            .in0(N__7752),
            .in1(N__5216),
            .in2(N__5205),
            .in3(N__5202),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9632),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_11_0 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_11_0  (
            .in0(N__6049),
            .in1(_gnd_net_),
            .in2(N__5670),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_10_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_10_11_1  (
            .in0(N__7056),
            .in1(N__6739),
            .in2(N__6674),
            .in3(N__6700),
            .lcout(\U712_CHIP_RAM.N_340 ),
            .ltout(\U712_CHIP_RAM.N_340_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_11_2 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__5381),
            .in2(N__5190),
            .in3(N__5697),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_10_11_3 .LUT_INIT=16'b0000100011001000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_10_11_3  (
            .in0(N__5168),
            .in1(N__7645),
            .in2(N__5187),
            .in3(N__5184),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9635),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_10_11_5 .LUT_INIT=16'b0000000000110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_10_11_5  (
            .in0(N__7472),
            .in1(N__5816),
            .in2(N__7362),
            .in3(N__5151),
            .lcout(\U712_CYCLE_TERM.N_312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_10_11_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(N__7420),
            .in2(_gnd_net_),
            .in3(N__6572),
            .lcout(\U712_CHIP_RAM.N_206 ),
            .ltout(\U712_CHIP_RAM.N_206_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_10_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_10_11_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_10_11_7  (
            .in0(N__6661),
            .in1(N__7229),
            .in2(N__5394),
            .in3(N__5723),
            .lcout(\U712_CHIP_RAM.N_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOJRU2_1_LC_10_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOJRU2_1_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOJRU2_1_LC_10_12_0 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOJRU2_1_LC_10_12_0  (
            .in0(N__7225),
            .in1(N__5340),
            .in2(N__7155),
            .in3(N__5391),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_12_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_12_1  (
            .in0(N__6050),
            .in1(N__5647),
            .in2(_gnd_net_),
            .in3(N__6128),
            .lcout(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_12_2  (
            .in0(N__6199),
            .in1(N__6178),
            .in2(N__5961),
            .in3(N__6217),
            .lcout(\U712_CHIP_RAM.N_323 ),
            .ltout(\U712_CHIP_RAM.N_323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_12_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5364),
            .in3(N__5645),
            .lcout(\U712_CHIP_RAM.N_327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_12_4 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_12_4  (
            .in0(N__6129),
            .in1(N__5361),
            .in2(N__5328),
            .in3(N__6250),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_10_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_10_12_5  (
            .in0(N__7272),
            .in1(N__7224),
            .in2(N__7146),
            .in3(N__6554),
            .lcout(\U712_CHIP_RAM.N_378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_12_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_12_6  (
            .in0(N__5646),
            .in1(N__7271),
            .in2(_gnd_net_),
            .in3(N__7123),
            .lcout(\U712_CHIP_RAM.N_335 ),
            .ltout(\U712_CHIP_RAM.N_335_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_10_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_10_12_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_10_12_7  (
            .in0(N__5339),
            .in1(_gnd_net_),
            .in2(N__5331),
            .in3(N__7223),
            .lcout(\U712_CHIP_RAM.N_280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_10_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_10_13_0 .LUT_INIT=16'b0001001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_10_13_0  (
            .in0(N__5474),
            .in1(N__5575),
            .in2(N__5456),
            .in3(N__5604),
            .lcout(\U712_CHIP_RAM.N_284 ),
            .ltout(\U712_CHIP_RAM.N_284_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_10_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_10_13_1 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_10_13_1  (
            .in0(N__5663),
            .in1(N__5959),
            .in2(N__5478),
            .in3(N__6085),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_10_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_10_13_2 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_10_13_2  (
            .in0(N__5475),
            .in1(N__5576),
            .in2(N__5457),
            .in3(N__6035),
            .lcout(\U712_CHIP_RAM.N_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_13_3 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_13_3  (
            .in0(N__5424),
            .in1(N__5985),
            .in2(N__5415),
            .in3(N__5926),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9642),
            .ce(N__6374),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_1_LC_10_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_1_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_1_LC_10_13_4 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_1_LC_10_13_4  (
            .in0(N__7755),
            .in1(N__6302),
            .in2(_gnd_net_),
            .in3(N__6747),
            .lcout(\U712_CHIP_RAM.N_218 ),
            .ltout(\U712_CHIP_RAM.N_218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQVN9G_2_LC_10_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQVN9G_2_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQVN9G_2_LC_10_13_5 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQVN9G_2_LC_10_13_5  (
            .in0(N__6134),
            .in1(_gnd_net_),
            .in2(N__5418),
            .in3(N__5408),
            .lcout(\U712_CHIP_RAM.N_181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(N__6291),
            .in2(_gnd_net_),
            .in3(N__5664),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a2_0_a5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_13_7 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_13_7  (
            .in0(N__5973),
            .in1(N__5927),
            .in2(N__5397),
            .in3(N__6086),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9642),
            .ce(N__6374),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_10_14_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_10_14_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_10_14_0  (
            .in0(N__6650),
            .in1(N__7757),
            .in2(_gnd_net_),
            .in3(N__5667),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_i_a5_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_14_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_14_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_14_1  (
            .in0(N__6562),
            .in1(N__7280),
            .in2(N__5685),
            .in3(N__7246),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_257_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_14_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_14_2 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_14_2  (
            .in0(N__6081),
            .in1(_gnd_net_),
            .in2(N__5682),
            .in3(N__5668),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_10_14_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_10_14_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_10_14_3  (
            .in0(N__7758),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6649),
            .lcout(\U712_CHIP_RAM.N_338 ),
            .ltout(\U712_CHIP_RAM.N_338_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_14_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_14_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_14_4  (
            .in0(N__7245),
            .in1(N__6749),
            .in2(N__5673),
            .in3(N__6561),
            .lcout(\U712_CHIP_RAM.N_254 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_10_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_10_14_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_10_14_5  (
            .in0(N__5666),
            .in1(N__6028),
            .in2(_gnd_net_),
            .in3(N__6080),
            .lcout(\U712_CHIP_RAM.N_284_2 ),
            .ltout(\U712_CHIP_RAM.N_284_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_14_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_14_6 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_14_6  (
            .in0(N__5598),
            .in1(N__5580),
            .in2(N__5553),
            .in3(N__5550),
            .lcout(\U712_CHIP_RAM.N_322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_14_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_14_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_14_7  (
            .in0(N__5735),
            .in1(N__5538),
            .in2(_gnd_net_),
            .in3(N__5528),
            .lcout(\U712_CHIP_RAM.N_256 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_0 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_0  (
            .in0(N__5499),
            .in1(N__9328),
            .in2(N__9200),
            .in3(N__9471),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_8_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_8_2  (
            .in0(N__9340),
            .in1(N__9195),
            .in2(N__5493),
            .in3(N__10236),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_9_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_9_1  (
            .in0(N__5898),
            .in1(N__5880),
            .in2(_gnd_net_),
            .in3(N__9136),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_9_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_9_6  (
            .in0(N__9135),
            .in1(N__5862),
            .in2(_gnd_net_),
            .in3(N__5841),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_11_10_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_11_10_0  (
            .in0(N__6058),
            .in1(N__6261),
            .in2(_gnd_net_),
            .in3(N__6156),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9629),
            .ce(N__5745),
            .sr(N__10785));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_11_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_11_1 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_11_1  (
            .in0(N__7444),
            .in1(N__5815),
            .in2(N__5787),
            .in3(N__7644),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_211_i_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_11_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_11_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_11_2  (
            .in0(N__10844),
            .in1(_gnd_net_),
            .in2(N__5763),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.N_211_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_11_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_11_11_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__10842),
            .in2(_gnd_net_),
            .in3(N__5751),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_1_LC_11_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_1_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_1_LC_11_11_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_1_LC_11_11_4  (
            .in0(N__7216),
            .in1(N__7122),
            .in2(_gnd_net_),
            .in3(N__6564),
            .lcout(\U712_CHIP_RAM.N_339 ),
            .ltout(\U712_CHIP_RAM.N_339_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_11_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_11_11_5 .LUT_INIT=16'b0011001101011111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_11_11_5  (
            .in0(N__6740),
            .in1(N__7217),
            .in2(N__5739),
            .in3(N__6675),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_11_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_11_11_6 .LUT_INIT=16'b1111111110000101;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_11_11_6  (
            .in0(N__6676),
            .in1(N__5730),
            .in2(N__5700),
            .in3(N__5696),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_11_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_11_11_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5988),
            .in3(N__10843),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_12_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__6563),
            .in2(_gnd_net_),
            .in3(N__5979),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_12_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_12_1  (
            .in0(N__5928),
            .in1(N__7141),
            .in2(_gnd_net_),
            .in3(N__5976),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__9636),
            .ce(N__6381),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_11_12_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_11_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__6657),
            .in2(_gnd_net_),
            .in3(N__5967),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_12_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_12_3  (
            .in0(N__5929),
            .in1(N__7236),
            .in2(_gnd_net_),
            .in3(N__5964),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__9636),
            .ce(N__6381),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_12_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_12_4  (
            .in0(N__5924),
            .in1(N__5960),
            .in2(_gnd_net_),
            .in3(N__5940),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__9636),
            .ce(N__6381),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_12_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_12_5  (
            .in0(N__5930),
            .in1(N__6180),
            .in2(_gnd_net_),
            .in3(N__5937),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__9636),
            .ce(N__6381),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_12_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_12_6  (
            .in0(N__5925),
            .in1(N__6201),
            .in2(_gnd_net_),
            .in3(N__5934),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__9636),
            .ce(N__6381),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_12_7  (
            .in0(N__5931),
            .in1(N__6219),
            .in2(_gnd_net_),
            .in3(N__6384),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9636),
            .ce(N__6381),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_11_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_11_13_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_1_LC_11_13_0  (
            .in0(N__6231),
            .in1(N__10040),
            .in2(_gnd_net_),
            .in3(N__6357),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_289_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_LC_11_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.BANK0_LC_11_13_1 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \U712_CHIP_RAM.BANK0_LC_11_13_1  (
            .in0(N__6314),
            .in1(N__6267),
            .in2(N__6339),
            .in3(N__6336),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9639),
            .ce(),
            .sr(N__10771));
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_11_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_11_13_2 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_2_LC_11_13_2  (
            .in0(N__6225),
            .in1(N__6303),
            .in2(N__6290),
            .in3(N__6748),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_11_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_11_13_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_11_13_3  (
            .in0(N__6036),
            .in1(N__6260),
            .in2(_gnd_net_),
            .in3(N__6133),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_11_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_11_13_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_11_13_4  (
            .in0(N__6633),
            .in1(N__7121),
            .in2(N__7237),
            .in3(N__6538),
            .lcout(\U712_CHIP_RAM.N_331 ),
            .ltout(\U712_CHIP_RAM.N_331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_7_LC_11_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_7_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_7_LC_11_13_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_7_LC_11_13_5  (
            .in0(N__6218),
            .in1(N__6200),
            .in2(N__6183),
            .in3(N__6179),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER15 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_7_LC_11_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_7_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_7_LC_11_13_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_7_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6093),
            .in3(N__7753),
            .lcout(\U712_CHIP_RAM.N_337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_14_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_14_2 .LUT_INIT=16'b1110010011101100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_14_2  (
            .in0(N__7754),
            .in1(N__6048),
            .in2(N__6483),
            .in3(N__7057),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9643),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_11_14_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_11_14_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_11_14_4  (
            .in0(N__7412),
            .in1(N__6656),
            .in2(N__6574),
            .in3(N__9321),
            .lcout(\U712_CHIP_RAM.CPU_TACK_7_iv_i_a5_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_15_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_15_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__6474),
            .in2(_gnd_net_),
            .in3(N__6467),
            .lcout(\U712_CHIP_RAM.un3_DMA_CYCLE_START ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_15_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_15_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_11_15_7  (
            .in0(N__6468),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7756),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9647),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_16_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_16_6 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_11_16_6  (
            .in0(N__7777),
            .in1(N__10624),
            .in2(_gnd_net_),
            .in3(N__10530),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9652),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_2_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_2_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_2_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_7_5  (
            .in0(N__7518),
            .in1(N__6441),
            .in2(_gnd_net_),
            .in3(N__7524),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9618),
            .ce(N__8080),
            .sr(N__10798));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_8_1 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_12_8_1  (
            .in0(N__8266),
            .in1(N__9405),
            .in2(N__8236),
            .in3(N__6423),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9621),
            .ce(N__8082),
            .sr(N__10788));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_8_6 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_12_8_6  (
            .in0(N__8226),
            .in1(N__8267),
            .in2(N__9507),
            .in3(N__6924),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9621),
            .ce(N__8082),
            .sr(N__10788));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_9_1 .LUT_INIT=16'b0000011000000111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_9_1  (
            .in0(N__9749),
            .in1(N__9128),
            .in2(N__8465),
            .in3(N__8390),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_9_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_9_2  (
            .in0(N__9294),
            .in1(N__9149),
            .in2(N__6933),
            .in3(N__9483),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_9_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__9293),
            .in2(_gnd_net_),
            .in3(N__9129),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_10_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_10_4  (
            .in0(N__9175),
            .in1(N__6918),
            .in2(_gnd_net_),
            .in3(N__6906),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_10_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_10_5  (
            .in0(N__9346),
            .in1(N__9176),
            .in2(N__6891),
            .in3(N__9003),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_10_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_10_6  (
            .in0(N__9307),
            .in1(N__6888),
            .in2(N__9199),
            .in3(N__10209),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_10_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_10_7  (
            .in0(N__6882),
            .in1(N__9306),
            .in2(_gnd_net_),
            .in3(N__9492),
            .lcout(\U712_CHIP_RAM.N_146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pll_RNI8MQ3_LC_12_11_2.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_12_11_2.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_12_11_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 pll_RNI8MQ3_LC_12_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6865),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_12_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_12_11_4 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_12_11_4  (
            .in0(N__7058),
            .in1(N__6753),
            .in2(N__6684),
            .in3(N__6702),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_12_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_12_11_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_12_11_6  (
            .in0(N__6701),
            .in1(N__7421),
            .in2(N__6683),
            .in3(N__9314),
            .lcout(\U712_CHIP_RAM.CLK_EN_6_0_a5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_12_11_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_12_11_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_12_11_7  (
            .in0(N__7471),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7352),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_12_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_12_12_6 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_LC_12_12_6  (
            .in0(N__9359),
            .in1(N__7145),
            .in2(N__7068),
            .in3(N__7422),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9631),
            .ce(N__7341),
            .sr(N__10769));
    defparam \U712_BYTE_ENABLE.N_118_i_LC_12_13_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_118_i_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_118_i_LC_12_13_0 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \U712_BYTE_ENABLE.N_118_i_LC_12_13_0  (
            .in0(N__10629),
            .in1(N__6962),
            .in2(N__6954),
            .in3(N__9387),
            .lcout(N_118_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_119_i_LC_12_13_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_119_i_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_119_i_LC_12_13_4 .LUT_INIT=16'b0101000111110011;
    LogicCell40 \U712_BYTE_ENABLE.N_119_i_LC_12_13_4  (
            .in0(N__6942),
            .in1(N__6963),
            .in2(N__10545),
            .in3(N__9388),
            .lcout(N_119_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_12_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_12_13_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_12_13_6  (
            .in0(N__7284),
            .in1(N__7235),
            .in2(N__7161),
            .in3(N__7074),
            .lcout(\U712_CHIP_RAM.N_287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a5_0_0_LC_12_13_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a5_0_0_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a5_0_0_LC_12_13_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a5_0_0_LC_12_13_7  (
            .in0(N__7059),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6998),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_a5_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UUBE_0_a2_LC_12_15_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UUBE_0_a2_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UUBE_0_a2_LC_12_15_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BYTE_ENABLE.UUBE_0_a2_LC_12_15_3  (
            .in0(N__8766),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8850),
            .lcout(\U712_BYTE_ENABLE.UUBE ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_i_o5_LC_12_16_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_i_o5_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_i_o5_LC_12_16_2 .LUT_INIT=16'b1111010101001111;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_i_o5_LC_12_16_2  (
            .in0(N__8842),
            .in1(N__8732),
            .in2(N__8685),
            .in3(N__8605),
            .lcout(\U712_BYTE_ENABLE.N_216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_6.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_6.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_18_6 (
            .in0(N__7742),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_12_20_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_12_20_7 .LUT_INIT=16'b0001000011111111;
    LogicCell40 \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_12_20_7  (
            .in0(N__8767),
            .in1(N__8579),
            .in2(N__8668),
            .in3(N__7838),
            .lcout(N_163),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_6_5 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_13_6_5  (
            .in0(N__8148),
            .in1(N__7563),
            .in2(N__9389),
            .in3(N__10428),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9619),
            .ce(N__8073),
            .sr(N__10813));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_7_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__9751),
            .in2(_gnd_net_),
            .in3(N__8404),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_7_1 .LUT_INIT=16'b0000010011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_7_1  (
            .in0(N__9371),
            .in1(N__8909),
            .in2(N__7527),
            .in3(N__9181),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_7_7 .LUT_INIT=16'b0000111011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_7_7  (
            .in0(N__9370),
            .in1(N__8910),
            .in2(N__8230),
            .in3(N__9180),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_8_6 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_8_6  (
            .in0(N__9204),
            .in1(N__8219),
            .in2(_gnd_net_),
            .in3(N__7512),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_8_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(N__7479),
            .in2(N__7503),
            .in3(N__7992),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9623),
            .ce(N__8085),
            .sr(N__10802));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_13_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_13_9_2 .LUT_INIT=16'b1101111111010101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_13_9_2  (
            .in0(N__8143),
            .in1(N__8016),
            .in2(N__9391),
            .in3(N__9528),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_9_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_9_3  (
            .in0(N__9750),
            .in1(N__9173),
            .in2(_gnd_net_),
            .in3(N__8403),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(\U712_CHIP_RAM.CMA_5_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_9_4 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_9_4  (
            .in0(N__9378),
            .in1(N__8015),
            .in2(N__7995),
            .in3(N__9527),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_9_6 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_9_6  (
            .in0(N__10847),
            .in1(N__7986),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_9_7  (
            .in0(N__7980),
            .in1(N__7959),
            .in2(_gnd_net_),
            .in3(N__9174),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_10_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_13_10_3  (
            .in0(N__8268),
            .in1(N__7851),
            .in2(N__8241),
            .in3(N__7941),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9630),
            .ce(N__8084),
            .sr(N__10786));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_10_4 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_13_10_4  (
            .in0(N__8234),
            .in1(N__8269),
            .in2(N__10131),
            .in3(N__7920),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9630),
            .ce(N__8084),
            .sr(N__10786));
    defparam \U712_CHIP_RAM.CLK_EN_LC_13_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_13_11_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_13_11_6 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_13_11_6  (
            .in0(N__7862),
            .in1(N__7893),
            .in2(_gnd_net_),
            .in3(N__7887),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9633),
            .ce(),
            .sr(N__10774));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_12_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_12_6  (
            .in0(N__8943),
            .in1(N__8991),
            .in2(_gnd_net_),
            .in3(N__10050),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9858),
            .ce(N__9817),
            .sr(N__10772));
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_LC_13_20_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_LC_13_20_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U712_BYTE_ENABLE.un1_UDSn_i_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(N__8768),
            .in2(_gnd_net_),
            .in3(N__7842),
            .lcout(U712_BYTE_ENABLE_un1_UDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WEn_LC_14_1_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_14_1_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_14_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_14_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8405),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9616),
            .ce(),
            .sr(N__10821));
    defparam \U712_CHIP_RAM.CASn_LC_14_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_14_4_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_14_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_14_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9203),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9617),
            .ce(),
            .sr(N__10819));
    defparam \U712_CHIP_RAM.CRCSn_LC_14_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_14_5_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_14_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_14_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8466),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9620),
            .ce(),
            .sr(N__10818));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_7  (
            .in0(N__9365),
            .in1(N__8475),
            .in2(N__9201),
            .in3(N__10332),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_7_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_14_7_3  (
            .in0(N__8464),
            .in1(N__9194),
            .in2(N__9764),
            .in3(N__8406),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9624),
            .ce(N__8081),
            .sr(N__10814));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_7_6 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_14_7_6  (
            .in0(N__8283),
            .in1(N__9516),
            .in2(N__8235),
            .in3(N__8310),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9624),
            .ce(N__8081),
            .sr(N__10814));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_8_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_14_8_0  (
            .in0(N__8282),
            .in1(N__9012),
            .in2(N__8237),
            .in3(N__9018),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9625),
            .ce(N__8083),
            .sr(N__10806));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_8_5 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_14_8_5  (
            .in0(N__8144),
            .in1(N__8127),
            .in2(N__9393),
            .in3(N__9867),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9625),
            .ce(N__8083),
            .sr(N__10806));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_9_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_9_7  (
            .in0(N__9390),
            .in1(N__9210),
            .in2(N__9202),
            .in3(N__10221),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_10_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_10_3  (
            .in0(N__10197),
            .in1(N__9967),
            .in2(_gnd_net_),
            .in3(N__10371),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9853),
            .ce(N__9819),
            .sr(N__10790));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_11_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_11_2  (
            .in0(N__8939),
            .in1(N__10044),
            .in2(_gnd_net_),
            .in3(N__9458),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__9816),
            .sr(N__10787));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_14_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_14_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_14_11_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_14_11_4  (
            .in0(N__8938),
            .in1(N__10043),
            .in2(_gnd_net_),
            .in3(N__8990),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__9816),
            .sr(N__10787));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_12_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_12_7  (
            .in0(N__9444),
            .in1(N__9993),
            .in2(_gnd_net_),
            .in3(N__8937),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9857),
            .ce(N__9820),
            .sr(N__10775));
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_14_19_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_14_19_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_BYTE_ENABLE.UUBE_i_LC_14_19_2  (
            .in0(N__8822),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8769),
            .lcout(U712_BYTE_ENABLE_UUBE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_215_i_LC_14_20_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_215_i_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_215_i_LC_14_20_0 .LUT_INIT=16'b0000010101110000;
    LogicCell40 \U712_BYTE_ENABLE.N_215_i_LC_14_20_0  (
            .in0(N__8847),
            .in1(N__8770),
            .in2(N__8682),
            .in3(N__8596),
            .lcout(N_215_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_217_i_LC_14_20_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_217_i_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_217_i_LC_14_20_2 .LUT_INIT=16'b0000110111010000;
    LogicCell40 \U712_BYTE_ENABLE.N_217_i_LC_14_20_2  (
            .in0(N__8849),
            .in1(N__8772),
            .in2(N__8684),
            .in3(N__8598),
            .lcout(N_217_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_216_i_LC_14_20_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_216_i_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_216_i_LC_14_20_6 .LUT_INIT=16'b0000101010110000;
    LogicCell40 \U712_BYTE_ENABLE.N_216_i_LC_14_20_6  (
            .in0(N__8848),
            .in1(N__8771),
            .in2(N__8683),
            .in3(N__8597),
            .lcout(N_216_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RASn_LC_15_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_15_5_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_15_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_15_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9765),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9622),
            .ce(),
            .sr(N__10820));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_9_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_9_3  (
            .in0(N__10416),
            .in1(N__10039),
            .in2(_gnd_net_),
            .in3(N__10369),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9854),
            .ce(N__9823),
            .sr(N__10807));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_9_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_9_4  (
            .in0(N__10320),
            .in1(_gnd_net_),
            .in2(N__10049),
            .in3(N__10415),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9854),
            .ce(N__9823),
            .sr(N__10807));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_9_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_9_5  (
            .in0(N__10284),
            .in1(N__10035),
            .in2(_gnd_net_),
            .in3(N__10319),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9854),
            .ce(N__9823),
            .sr(N__10807));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_10_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_10_4  (
            .in0(N__10034),
            .in1(N__10196),
            .in2(_gnd_net_),
            .in3(N__10370),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__9822),
            .sr(N__10803));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_10_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_10_5  (
            .in0(N__10313),
            .in1(N__10033),
            .in2(_gnd_net_),
            .in3(N__10408),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__9822),
            .sr(N__10803));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_10_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_10_7  (
            .in0(N__9459),
            .in1(N__10032),
            .in2(_gnd_net_),
            .in3(N__10283),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__9822),
            .sr(N__10803));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_11_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_11_2  (
            .in0(N__9457),
            .in1(N__10042),
            .in2(_gnd_net_),
            .in3(N__10275),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9855),
            .ce(N__9818),
            .sr(N__10791));
    defparam \U712_CHIP_RAM.DMA_A20_LC_15_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A20_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A20_LC_15_13_3 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A20_LC_15_13_3  (
            .in0(N__9992),
            .in1(N__10464),
            .in2(N__10118),
            .in3(N__10442),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .ce(),
            .sr(N__10776));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_8_3  (
            .in0(N__10031),
            .in1(N__10119),
            .in2(_gnd_net_),
            .in3(N__10167),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9856),
            .ce(N__9827),
            .sr(N__10817));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_16_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_16_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_16_9_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_16_9_6  (
            .in0(N__10414),
            .in1(_gnd_net_),
            .in2(N__10048),
            .in3(N__10362),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__9825),
            .sr(N__10815));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_16_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_16_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_16_9_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_16_9_7  (
            .in0(N__10306),
            .in1(N__10027),
            .in2(_gnd_net_),
            .in3(N__10282),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__9825),
            .sr(N__10815));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_16_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_16_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_16_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_16_10_5  (
            .in0(N__10165),
            .in1(N__10195),
            .in2(_gnd_net_),
            .in3(N__10026),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__9824),
            .sr(N__10808));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_11_7  (
            .in0(N__9944),
            .in1(N__10114),
            .in2(_gnd_net_),
            .in3(N__10166),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__9821),
            .sr(N__10804));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_10_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_10_6  (
            .in0(N__10194),
            .in1(N__10041),
            .in2(_gnd_net_),
            .in3(N__10164),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9852),
            .ce(N__9826),
            .sr(N__10816));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_8_5  (
            .in0(N__10093),
            .in1(N__10059),
            .in2(_gnd_net_),
            .in3(N__10011),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9851),
            .ce(N__9828),
            .sr(N__10822));
    defparam \U712_BUFFERS.un1_DRDENn_0_a5_LC_24_19_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a5_LC_24_19_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a5_LC_24_19_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a5_LC_24_19_5  (
            .in0(N__10674),
            .in1(N__10581),
            .in2(_gnd_net_),
            .in3(N__10499),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

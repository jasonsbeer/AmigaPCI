-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     May 31 2025 14:05:17

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    TT : in std_logic_vector(1 downto 0);
    TM : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(31 downto 1);
    D : out std_logic_vector(7 downto 0);
    TICK60 : out std_logic;
    CIACS0n : out std_logic;
    CLK6 : in std_logic;
    CLK_CIA : out std_logic;
    BUFENn : out std_logic;
    RnW : in std_logic;
    CIACS1n : out std_logic;
    TICK50 : out std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : out std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    REGSPACEn : out std_logic;
    TSn : in std_logic;
    RTC_ENn : out std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    TACKn : inout std_logic;
    ROMENn : out std_logic;
    PORTSIZE : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__7928\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2920\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_26\ : std_logic;
signal \A_c_25\ : std_logic;
signal \A_c_24\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_\ : std_logic;
signal \A_c_31\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_28\ : std_logic;
signal \A_c_29\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACE_0Z0Z_1_cascade_\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_5\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_0_cascade_\ : std_logic;
signal \RnW_c\ : std_logic;
signal \D_1_i\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RTC_ENn_i\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5\ : std_logic;
signal \U409_ADDRESS_DECODE_LOWROM_3_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOVECTOR_3\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOVECTOR_2\ : std_logic;
signal \U409_ADDRESS_DECODE_LOWROM_2_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_45\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2Z0Z_1_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_20\ : std_logic;
signal \A_c_19\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_\ : std_logic;
signal \TM_c_1\ : std_logic;
signal \TM_c_0\ : std_logic;
signal \A_c_23\ : std_logic;
signal \A_c_22\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn_i\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.un2_REGSPACEn_0_0\ : std_logic;
signal \U409_ADDRESS_DECODE.REG_SPACE_3_0\ : std_logic;
signal \U409_ADDRESS_DECODE.REG_SPACEZ0Z_2\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RTC_ENn\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_OUTnC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6\ : std_logic;
signal \U409_TRANSFER_ACK.N_35\ : std_logic;
signal \ROMENn_c\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_47\ : std_logic;
signal \U409_TRANSFER_ACK.N_142\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\ : std_logic;
signal \A_c_21\ : std_logic;
signal \OVL_c\ : std_logic;
signal \U409_ADDRESS_DECODE_LOWROM_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_2_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5\ : std_logic;
signal \U409_ADDRESS_DECODE_ROMEN_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_23\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_1_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_35_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_29\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.N_36\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn\ : std_logic;
signal \BUFENn_c\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.i6_mux_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_9_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TRANSFER_ACK.N_4\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_5\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \U409_TRANSFER_ACK.m8_ns_1\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.TICK603_8\ : std_logic;
signal \U409_TICK.TICK603_11_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.TICK603_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_0C_net\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \AUTOCONFIG_SPACE\ : std_logic;
signal \TCIn_1_i\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS1n_i\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \CIA_ENABLE\ : std_logic;
signal \A_c_12\ : std_logic;
signal \CIA_ENABLE_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS0n_i\ : std_logic;
signal \U409_TICK.TICK503_11_cascade_\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \U409_TICK.TICK503_8\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \U409_CIA.CLK_CIA6_3_cascade_\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_\ : std_logic;
signal \CIA_SPACE\ : std_logic;
signal \U409_CIA.VMA_RNOZ0Z_0_cascade_\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \CLK_CIA_c\ : std_logic;
signal \U409_CIA.CLK_CIA_r_1_0\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_0\ : std_logic;
signal \U409_CIA.CLK_CIA6_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_6\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_5\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_6\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_7\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \D_wire\ : std_logic_vector(7 downto 0);
signal \RTC_ENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \TM_wire\ : std_logic_vector(1 downto 0);
signal \CLK_CIA_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \ROMENn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \CIACS0n_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \CIACS1n_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    \TT_wire\ <= TT;
    D <= \D_wire\;
    RTC_ENn <= \RTC_ENn_wire\;
    \A_wire\ <= A;
    \TM_wire\ <= TM;
    CLK_CIA <= \CLK_CIA_wire\;
    RAMSPACEn <= \RAMSPACEn_wire\;
    ROMENn <= \ROMENn_wire\;
    TBIn <= \TBIn_wire\;
    \TSn_wire\ <= TSn;
    BUFENn <= \BUFENn_wire\;
    PORTSIZE <= \PORTSIZE_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    CIACS0n <= \CIACS0n_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TCIn <= \TCIn_wire\;
    \RnW_wire\ <= RnW;
    TICK60 <= \TICK60_wire\;
    CIACS1n <= \CIACS1n_wire\;
    REGSPACEn <= \REGSPACEn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__5548\,
            RESETB => \N__4699\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__7926\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7928\,
            DIN => \N__7927\,
            DOUT => \N__7926\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7928\,
            PADOUT => \N__7927\,
            PADIN => \N__7926\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__7916\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7918\,
            DIN => \N__7917\,
            DOUT => \N__7916\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7918\,
            PADOUT => \N__7917\,
            PADIN => \N__7916\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7907\,
            DIN => \N__7906\,
            DOUT => \N__7905\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7907\,
            PADOUT => \N__7906\,
            PADIN => \N__7905\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7898\,
            DIN => \N__7897\,
            DOUT => \N__7896\,
            PACKAGEPIN => \D_wire\(6)
        );

    \D_obuft_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7898\,
            PADOUT => \N__7897\,
            PADIN => \N__7896\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3324\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RTC_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7889\,
            DIN => \N__7888\,
            DOUT => \N__7887\,
            PACKAGEPIN => \RTC_ENn_wire\
        );

    \RTC_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7889\,
            PADOUT => \N__7888\,
            PADIN => \N__7887\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3253\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7880\,
            DIN => \N__7879\,
            DOUT => \N__7878\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7880\,
            PADOUT => \N__7879\,
            PADIN => \N__7878\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7871\,
            DIN => \N__7870\,
            DOUT => \N__7869\,
            PACKAGEPIN => \D_wire\(5)
        );

    \D_obuft_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7871\,
            PADOUT => \N__7870\,
            PADIN => \N__7869\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3323\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7862\,
            DIN => \N__7861\,
            DOUT => \N__7860\,
            PACKAGEPIN => \TM_wire\(1)
        );

    \TM_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7862\,
            PADOUT => \N__7861\,
            PADIN => \N__7860\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7853\,
            DIN => \N__7852\,
            DOUT => \N__7851\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7853\,
            PADOUT => \N__7852\,
            PADIN => \N__7851\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_CIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7844\,
            DIN => \N__7843\,
            DOUT => \N__7842\,
            PACKAGEPIN => \CLK_CIA_wire\
        );

    \CLK_CIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7844\,
            PADOUT => \N__7843\,
            PADIN => \N__7842\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7183\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7835\,
            DIN => \N__7834\,
            DOUT => \N__7833\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7835\,
            PADOUT => \N__7834\,
            PADIN => \N__7833\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7826\,
            DIN => \N__7825\,
            DOUT => \N__7824\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7826\,
            PADOUT => \N__7825\,
            PADIN => \N__7824\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4468\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7817\,
            DIN => \N__7816\,
            DOUT => \N__7815\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7817\,
            PADOUT => \N__7816\,
            PADIN => \N__7815\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6378\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__4243\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7808\,
            DIN => \N__7807\,
            DOUT => \N__7806\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7808\,
            PADOUT => \N__7807\,
            PADIN => \N__7806\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7799\,
            DIN => \N__7798\,
            DOUT => \N__7797\,
            PACKAGEPIN => \ROMENn_wire\
        );

    \ROMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7799\,
            PADOUT => \N__7798\,
            PADIN => \N__7797\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4123\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7790\,
            DIN => \N__7789\,
            DOUT => \N__7788\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7790\,
            PADOUT => \N__7789\,
            PADIN => \N__7788\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6382\,
            DIN0 => OPEN,
            DOUT0 => \N__4238\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7781\,
            DIN => \N__7780\,
            DOUT => \N__7779\,
            PACKAGEPIN => \D_wire\(0)
        );

    \D_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7781\,
            PADOUT => \N__7780\,
            PADIN => \N__7779\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3308\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7772\,
            DIN => \N__7771\,
            DOUT => \N__7770\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7772\,
            PADOUT => \N__7771\,
            PADIN => \N__7770\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7763\,
            DIN => \N__7762\,
            DOUT => \N__7761\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7763\,
            PADOUT => \N__7762\,
            PADIN => \N__7761\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7754\,
            DIN => \N__7753\,
            DOUT => \N__7752\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7754\,
            PADOUT => \N__7753\,
            PADIN => \N__7752\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5389\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7745\,
            DIN => \N__7744\,
            DOUT => \N__7743\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7745\,
            PADOUT => \N__7744\,
            PADIN => \N__7743\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3751\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7736\,
            DIN => \N__7735\,
            DOUT => \N__7734\,
            PACKAGEPIN => \D_wire\(7)
        );

    \D_obuft_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7736\,
            PADOUT => \N__7735\,
            PADIN => \N__7734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3328\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7727\,
            DIN => \N__7726\,
            DOUT => \N__7725\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7727\,
            PADOUT => \N__7726\,
            PADIN => \N__7725\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7718\,
            DIN => \N__7717\,
            DOUT => \N__7716\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7718\,
            PADOUT => \N__7717\,
            PADIN => \N__7716\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7709\,
            DIN => \N__7708\,
            DOUT => \N__7707\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7709\,
            PADOUT => \N__7708\,
            PADIN => \N__7707\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7700\,
            DIN => \N__7699\,
            DOUT => \N__7698\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7700\,
            PADOUT => \N__7699\,
            PADIN => \N__7698\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7691\,
            DIN => \N__7690\,
            DOUT => \N__7689\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7691\,
            PADOUT => \N__7690\,
            PADIN => \N__7689\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7682\,
            DIN => \N__7681\,
            DOUT => \N__7680\,
            PACKAGEPIN => \D_wire\(2)
        );

    \D_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7682\,
            PADOUT => \N__7681\,
            PADIN => \N__7680\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3275\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7673\,
            DIN => \N__7672\,
            DOUT => \N__7671\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7673\,
            PADOUT => \N__7672\,
            PADIN => \N__7671\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7664\,
            DIN => \N__7663\,
            DOUT => \N__7662\,
            PACKAGEPIN => \TM_wire\(0)
        );

    \TM_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7664\,
            PADOUT => \N__7663\,
            PADIN => \N__7662\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7655\,
            DIN => \N__7654\,
            DOUT => \N__7653\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7655\,
            PADOUT => \N__7654\,
            PADIN => \N__7653\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7646\,
            DIN => \N__7645\,
            DOUT => \N__7644\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7646\,
            PADOUT => \N__7645\,
            PADIN => \N__7644\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7637\,
            DIN => \N__7636\,
            DOUT => \N__7635\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7637\,
            PADOUT => \N__7636\,
            PADIN => \N__7635\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7628\,
            DIN => \N__7627\,
            DOUT => \N__7626\,
            PACKAGEPIN => \D_wire\(1)
        );

    \D_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7628\,
            PADOUT => \N__7627\,
            PADIN => \N__7626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3307\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7619\,
            DIN => \N__7618\,
            DOUT => \N__7617\,
            PACKAGEPIN => \CIACS0n_wire\
        );

    \CIACS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7619\,
            PADOUT => \N__7618\,
            PADIN => \N__7617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6088\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7610\,
            DIN => \N__7609\,
            DOUT => \N__7608\,
            PACKAGEPIN => \D_wire\(4)
        );

    \D_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7610\,
            PADOUT => \N__7609\,
            PADIN => \N__7608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3322\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7601\,
            DIN => \N__7600\,
            DOUT => \N__7599\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7601\,
            PADOUT => \N__7600\,
            PADIN => \N__7599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7138\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7592\,
            DIN => \N__7591\,
            DOUT => \N__7590\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7592\,
            PADOUT => \N__7591\,
            PADIN => \N__7590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7583\,
            DIN => \N__7582\,
            DOUT => \N__7581\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7583\,
            PADOUT => \N__7582\,
            PADIN => \N__7581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7574\,
            DIN => \N__7573\,
            DOUT => \N__7572\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7574\,
            PADOUT => \N__7573\,
            PADIN => \N__7572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7565\,
            DIN => \N__7564\,
            DOUT => \N__7563\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7565\,
            PADOUT => \N__7564\,
            PADIN => \N__7563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7556\,
            DIN => \N__7555\,
            DOUT => \N__7554\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7556\,
            PADOUT => \N__7555\,
            PADIN => \N__7554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6295\,
            DIN0 => OPEN,
            DOUT0 => \N__4239\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7547\,
            DIN => \N__7546\,
            DOUT => \N__7545\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7547\,
            PADOUT => \N__7546\,
            PADIN => \N__7545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7538\,
            DIN => \N__7537\,
            DOUT => \N__7536\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7538\,
            PADOUT => \N__7537\,
            PADIN => \N__7536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7529\,
            DIN => \N__7528\,
            DOUT => \N__7527\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7529\,
            PADOUT => \N__7528\,
            PADIN => \N__7527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5662\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7520\,
            DIN => \N__7519\,
            DOUT => \N__7518\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7520\,
            PADOUT => \N__7519\,
            PADIN => \N__7518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7511\,
            DIN => \N__7510\,
            DOUT => \N__7509\,
            PACKAGEPIN => \D_wire\(3)
        );

    \D_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7511\,
            PADOUT => \N__7510\,
            PADIN => \N__7509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3309\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7502\,
            DIN => \N__7501\,
            DOUT => \N__7500\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7502\,
            PADOUT => \N__7501\,
            PADIN => \N__7500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7493\,
            DIN => \N__7492\,
            DOUT => \N__7491\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7493\,
            PADOUT => \N__7492\,
            PADIN => \N__7491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7484\,
            DIN => \N__7483\,
            DOUT => \N__7482\,
            PACKAGEPIN => \CIACS1n_wire\
        );

    \CIACS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7484\,
            PADOUT => \N__7483\,
            PADIN => \N__7482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6265\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7475\,
            DIN => \N__7474\,
            DOUT => \N__7473\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7475\,
            PADOUT => \N__7474\,
            PADIN => \N__7473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3883\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1767\ : InMux
    port map (
            O => \N__7456\,
            I => \N__7451\
        );

    \I__1766\ : InMux
    port map (
            O => \N__7455\,
            I => \N__7448\
        );

    \I__1765\ : InMux
    port map (
            O => \N__7454\,
            I => \N__7445\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__7451\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__7448\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__7445\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1761\ : InMux
    port map (
            O => \N__7438\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\
        );

    \I__1760\ : InMux
    port map (
            O => \N__7435\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\
        );

    \I__1759\ : InMux
    port map (
            O => \N__7432\,
            I => \N__7427\
        );

    \I__1758\ : InMux
    port map (
            O => \N__7431\,
            I => \N__7422\
        );

    \I__1757\ : InMux
    port map (
            O => \N__7430\,
            I => \N__7422\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__7427\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__7422\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__7417\,
            I => \N__7409\
        );

    \I__1753\ : InMux
    port map (
            O => \N__7416\,
            I => \N__7406\
        );

    \I__1752\ : InMux
    port map (
            O => \N__7415\,
            I => \N__7403\
        );

    \I__1751\ : InMux
    port map (
            O => \N__7414\,
            I => \N__7398\
        );

    \I__1750\ : InMux
    port map (
            O => \N__7413\,
            I => \N__7398\
        );

    \I__1749\ : InMux
    port map (
            O => \N__7412\,
            I => \N__7393\
        );

    \I__1748\ : InMux
    port map (
            O => \N__7409\,
            I => \N__7393\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__7406\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__7403\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__7398\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__7393\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1743\ : ClkMux
    port map (
            O => \N__7384\,
            I => \N__7375\
        );

    \I__1742\ : ClkMux
    port map (
            O => \N__7383\,
            I => \N__7375\
        );

    \I__1741\ : ClkMux
    port map (
            O => \N__7382\,
            I => \N__7375\
        );

    \I__1740\ : GlobalMux
    port map (
            O => \N__7375\,
            I => \N__7372\
        );

    \I__1739\ : gio2CtrlBuf
    port map (
            O => \N__7372\,
            I => \CLK28_IN_c_g\
        );

    \I__1738\ : InMux
    port map (
            O => \N__7369\,
            I => \N__7366\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__7366\,
            I => \U409_CIA.CIA_CLK_COUNT11_2\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__7363\,
            I => \N__7360\
        );

    \I__1735\ : InMux
    port map (
            O => \N__7360\,
            I => \N__7356\
        );

    \I__1734\ : InMux
    port map (
            O => \N__7359\,
            I => \N__7353\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__7356\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__7353\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0\
        );

    \I__1731\ : InMux
    port map (
            O => \N__7348\,
            I => \N__7341\
        );

    \I__1730\ : InMux
    port map (
            O => \N__7347\,
            I => \N__7341\
        );

    \I__1729\ : InMux
    port map (
            O => \N__7346\,
            I => \N__7338\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__7341\,
            I => \U409_CIA.CLK_CIA6_4\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__7338\,
            I => \U409_CIA.CLK_CIA6_4\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__7333\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_cascade_\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__7330\,
            I => \N__7327\
        );

    \I__1724\ : InMux
    port map (
            O => \N__7327\,
            I => \N__7319\
        );

    \I__1723\ : InMux
    port map (
            O => \N__7326\,
            I => \N__7314\
        );

    \I__1722\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7314\
        );

    \I__1721\ : InMux
    port map (
            O => \N__7324\,
            I => \N__7309\
        );

    \I__1720\ : InMux
    port map (
            O => \N__7323\,
            I => \N__7309\
        );

    \I__1719\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7306\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__7319\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__7314\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__7309\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__7306\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1714\ : InMux
    port map (
            O => \N__7297\,
            I => \N__7291\
        );

    \I__1713\ : InMux
    port map (
            O => \N__7296\,
            I => \N__7286\
        );

    \I__1712\ : InMux
    port map (
            O => \N__7295\,
            I => \N__7286\
        );

    \I__1711\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7283\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__7291\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__7286\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__7283\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1707\ : InMux
    port map (
            O => \N__7276\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__1706\ : InMux
    port map (
            O => \N__7273\,
            I => \N__7267\
        );

    \I__1705\ : InMux
    port map (
            O => \N__7272\,
            I => \N__7262\
        );

    \I__1704\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7262\
        );

    \I__1703\ : InMux
    port map (
            O => \N__7270\,
            I => \N__7259\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__7267\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__7262\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__7259\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1699\ : InMux
    port map (
            O => \N__7252\,
            I => \N__7249\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__7249\,
            I => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3\
        );

    \I__1697\ : InMux
    port map (
            O => \N__7246\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__1696\ : InMux
    port map (
            O => \N__7243\,
            I => \N__7235\
        );

    \I__1695\ : InMux
    port map (
            O => \N__7242\,
            I => \N__7235\
        );

    \I__1694\ : InMux
    port map (
            O => \N__7241\,
            I => \N__7232\
        );

    \I__1693\ : InMux
    port map (
            O => \N__7240\,
            I => \N__7229\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__7235\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__7232\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__7229\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1689\ : InMux
    port map (
            O => \N__7222\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__7219\,
            I => \N__7215\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__7218\,
            I => \N__7210\
        );

    \I__1686\ : InMux
    port map (
            O => \N__7215\,
            I => \N__7207\
        );

    \I__1685\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7204\
        );

    \I__1684\ : InMux
    port map (
            O => \N__7213\,
            I => \N__7199\
        );

    \I__1683\ : InMux
    port map (
            O => \N__7210\,
            I => \N__7199\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__7207\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__7204\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__7199\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1679\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7189\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__7189\,
            I => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5\
        );

    \I__1677\ : InMux
    port map (
            O => \N__7186\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__1676\ : IoInMux
    port map (
            O => \N__7183\,
            I => \N__7180\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__7180\,
            I => \N__7177\
        );

    \I__1674\ : Span4Mux_s3_v
    port map (
            O => \N__7177\,
            I => \N__7174\
        );

    \I__1673\ : Span4Mux_v
    port map (
            O => \N__7174\,
            I => \N__7171\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__7171\,
            I => \N__7167\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__7170\,
            I => \N__7162\
        );

    \I__1670\ : Span4Mux_v
    port map (
            O => \N__7167\,
            I => \N__7159\
        );

    \I__1669\ : InMux
    port map (
            O => \N__7166\,
            I => \N__7156\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7165\,
            I => \N__7151\
        );

    \I__1667\ : InMux
    port map (
            O => \N__7162\,
            I => \N__7151\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__7159\,
            I => \CLK_CIA_c\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__7156\,
            I => \CLK_CIA_c\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__7151\,
            I => \CLK_CIA_c\
        );

    \I__1663\ : InMux
    port map (
            O => \N__7144\,
            I => \N__7141\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7141\,
            I => \U409_CIA.CLK_CIA_r_1_0\
        );

    \I__1661\ : IoInMux
    port map (
            O => \N__7138\,
            I => \N__7135\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7135\,
            I => \N__7132\
        );

    \I__1659\ : Span4Mux_s3_v
    port map (
            O => \N__7132\,
            I => \N__7129\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__7129\,
            I => \N__7126\
        );

    \I__1657\ : Span4Mux_v
    port map (
            O => \N__7126\,
            I => \N__7123\
        );

    \I__1656\ : Span4Mux_h
    port map (
            O => \N__7123\,
            I => \N__7119\
        );

    \I__1655\ : InMux
    port map (
            O => \N__7122\,
            I => \N__7116\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__7119\,
            I => \TICK50_c\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__7116\,
            I => \TICK50_c\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__7111\,
            I => \N__7108\
        );

    \I__1651\ : InMux
    port map (
            O => \N__7108\,
            I => \N__7105\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__7105\,
            I => \N__7102\
        );

    \I__1649\ : Span4Mux_h
    port map (
            O => \N__7102\,
            I => \N__7099\
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__7099\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__7096\,
            I => \N__7093\
        );

    \I__1646\ : InMux
    port map (
            O => \N__7093\,
            I => \N__7089\
        );

    \I__1645\ : InMux
    port map (
            O => \N__7092\,
            I => \N__7086\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7089\,
            I => \N__7083\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7086\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__7083\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1641\ : InMux
    port map (
            O => \N__7078\,
            I => \N__7075\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__7075\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__1639\ : InMux
    port map (
            O => \N__7072\,
            I => \N__7068\
        );

    \I__1638\ : InMux
    port map (
            O => \N__7071\,
            I => \N__7065\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__7068\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__7065\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1635\ : InMux
    port map (
            O => \N__7060\,
            I => \N__7056\
        );

    \I__1634\ : InMux
    port map (
            O => \N__7059\,
            I => \N__7053\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7056\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__7053\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__7048\,
            I => \N__7045\
        );

    \I__1630\ : InMux
    port map (
            O => \N__7045\,
            I => \N__7041\
        );

    \I__1629\ : InMux
    port map (
            O => \N__7044\,
            I => \N__7038\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__7041\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__7038\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__7033\,
            I => \N__7027\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__7032\,
            I => \N__7024\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__7031\,
            I => \N__7020\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__7030\,
            I => \N__7015\
        );

    \I__1622\ : InMux
    port map (
            O => \N__7027\,
            I => \N__7011\
        );

    \I__1621\ : InMux
    port map (
            O => \N__7024\,
            I => \N__7008\
        );

    \I__1620\ : InMux
    port map (
            O => \N__7023\,
            I => \N__7003\
        );

    \I__1619\ : InMux
    port map (
            O => \N__7020\,
            I => \N__7003\
        );

    \I__1618\ : InMux
    port map (
            O => \N__7019\,
            I => \N__6994\
        );

    \I__1617\ : InMux
    port map (
            O => \N__7018\,
            I => \N__6994\
        );

    \I__1616\ : InMux
    port map (
            O => \N__7015\,
            I => \N__6994\
        );

    \I__1615\ : InMux
    port map (
            O => \N__7014\,
            I => \N__6994\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__7011\,
            I => \N__6991\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__7008\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__7003\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__6994\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1610\ : Odrv4
    port map (
            O => \N__6991\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1609\ : InMux
    port map (
            O => \N__6982\,
            I => \N__6972\
        );

    \I__1608\ : InMux
    port map (
            O => \N__6981\,
            I => \N__6967\
        );

    \I__1607\ : InMux
    port map (
            O => \N__6980\,
            I => \N__6967\
        );

    \I__1606\ : InMux
    port map (
            O => \N__6979\,
            I => \N__6962\
        );

    \I__1605\ : InMux
    port map (
            O => \N__6978\,
            I => \N__6962\
        );

    \I__1604\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6955\
        );

    \I__1603\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6955\
        );

    \I__1602\ : InMux
    port map (
            O => \N__6975\,
            I => \N__6955\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__6972\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__6967\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__6962\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__6955\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1597\ : InMux
    port map (
            O => \N__6946\,
            I => \N__6932\
        );

    \I__1596\ : InMux
    port map (
            O => \N__6945\,
            I => \N__6932\
        );

    \I__1595\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6932\
        );

    \I__1594\ : InMux
    port map (
            O => \N__6943\,
            I => \N__6927\
        );

    \I__1593\ : InMux
    port map (
            O => \N__6942\,
            I => \N__6927\
        );

    \I__1592\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6924\
        );

    \I__1591\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6919\
        );

    \I__1590\ : InMux
    port map (
            O => \N__6939\,
            I => \N__6919\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__6932\,
            I => \N__6916\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__6927\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__6924\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__6919\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__6916\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__6907\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__1583\ : InMux
    port map (
            O => \N__6904\,
            I => \N__6901\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__6901\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__1581\ : InMux
    port map (
            O => \N__6898\,
            I => \N__6894\
        );

    \I__1580\ : InMux
    port map (
            O => \N__6897\,
            I => \N__6891\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__6894\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__6891\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1577\ : ClkMux
    port map (
            O => \N__6886\,
            I => \N__6853\
        );

    \I__1576\ : ClkMux
    port map (
            O => \N__6885\,
            I => \N__6853\
        );

    \I__1575\ : ClkMux
    port map (
            O => \N__6884\,
            I => \N__6853\
        );

    \I__1574\ : ClkMux
    port map (
            O => \N__6883\,
            I => \N__6853\
        );

    \I__1573\ : ClkMux
    port map (
            O => \N__6882\,
            I => \N__6853\
        );

    \I__1572\ : ClkMux
    port map (
            O => \N__6881\,
            I => \N__6853\
        );

    \I__1571\ : ClkMux
    port map (
            O => \N__6880\,
            I => \N__6853\
        );

    \I__1570\ : ClkMux
    port map (
            O => \N__6879\,
            I => \N__6853\
        );

    \I__1569\ : ClkMux
    port map (
            O => \N__6878\,
            I => \N__6853\
        );

    \I__1568\ : ClkMux
    port map (
            O => \N__6877\,
            I => \N__6853\
        );

    \I__1567\ : ClkMux
    port map (
            O => \N__6876\,
            I => \N__6853\
        );

    \I__1566\ : GlobalMux
    port map (
            O => \N__6853\,
            I => \N__6850\
        );

    \I__1565\ : gio2CtrlBuf
    port map (
            O => \N__6850\,
            I => \CLK6_c_g\
        );

    \I__1564\ : InMux
    port map (
            O => \N__6847\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__1563\ : InMux
    port map (
            O => \N__6844\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__1562\ : InMux
    port map (
            O => \N__6841\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__1561\ : InMux
    port map (
            O => \N__6838\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__1560\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6831\
        );

    \I__1559\ : InMux
    port map (
            O => \N__6834\,
            I => \N__6828\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__6831\,
            I => \N__6825\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__6828\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__1556\ : Odrv4
    port map (
            O => \N__6825\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__6820\,
            I => \U409_CIA.CLK_CIA6_3_cascade_\
        );

    \I__1554\ : CascadeMux
    port map (
            O => \N__6817\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_\
        );

    \I__1553\ : InMux
    port map (
            O => \N__6814\,
            I => \N__6811\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__6811\,
            I => \N__6807\
        );

    \I__1551\ : InMux
    port map (
            O => \N__6810\,
            I => \N__6804\
        );

    \I__1550\ : Span4Mux_v
    port map (
            O => \N__6807\,
            I => \N__6800\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__6804\,
            I => \N__6797\
        );

    \I__1548\ : InMux
    port map (
            O => \N__6803\,
            I => \N__6794\
        );

    \I__1547\ : Span4Mux_h
    port map (
            O => \N__6800\,
            I => \N__6791\
        );

    \I__1546\ : Span12Mux_h
    port map (
            O => \N__6797\,
            I => \N__6788\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__6794\,
            I => \N__6785\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__6791\,
            I => \CIA_SPACE\
        );

    \I__1543\ : Odrv12
    port map (
            O => \N__6788\,
            I => \CIA_SPACE\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__6785\,
            I => \CIA_SPACE\
        );

    \I__1541\ : CascadeMux
    port map (
            O => \N__6778\,
            I => \U409_CIA.VMA_RNOZ0Z_0_cascade_\
        );

    \I__1540\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6771\
        );

    \I__1539\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6768\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__6771\,
            I => \N__6765\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__6768\,
            I => \N__6761\
        );

    \I__1536\ : Span4Mux_v
    port map (
            O => \N__6765\,
            I => \N__6758\
        );

    \I__1535\ : InMux
    port map (
            O => \N__6764\,
            I => \N__6755\
        );

    \I__1534\ : Odrv12
    port map (
            O => \N__6761\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__6758\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__6755\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1531\ : InMux
    port map (
            O => \N__6748\,
            I => \N__6744\
        );

    \I__1530\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6741\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__6744\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__6741\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__1527\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6733\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__6733\,
            I => \N__6730\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__6730\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__1524\ : InMux
    port map (
            O => \N__6727\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__1523\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6720\
        );

    \I__1522\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6717\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__6720\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__6717\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__6712\,
            I => \N__6709\
        );

    \I__1518\ : InMux
    port map (
            O => \N__6709\,
            I => \N__6706\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__6706\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__1516\ : InMux
    port map (
            O => \N__6703\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__1515\ : InMux
    port map (
            O => \N__6700\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__6697\,
            I => \N__6694\
        );

    \I__1513\ : InMux
    port map (
            O => \N__6694\,
            I => \N__6690\
        );

    \I__1512\ : InMux
    port map (
            O => \N__6693\,
            I => \N__6687\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__6690\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__6687\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__1509\ : InMux
    port map (
            O => \N__6682\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__6679\,
            I => \N__6675\
        );

    \I__1507\ : InMux
    port map (
            O => \N__6678\,
            I => \N__6672\
        );

    \I__1506\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6669\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__6672\,
            I => \N__6666\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__6669\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__1503\ : Odrv4
    port map (
            O => \N__6666\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__1502\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6658\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__6658\,
            I => \N__6655\
        );

    \I__1500\ : Odrv4
    port map (
            O => \N__6655\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__1499\ : InMux
    port map (
            O => \N__6652\,
            I => \bfn_14_10_0_\
        );

    \I__1498\ : InMux
    port map (
            O => \N__6649\,
            I => \N__6646\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__6646\,
            I => \N__6642\
        );

    \I__1496\ : InMux
    port map (
            O => \N__6645\,
            I => \N__6639\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__6642\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__6639\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__1493\ : InMux
    port map (
            O => \N__6634\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__1492\ : InMux
    port map (
            O => \N__6631\,
            I => \N__6627\
        );

    \I__1491\ : InMux
    port map (
            O => \N__6630\,
            I => \N__6624\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__6627\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__6624\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__1488\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6616\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__6616\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__1486\ : InMux
    port map (
            O => \N__6613\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__1485\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6607\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__6607\,
            I => \N__6603\
        );

    \I__1483\ : InMux
    port map (
            O => \N__6606\,
            I => \N__6600\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__6603\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__6600\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__1480\ : InMux
    port map (
            O => \N__6595\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__1479\ : CascadeMux
    port map (
            O => \N__6592\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__1478\ : InMux
    port map (
            O => \N__6589\,
            I => \N__6586\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__6586\,
            I => \U409_TICK.TICK503_8\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__6583\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__1475\ : InMux
    port map (
            O => \N__6580\,
            I => \N__6574\
        );

    \I__1474\ : InMux
    port map (
            O => \N__6579\,
            I => \N__6569\
        );

    \I__1473\ : InMux
    port map (
            O => \N__6578\,
            I => \N__6569\
        );

    \I__1472\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6566\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__6574\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__6569\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__6566\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__6559\,
            I => \N__6554\
        );

    \I__1467\ : InMux
    port map (
            O => \N__6558\,
            I => \N__6551\
        );

    \I__1466\ : InMux
    port map (
            O => \N__6557\,
            I => \N__6548\
        );

    \I__1465\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6545\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__6551\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__6548\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__6545\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1461\ : InMux
    port map (
            O => \N__6538\,
            I => \N__6534\
        );

    \I__1460\ : InMux
    port map (
            O => \N__6537\,
            I => \N__6531\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__6534\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__6531\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__1457\ : InMux
    port map (
            O => \N__6526\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__1456\ : InMux
    port map (
            O => \N__6523\,
            I => \N__6519\
        );

    \I__1455\ : InMux
    port map (
            O => \N__6522\,
            I => \N__6516\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__6519\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__6516\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__1452\ : InMux
    port map (
            O => \N__6511\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__1451\ : InMux
    port map (
            O => \N__6508\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__1450\ : InMux
    port map (
            O => \N__6505\,
            I => \N__6502\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__6502\,
            I => \N__6496\
        );

    \I__1448\ : InMux
    port map (
            O => \N__6501\,
            I => \N__6491\
        );

    \I__1447\ : InMux
    port map (
            O => \N__6500\,
            I => \N__6491\
        );

    \I__1446\ : InMux
    port map (
            O => \N__6499\,
            I => \N__6488\
        );

    \I__1445\ : Span4Mux_h
    port map (
            O => \N__6496\,
            I => \N__6485\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__6491\,
            I => \N__6482\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__6488\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__6485\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1441\ : Odrv4
    port map (
            O => \N__6482\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1440\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6472\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__6472\,
            I => \N__6467\
        );

    \I__1438\ : InMux
    port map (
            O => \N__6471\,
            I => \N__6462\
        );

    \I__1437\ : InMux
    port map (
            O => \N__6470\,
            I => \N__6462\
        );

    \I__1436\ : Span4Mux_h
    port map (
            O => \N__6467\,
            I => \N__6459\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__6462\,
            I => \N__6456\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__6459\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__1433\ : Odrv12
    port map (
            O => \N__6456\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__1432\ : SRMux
    port map (
            O => \N__6451\,
            I => \N__6447\
        );

    \I__1431\ : SRMux
    port map (
            O => \N__6450\,
            I => \N__6443\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6447\,
            I => \N__6438\
        );

    \I__1429\ : SRMux
    port map (
            O => \N__6446\,
            I => \N__6435\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__6443\,
            I => \N__6431\
        );

    \I__1427\ : SRMux
    port map (
            O => \N__6442\,
            I => \N__6428\
        );

    \I__1426\ : SRMux
    port map (
            O => \N__6441\,
            I => \N__6425\
        );

    \I__1425\ : Span4Mux_v
    port map (
            O => \N__6438\,
            I => \N__6420\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__6435\,
            I => \N__6420\
        );

    \I__1423\ : SRMux
    port map (
            O => \N__6434\,
            I => \N__6417\
        );

    \I__1422\ : Span4Mux_h
    port map (
            O => \N__6431\,
            I => \N__6412\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__6428\,
            I => \N__6412\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__6425\,
            I => \N__6409\
        );

    \I__1419\ : Span4Mux_v
    port map (
            O => \N__6420\,
            I => \N__6403\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__6417\,
            I => \N__6403\
        );

    \I__1417\ : Span4Mux_v
    port map (
            O => \N__6412\,
            I => \N__6400\
        );

    \I__1416\ : Span4Mux_h
    port map (
            O => \N__6409\,
            I => \N__6397\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6408\,
            I => \N__6394\
        );

    \I__1414\ : Span4Mux_v
    port map (
            O => \N__6403\,
            I => \N__6391\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__6400\,
            I => \RESETn_c_i\
        );

    \I__1412\ : Odrv4
    port map (
            O => \N__6397\,
            I => \RESETn_c_i\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6394\,
            I => \RESETn_c_i\
        );

    \I__1410\ : Odrv4
    port map (
            O => \N__6391\,
            I => \RESETn_c_i\
        );

    \I__1409\ : IoInMux
    port map (
            O => \N__6382\,
            I => \N__6379\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__6379\,
            I => \N__6375\
        );

    \I__1407\ : IoInMux
    port map (
            O => \N__6378\,
            I => \N__6372\
        );

    \I__1406\ : IoSpan4Mux
    port map (
            O => \N__6375\,
            I => \N__6367\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__6372\,
            I => \N__6367\
        );

    \I__1404\ : IoSpan4Mux
    port map (
            O => \N__6367\,
            I => \N__6364\
        );

    \I__1403\ : Span4Mux_s2_v
    port map (
            O => \N__6364\,
            I => \N__6361\
        );

    \I__1402\ : Sp12to4
    port map (
            O => \N__6361\,
            I => \N__6357\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6360\,
            I => \N__6354\
        );

    \I__1400\ : Span12Mux_s10_v
    port map (
            O => \N__6357\,
            I => \N__6348\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__6354\,
            I => \N__6348\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__6353\,
            I => \N__6345\
        );

    \I__1397\ : Span12Mux_h
    port map (
            O => \N__6348\,
            I => \N__6342\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6345\,
            I => \N__6339\
        );

    \I__1395\ : Odrv12
    port map (
            O => \N__6342\,
            I => \TACK_EN\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6339\,
            I => \TACK_EN\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6334\,
            I => \N__6330\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6333\,
            I => \N__6327\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6330\,
            I => \N__6323\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6327\,
            I => \N__6320\
        );

    \I__1389\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6317\
        );

    \I__1388\ : Span4Mux_v
    port map (
            O => \N__6323\,
            I => \N__6314\
        );

    \I__1387\ : Span4Mux_v
    port map (
            O => \N__6320\,
            I => \N__6311\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__6317\,
            I => \N__6308\
        );

    \I__1385\ : Sp12to4
    port map (
            O => \N__6314\,
            I => \N__6305\
        );

    \I__1384\ : Span4Mux_h
    port map (
            O => \N__6311\,
            I => \N__6300\
        );

    \I__1383\ : Span4Mux_v
    port map (
            O => \N__6308\,
            I => \N__6300\
        );

    \I__1382\ : Odrv12
    port map (
            O => \N__6305\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__6300\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__1380\ : IoInMux
    port map (
            O => \N__6295\,
            I => \N__6292\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6292\,
            I => \N__6289\
        );

    \I__1378\ : Span12Mux_s1_v
    port map (
            O => \N__6289\,
            I => \N__6286\
        );

    \I__1377\ : Span12Mux_h
    port map (
            O => \N__6286\,
            I => \N__6283\
        );

    \I__1376\ : Odrv12
    port map (
            O => \N__6283\,
            I => \TCIn_1_i\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6280\,
            I => \N__6277\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__6277\,
            I => \N__6274\
        );

    \I__1373\ : Span12Mux_v
    port map (
            O => \N__6274\,
            I => \N__6271\
        );

    \I__1372\ : Span12Mux_h
    port map (
            O => \N__6271\,
            I => \N__6268\
        );

    \I__1371\ : Odrv12
    port map (
            O => \N__6268\,
            I => \A_c_13\
        );

    \I__1370\ : IoInMux
    port map (
            O => \N__6265\,
            I => \N__6262\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__6262\,
            I => \N__6259\
        );

    \I__1368\ : Span4Mux_s2_h
    port map (
            O => \N__6259\,
            I => \N__6256\
        );

    \I__1367\ : Span4Mux_h
    port map (
            O => \N__6256\,
            I => \N__6253\
        );

    \I__1366\ : Sp12to4
    port map (
            O => \N__6253\,
            I => \N__6250\
        );

    \I__1365\ : Span12Mux_s9_v
    port map (
            O => \N__6250\,
            I => \N__6247\
        );

    \I__1364\ : Odrv12
    port map (
            O => \N__6247\,
            I => \U409_ADDRESS_DECODE_un1_CIACS1n_i\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6244\,
            I => \N__6239\
        );

    \I__1362\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6236\
        );

    \I__1361\ : InMux
    port map (
            O => \N__6242\,
            I => \N__6233\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__6239\,
            I => \N__6227\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__6236\,
            I => \N__6227\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__6233\,
            I => \N__6222\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__6232\,
            I => \N__6219\
        );

    \I__1356\ : Span4Mux_v
    port map (
            O => \N__6227\,
            I => \N__6216\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6226\,
            I => \N__6213\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__6225\,
            I => \N__6209\
        );

    \I__1353\ : Span4Mux_v
    port map (
            O => \N__6222\,
            I => \N__6204\
        );

    \I__1352\ : InMux
    port map (
            O => \N__6219\,
            I => \N__6201\
        );

    \I__1351\ : Span4Mux_h
    port map (
            O => \N__6216\,
            I => \N__6196\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6213\,
            I => \N__6196\
        );

    \I__1349\ : InMux
    port map (
            O => \N__6212\,
            I => \N__6189\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6209\,
            I => \N__6189\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6208\,
            I => \N__6189\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6207\,
            I => \N__6182\
        );

    \I__1345\ : Span4Mux_h
    port map (
            O => \N__6204\,
            I => \N__6179\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__6201\,
            I => \N__6176\
        );

    \I__1343\ : Span4Mux_v
    port map (
            O => \N__6196\,
            I => \N__6171\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6189\,
            I => \N__6171\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6188\,
            I => \N__6168\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6187\,
            I => \N__6165\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6186\,
            I => \N__6162\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6159\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6182\,
            I => \N__6156\
        );

    \I__1336\ : Span4Mux_h
    port map (
            O => \N__6179\,
            I => \N__6151\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__6176\,
            I => \N__6151\
        );

    \I__1334\ : Span4Mux_h
    port map (
            O => \N__6171\,
            I => \N__6142\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__6168\,
            I => \N__6142\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6165\,
            I => \N__6142\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__6162\,
            I => \N__6142\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__6159\,
            I => \N__6139\
        );

    \I__1329\ : Span12Mux_h
    port map (
            O => \N__6156\,
            I => \N__6134\
        );

    \I__1328\ : Sp12to4
    port map (
            O => \N__6151\,
            I => \N__6134\
        );

    \I__1327\ : Span4Mux_v
    port map (
            O => \N__6142\,
            I => \N__6131\
        );

    \I__1326\ : Span4Mux_v
    port map (
            O => \N__6139\,
            I => \N__6128\
        );

    \I__1325\ : Span12Mux_v
    port map (
            O => \N__6134\,
            I => \N__6121\
        );

    \I__1324\ : Sp12to4
    port map (
            O => \N__6131\,
            I => \N__6121\
        );

    \I__1323\ : Sp12to4
    port map (
            O => \N__6128\,
            I => \N__6121\
        );

    \I__1322\ : Span12Mux_h
    port map (
            O => \N__6121\,
            I => \N__6118\
        );

    \I__1321\ : Odrv12
    port map (
            O => \N__6118\,
            I => \RESETn_c\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6115\,
            I => \N__6112\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6112\,
            I => \CIA_ENABLE\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6109\,
            I => \N__6106\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6106\,
            I => \N__6103\
        );

    \I__1316\ : Span4Mux_v
    port map (
            O => \N__6103\,
            I => \N__6100\
        );

    \I__1315\ : Sp12to4
    port map (
            O => \N__6100\,
            I => \N__6097\
        );

    \I__1314\ : Span12Mux_h
    port map (
            O => \N__6097\,
            I => \N__6094\
        );

    \I__1313\ : Odrv12
    port map (
            O => \N__6094\,
            I => \A_c_12\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__6091\,
            I => \CIA_ENABLE_cascade_\
        );

    \I__1311\ : IoInMux
    port map (
            O => \N__6088\,
            I => \N__6085\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__6085\,
            I => \N__6082\
        );

    \I__1309\ : IoSpan4Mux
    port map (
            O => \N__6082\,
            I => \N__6079\
        );

    \I__1308\ : Sp12to4
    port map (
            O => \N__6079\,
            I => \N__6076\
        );

    \I__1307\ : Span12Mux_s7_v
    port map (
            O => \N__6076\,
            I => \N__6073\
        );

    \I__1306\ : Span12Mux_h
    port map (
            O => \N__6073\,
            I => \N__6070\
        );

    \I__1305\ : Odrv12
    port map (
            O => \N__6070\,
            I => \U409_ADDRESS_DECODE_un1_CIACS0n_i\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__6067\,
            I => \U409_TICK.TICK503_11_cascade_\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6064\,
            I => \N__6060\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6063\,
            I => \N__6057\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__6060\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6057\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6048\
        );

    \I__1298\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6045\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6048\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__6045\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__6040\,
            I => \N__6035\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__6039\,
            I => \N__6032\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6029\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6026\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6032\,
            I => \N__6023\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__6029\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6026\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6023\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6016\,
            I => \N__6012\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6015\,
            I => \N__6009\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__6012\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__6009\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6004\,
            I => \N__6000\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6003\,
            I => \N__5997\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6000\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__5997\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5992\,
            I => \N__5989\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5989\,
            I => \U409_TICK.TICK603_8\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__5986\,
            I => \U409_TICK.TICK603_11_cascade_\
        );

    \I__1276\ : InMux
    port map (
            O => \N__5983\,
            I => \N__5979\
        );

    \I__1275\ : InMux
    port map (
            O => \N__5982\,
            I => \N__5976\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__5979\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__5976\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__5971\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__1271\ : InMux
    port map (
            O => \N__5968\,
            I => \N__5965\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__5965\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5962\,
            I => \N__5958\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5961\,
            I => \N__5955\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__5958\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__5955\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5950\,
            I => \N__5946\
        );

    \I__1264\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5943\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5946\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__5943\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__5938\,
            I => \N__5935\
        );

    \I__1260\ : InMux
    port map (
            O => \N__5935\,
            I => \N__5931\
        );

    \I__1259\ : InMux
    port map (
            O => \N__5934\,
            I => \N__5928\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__5931\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5928\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__5923\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5920\,
            I => \N__5917\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__5917\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5914\,
            I => \N__5910\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5913\,
            I => \N__5907\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__5910\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__5907\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5898\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5901\,
            I => \N__5895\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__5898\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__5895\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5890\,
            I => \N__5886\
        );

    \I__1244\ : InMux
    port map (
            O => \N__5889\,
            I => \N__5883\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__5886\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5883\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__5878\,
            I => \N__5875\
        );

    \I__1240\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5871\
        );

    \I__1239\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5868\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__5871\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__5868\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__5863\,
            I => \U409_TICK.TICK603_10_cascade_\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5857\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5857\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__1233\ : InMux
    port map (
            O => \N__5854\,
            I => \N__5850\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5853\,
            I => \N__5847\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__5850\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5847\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5833\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5828\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5828\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5823\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5823\
        );

    \I__1224\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5818\
        );

    \I__1223\ : InMux
    port map (
            O => \N__5836\,
            I => \N__5818\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__5833\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5828\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__5823\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5818\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__5809\,
            I => \N__5805\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__5808\,
            I => \N__5802\
        );

    \I__1216\ : InMux
    port map (
            O => \N__5805\,
            I => \N__5794\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5789\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5789\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5784\
        );

    \I__1212\ : InMux
    port map (
            O => \N__5799\,
            I => \N__5784\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5779\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5779\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__5794\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__5789\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__5784\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__5779\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5770\,
            I => \N__5762\
        );

    \I__1204\ : CascadeMux
    port map (
            O => \N__5769\,
            I => \N__5759\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__5768\,
            I => \N__5755\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5767\,
            I => \N__5750\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5766\,
            I => \N__5750\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5765\,
            I => \N__5747\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5762\,
            I => \N__5744\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5759\,
            I => \N__5739\
        );

    \I__1197\ : InMux
    port map (
            O => \N__5758\,
            I => \N__5739\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5755\,
            I => \N__5736\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5750\,
            I => \N__5733\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5747\,
            I => \N__5730\
        );

    \I__1193\ : Odrv12
    port map (
            O => \N__5744\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5739\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__5736\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1190\ : Odrv4
    port map (
            O => \N__5733\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1189\ : Odrv4
    port map (
            O => \N__5730\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5716\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5716\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5713\,
            I => \N__5709\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5712\,
            I => \N__5706\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__5709\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5706\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__5701\,
            I => \N__5698\
        );

    \I__1181\ : InMux
    port map (
            O => \N__5698\,
            I => \N__5693\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5697\,
            I => \N__5690\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__5696\,
            I => \N__5685\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5693\,
            I => \N__5680\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__5690\,
            I => \N__5680\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5673\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5688\,
            I => \N__5673\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5685\,
            I => \N__5673\
        );

    \I__1173\ : Span4Mux_h
    port map (
            O => \N__5680\,
            I => \N__5670\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__5673\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1171\ : Odrv4
    port map (
            O => \N__5670\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__5665\,
            I => \U409_TRANSFER_ACK.N_9_cascade_\
        );

    \I__1169\ : IoInMux
    port map (
            O => \N__5662\,
            I => \N__5659\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__5659\,
            I => \N__5656\
        );

    \I__1167\ : Span4Mux_s3_v
    port map (
            O => \N__5656\,
            I => \N__5653\
        );

    \I__1166\ : Span4Mux_v
    port map (
            O => \N__5653\,
            I => \N__5650\
        );

    \I__1165\ : Span4Mux_v
    port map (
            O => \N__5650\,
            I => \N__5647\
        );

    \I__1164\ : Span4Mux_h
    port map (
            O => \N__5647\,
            I => \N__5643\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5646\,
            I => \N__5640\
        );

    \I__1162\ : Odrv4
    port map (
            O => \N__5643\,
            I => \TICK60_c\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5640\,
            I => \TICK60_c\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5635\,
            I => \N__5632\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5632\,
            I => \U409_TRANSFER_ACK.N_4\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5629\,
            I => \N__5626\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5626\,
            I => \N__5622\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__5625\,
            I => \N__5618\
        );

    \I__1155\ : Span4Mux_h
    port map (
            O => \N__5622\,
            I => \N__5614\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5621\,
            I => \N__5609\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5609\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5606\
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__5614\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5609\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5606\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5599\,
            I => \N__5592\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5598\,
            I => \N__5592\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5589\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5592\,
            I => \N__5584\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__5589\,
            I => \N__5584\
        );

    \I__1143\ : Odrv4
    port map (
            O => \N__5584\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__5581\,
            I => \U409_TRANSFER_ACK.N_4_cascade_\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5578\,
            I => \N__5572\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5577\,
            I => \N__5569\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5576\,
            I => \N__5564\
        );

    \I__1138\ : InMux
    port map (
            O => \N__5575\,
            I => \N__5564\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5572\,
            I => \N__5561\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__5569\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5564\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__5561\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5554\,
            I => \N__5551\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__5551\,
            I => \U409_TRANSFER_ACK.N_5\
        );

    \I__1131\ : IoInMux
    port map (
            O => \N__5548\,
            I => \N__5543\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__5547\,
            I => \N__5538\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__5546\,
            I => \N__5535\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5543\,
            I => \N__5531\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__5542\,
            I => \N__5528\
        );

    \I__1126\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5524\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5538\,
            I => \N__5521\
        );

    \I__1124\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5518\
        );

    \I__1123\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5515\
        );

    \I__1122\ : IoSpan4Mux
    port map (
            O => \N__5531\,
            I => \N__5512\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5528\,
            I => \N__5507\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5507\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__5524\,
            I => \N__5500\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5521\,
            I => \N__5500\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__5518\,
            I => \N__5500\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5515\,
            I => \N__5497\
        );

    \I__1115\ : Span4Mux_s0_v
    port map (
            O => \N__5512\,
            I => \N__5493\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__5507\,
            I => \N__5490\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__5500\,
            I => \N__5487\
        );

    \I__1112\ : Span4Mux_v
    port map (
            O => \N__5497\,
            I => \N__5484\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5496\,
            I => \N__5481\
        );

    \I__1110\ : Sp12to4
    port map (
            O => \N__5493\,
            I => \N__5478\
        );

    \I__1109\ : Span4Mux_h
    port map (
            O => \N__5490\,
            I => \N__5475\
        );

    \I__1108\ : Sp12to4
    port map (
            O => \N__5487\,
            I => \N__5470\
        );

    \I__1107\ : Sp12to4
    port map (
            O => \N__5484\,
            I => \N__5470\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__5481\,
            I => \N__5467\
        );

    \I__1105\ : Span12Mux_v
    port map (
            O => \N__5478\,
            I => \N__5458\
        );

    \I__1104\ : Sp12to4
    port map (
            O => \N__5475\,
            I => \N__5458\
        );

    \I__1103\ : Span12Mux_h
    port map (
            O => \N__5470\,
            I => \N__5458\
        );

    \I__1102\ : Span12Mux_h
    port map (
            O => \N__5467\,
            I => \N__5458\
        );

    \I__1101\ : Span12Mux_v
    port map (
            O => \N__5458\,
            I => \N__5455\
        );

    \I__1100\ : Odrv12
    port map (
            O => \N__5455\,
            I => \CLK40_IN_c\
        );

    \I__1099\ : InMux
    port map (
            O => \N__5452\,
            I => \N__5449\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5449\,
            I => \U409_TRANSFER_ACK.m8_ns_1\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5443\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5443\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__1095\ : InMux
    port map (
            O => \N__5440\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5437\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5434\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__1092\ : InMux
    port map (
            O => \N__5431\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5428\,
            I => \N__5424\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5427\,
            I => \N__5421\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5424\,
            I => \N__5416\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5421\,
            I => \N__5416\
        );

    \I__1087\ : Span4Mux_v
    port map (
            O => \N__5416\,
            I => \N__5413\
        );

    \I__1086\ : Odrv4
    port map (
            O => \N__5413\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn\
        );

    \I__1085\ : InMux
    port map (
            O => \N__5410\,
            I => \N__5406\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5409\,
            I => \N__5403\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__5406\,
            I => \N__5397\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__5403\,
            I => \N__5397\
        );

    \I__1081\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5394\
        );

    \I__1080\ : Odrv12
    port map (
            O => \N__5397\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__5394\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__1078\ : IoInMux
    port map (
            O => \N__5389\,
            I => \N__5386\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5386\,
            I => \N__5383\
        );

    \I__1076\ : IoSpan4Mux
    port map (
            O => \N__5383\,
            I => \N__5380\
        );

    \I__1075\ : Span4Mux_s2_v
    port map (
            O => \N__5380\,
            I => \N__5377\
        );

    \I__1074\ : Sp12to4
    port map (
            O => \N__5377\,
            I => \N__5374\
        );

    \I__1073\ : Span12Mux_s10_v
    port map (
            O => \N__5374\,
            I => \N__5371\
        );

    \I__1072\ : Odrv12
    port map (
            O => \N__5371\,
            I => \BUFENn_c\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__5368\,
            I => \U409_TRANSFER_ACK.i6_mux_0_cascade_\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5365\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__1069\ : InMux
    port map (
            O => \N__5362\,
            I => \N__5358\
        );

    \I__1068\ : InMux
    port map (
            O => \N__5361\,
            I => \N__5355\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__5358\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5355\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5350\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__1064\ : InMux
    port map (
            O => \N__5347\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5344\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5338\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5338\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5335\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__1059\ : InMux
    port map (
            O => \N__5332\,
            I => \bfn_12_10_0_\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5329\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5326\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5323\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5320\,
            I => \N__5314\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5319\,
            I => \N__5309\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5318\,
            I => \N__5309\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5317\,
            I => \N__5306\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__5314\,
            I => \N__5296\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__5309\,
            I => \N__5296\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__5306\,
            I => \N__5296\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5305\,
            I => \N__5293\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5304\,
            I => \N__5290\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5287\
        );

    \I__1045\ : Span4Mux_v
    port map (
            O => \N__5296\,
            I => \N__5282\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__5293\,
            I => \N__5282\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5290\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5287\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__5282\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1040\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5270\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__5274\,
            I => \N__5265\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5261\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__5270\,
            I => \N__5258\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5255\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5252\
        );

    \I__1034\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5246\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5246\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5261\,
            I => \N__5241\
        );

    \I__1031\ : Span4Mux_v
    port map (
            O => \N__5258\,
            I => \N__5241\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5255\,
            I => \N__5236\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5252\,
            I => \N__5236\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5251\,
            I => \N__5233\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5246\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1026\ : Odrv4
    port map (
            O => \N__5241\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1025\ : Odrv4
    port map (
            O => \N__5236\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__5233\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__5224\,
            I => \N__5220\
        );

    \I__1022\ : CascadeMux
    port map (
            O => \N__5223\,
            I => \N__5216\
        );

    \I__1021\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5206\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5219\,
            I => \N__5206\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5216\,
            I => \N__5206\
        );

    \I__1018\ : InMux
    port map (
            O => \N__5215\,
            I => \N__5203\
        );

    \I__1017\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5198\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__5213\,
            I => \N__5195\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5206\,
            I => \N__5190\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5203\,
            I => \N__5190\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5185\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5185\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__5198\,
            I => \N__5182\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5195\,
            I => \N__5179\
        );

    \I__1009\ : Span4Mux_v
    port map (
            O => \N__5190\,
            I => \N__5176\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5185\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1007\ : Odrv4
    port map (
            O => \N__5182\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__5179\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__5176\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5167\,
            I => \N__5164\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5164\,
            I => \N__5157\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5163\,
            I => \N__5154\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5162\,
            I => \N__5151\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5145\
        );

    \I__999\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5145\
        );

    \I__998\ : Span4Mux_h
    port map (
            O => \N__5157\,
            I => \N__5142\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5154\,
            I => \N__5137\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5151\,
            I => \N__5137\
        );

    \I__995\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5134\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5145\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__5142\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__992\ : Odrv4
    port map (
            O => \N__5137\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5134\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__990\ : InMux
    port map (
            O => \N__5125\,
            I => \N__5122\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__5122\,
            I => \N__5119\
        );

    \I__988\ : Odrv4
    port map (
            O => \N__5119\,
            I => \U409_TRANSFER_ACK.N_36\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__5116\,
            I => \N__5113\
        );

    \I__986\ : InMux
    port map (
            O => \N__5113\,
            I => \N__5103\
        );

    \I__985\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5103\
        );

    \I__984\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5103\
        );

    \I__983\ : InMux
    port map (
            O => \N__5110\,
            I => \N__5100\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5103\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5100\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__980\ : InMux
    port map (
            O => \N__5095\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__979\ : InMux
    port map (
            O => \N__5092\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__5089\,
            I => \N__5083\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__5088\,
            I => \N__5080\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__5087\,
            I => \N__5077\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__5086\,
            I => \N__5074\
        );

    \I__974\ : InMux
    port map (
            O => \N__5083\,
            I => \N__5062\
        );

    \I__973\ : InMux
    port map (
            O => \N__5080\,
            I => \N__5062\
        );

    \I__972\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5062\
        );

    \I__971\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5062\
        );

    \I__970\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5062\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__5062\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__5059\,
            I => \N__5053\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__5058\,
            I => \N__5050\
        );

    \I__966\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5047\
        );

    \I__965\ : InMux
    port map (
            O => \N__5056\,
            I => \N__5044\
        );

    \I__964\ : InMux
    port map (
            O => \N__5053\,
            I => \N__5041\
        );

    \I__963\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5038\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5047\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__5044\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__5041\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__5038\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__958\ : InMux
    port map (
            O => \N__5029\,
            I => \N__5023\
        );

    \I__957\ : InMux
    port map (
            O => \N__5028\,
            I => \N__5020\
        );

    \I__956\ : InMux
    port map (
            O => \N__5027\,
            I => \N__5015\
        );

    \I__955\ : InMux
    port map (
            O => \N__5026\,
            I => \N__5015\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5023\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5020\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__5015\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__951\ : InMux
    port map (
            O => \N__5008\,
            I => \N__5002\
        );

    \I__950\ : InMux
    port map (
            O => \N__5007\,
            I => \N__5002\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5002\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__948\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4988\
        );

    \I__947\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4988\
        );

    \I__946\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4985\
        );

    \I__945\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4982\
        );

    \I__944\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4979\
        );

    \I__943\ : InMux
    port map (
            O => \N__4994\,
            I => \N__4974\
        );

    \I__942\ : InMux
    port map (
            O => \N__4993\,
            I => \N__4974\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__4988\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4985\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4982\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4979\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__4974\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__936\ : InMux
    port map (
            O => \N__4963\,
            I => \N__4958\
        );

    \I__935\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4955\
        );

    \I__934\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4952\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4958\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4955\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4952\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__930\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4937\
        );

    \I__929\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4937\
        );

    \I__928\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4934\
        );

    \I__927\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4931\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4937\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4934\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4931\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__923\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4919\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__4923\,
            I => \N__4916\
        );

    \I__921\ : InMux
    port map (
            O => \N__4922\,
            I => \N__4913\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4919\,
            I => \N__4910\
        );

    \I__919\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4907\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4913\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__917\ : Odrv4
    port map (
            O => \N__4910\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4907\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__915\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4892\
        );

    \I__914\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4892\
        );

    \I__913\ : InMux
    port map (
            O => \N__4898\,
            I => \N__4887\
        );

    \I__912\ : InMux
    port map (
            O => \N__4897\,
            I => \N__4884\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4892\,
            I => \N__4881\
        );

    \I__910\ : InMux
    port map (
            O => \N__4891\,
            I => \N__4876\
        );

    \I__909\ : InMux
    port map (
            O => \N__4890\,
            I => \N__4876\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4887\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4884\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__906\ : Odrv4
    port map (
            O => \N__4881\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4876\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__4867\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\
        );

    \I__903\ : InMux
    port map (
            O => \N__4864\,
            I => \N__4857\
        );

    \I__902\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4852\
        );

    \I__901\ : InMux
    port map (
            O => \N__4862\,
            I => \N__4852\
        );

    \I__900\ : InMux
    port map (
            O => \N__4861\,
            I => \N__4847\
        );

    \I__899\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4847\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4857\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4852\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4847\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__895\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4837\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4837\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5\
        );

    \I__893\ : InMux
    port map (
            O => \N__4834\,
            I => \N__4831\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4831\,
            I => \N__4826\
        );

    \I__891\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4823\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__4829\,
            I => \N__4820\
        );

    \I__889\ : Span4Mux_h
    port map (
            O => \N__4826\,
            I => \N__4815\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4823\,
            I => \N__4815\
        );

    \I__887\ : InMux
    port map (
            O => \N__4820\,
            I => \N__4812\
        );

    \I__886\ : Span4Mux_h
    port map (
            O => \N__4815\,
            I => \N__4806\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4812\,
            I => \N__4806\
        );

    \I__884\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4803\
        );

    \I__883\ : Span4Mux_v
    port map (
            O => \N__4806\,
            I => \N__4798\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4803\,
            I => \N__4798\
        );

    \I__881\ : Span4Mux_h
    port map (
            O => \N__4798\,
            I => \N__4795\
        );

    \I__880\ : Odrv4
    port map (
            O => \N__4795\,
            I => \U409_ADDRESS_DECODE_ROMEN_1\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__4792\,
            I => \N__4789\
        );

    \I__878\ : InMux
    port map (
            O => \N__4789\,
            I => \N__4785\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__4788\,
            I => \N__4782\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4785\,
            I => \N__4779\
        );

    \I__875\ : InMux
    port map (
            O => \N__4782\,
            I => \N__4776\
        );

    \I__874\ : Span4Mux_h
    port map (
            O => \N__4779\,
            I => \N__4771\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4776\,
            I => \N__4771\
        );

    \I__872\ : Span4Mux_h
    port map (
            O => \N__4771\,
            I => \N__4768\
        );

    \I__871\ : Odrv4
    port map (
            O => \N__4768\,
            I => \U409_TRANSFER_ACK.N_23\
        );

    \I__870\ : InMux
    port map (
            O => \N__4765\,
            I => \N__4762\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4762\,
            I => \N__4759\
        );

    \I__868\ : Sp12to4
    port map (
            O => \N__4759\,
            I => \N__4756\
        );

    \I__867\ : Span12Mux_s9_v
    port map (
            O => \N__4756\,
            I => \N__4753\
        );

    \I__866\ : Span12Mux_h
    port map (
            O => \N__4753\,
            I => \N__4750\
        );

    \I__865\ : Odrv12
    port map (
            O => \N__4750\,
            I => \TACKn_in\
        );

    \I__864\ : SRMux
    port map (
            O => \N__4747\,
            I => \N__4743\
        );

    \I__863\ : SRMux
    port map (
            O => \N__4746\,
            I => \N__4740\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4743\,
            I => \N__4736\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4740\,
            I => \N__4733\
        );

    \I__860\ : SRMux
    port map (
            O => \N__4739\,
            I => \N__4730\
        );

    \I__859\ : Span4Mux_h
    port map (
            O => \N__4736\,
            I => \N__4727\
        );

    \I__858\ : Span4Mux_h
    port map (
            O => \N__4733\,
            I => \N__4722\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4730\,
            I => \N__4722\
        );

    \I__856\ : Span4Mux_v
    port map (
            O => \N__4727\,
            I => \N__4716\
        );

    \I__855\ : Span4Mux_v
    port map (
            O => \N__4722\,
            I => \N__4716\
        );

    \I__854\ : SRMux
    port map (
            O => \N__4721\,
            I => \N__4713\
        );

    \I__853\ : Span4Mux_v
    port map (
            O => \N__4716\,
            I => \N__4708\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__4713\,
            I => \N__4708\
        );

    \I__851\ : Span4Mux_v
    port map (
            O => \N__4708\,
            I => \N__4705\
        );

    \I__850\ : Span4Mux_v
    port map (
            O => \N__4705\,
            I => \N__4702\
        );

    \I__849\ : Odrv4
    port map (
            O => \N__4702\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__848\ : IoInMux
    port map (
            O => \N__4699\,
            I => \N__4696\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4696\,
            I => \N__4693\
        );

    \I__846\ : Span4Mux_s2_v
    port map (
            O => \N__4693\,
            I => \N__4690\
        );

    \I__845\ : Span4Mux_v
    port map (
            O => \N__4690\,
            I => \N__4687\
        );

    \I__844\ : Odrv4
    port map (
            O => \N__4687\,
            I => \CONSTANT_ONE_NET\
        );

    \I__843\ : InMux
    port map (
            O => \N__4684\,
            I => \N__4681\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4681\,
            I => \N__4678\
        );

    \I__841\ : Odrv4
    port map (
            O => \N__4678\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_1_0\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__4675\,
            I => \N__4672\
        );

    \I__839\ : InMux
    port map (
            O => \N__4672\,
            I => \N__4669\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4669\,
            I => \N__4665\
        );

    \I__837\ : InMux
    port map (
            O => \N__4668\,
            I => \N__4662\
        );

    \I__836\ : Span4Mux_v
    port map (
            O => \N__4665\,
            I => \N__4657\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4662\,
            I => \N__4657\
        );

    \I__834\ : Odrv4
    port map (
            O => \N__4657\,
            I => \U409_TRANSFER_ACK.N_35_1\
        );

    \I__833\ : InMux
    port map (
            O => \N__4654\,
            I => \N__4651\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4651\,
            I => \N__4648\
        );

    \I__831\ : Odrv12
    port map (
            O => \N__4648\,
            I => \U409_TRANSFER_ACK.N_29\
        );

    \I__830\ : CascadeMux
    port map (
            O => \N__4645\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_3_cascade_\
        );

    \I__829\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4639\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4639\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__827\ : InMux
    port map (
            O => \N__4636\,
            I => \N__4630\
        );

    \I__826\ : InMux
    port map (
            O => \N__4635\,
            I => \N__4630\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4630\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__4627\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_2_cascade_\
        );

    \I__823\ : InMux
    port map (
            O => \N__4624\,
            I => \N__4620\
        );

    \I__822\ : InMux
    port map (
            O => \N__4623\,
            I => \N__4617\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4620\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4617\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__819\ : InMux
    port map (
            O => \N__4612\,
            I => \N__4609\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4609\,
            I => \N__4605\
        );

    \I__817\ : InMux
    port map (
            O => \N__4608\,
            I => \N__4600\
        );

    \I__816\ : Span4Mux_v
    port map (
            O => \N__4605\,
            I => \N__4597\
        );

    \I__815\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4592\
        );

    \I__814\ : InMux
    port map (
            O => \N__4603\,
            I => \N__4592\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__4600\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__812\ : Odrv4
    port map (
            O => \N__4597\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4592\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__810\ : InMux
    port map (
            O => \N__4585\,
            I => \N__4582\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4582\,
            I => \N__4579\
        );

    \I__808\ : Odrv4
    port map (
            O => \N__4579\,
            I => \U409_TRANSFER_ACK.N_47\
        );

    \I__807\ : InMux
    port map (
            O => \N__4576\,
            I => \N__4573\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4573\,
            I => \U409_TRANSFER_ACK.N_142\
        );

    \I__805\ : InMux
    port map (
            O => \N__4570\,
            I => \N__4564\
        );

    \I__804\ : InMux
    port map (
            O => \N__4569\,
            I => \N__4564\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4564\,
            I => \N__4561\
        );

    \I__802\ : Span12Mux_v
    port map (
            O => \N__4561\,
            I => \N__4558\
        );

    \I__801\ : Odrv12
    port map (
            O => \N__4558\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_0\
        );

    \I__800\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4550\
        );

    \I__799\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4547\
        );

    \I__798\ : CascadeMux
    port map (
            O => \N__4553\,
            I => \N__4544\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4550\,
            I => \N__4538\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4547\,
            I => \N__4538\
        );

    \I__795\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4533\
        );

    \I__794\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4533\
        );

    \I__793\ : Span4Mux_v
    port map (
            O => \N__4538\,
            I => \N__4527\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4533\,
            I => \N__4527\
        );

    \I__791\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4524\
        );

    \I__790\ : Span4Mux_v
    port map (
            O => \N__4527\,
            I => \N__4521\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__4524\,
            I => \N__4518\
        );

    \I__788\ : Sp12to4
    port map (
            O => \N__4521\,
            I => \N__4515\
        );

    \I__787\ : Span12Mux_h
    port map (
            O => \N__4518\,
            I => \N__4512\
        );

    \I__786\ : Span12Mux_h
    port map (
            O => \N__4515\,
            I => \N__4509\
        );

    \I__785\ : Span12Mux_v
    port map (
            O => \N__4512\,
            I => \N__4506\
        );

    \I__784\ : Span12Mux_v
    port map (
            O => \N__4509\,
            I => \N__4503\
        );

    \I__783\ : Odrv12
    port map (
            O => \N__4506\,
            I => \TSn_c\
        );

    \I__782\ : Odrv12
    port map (
            O => \N__4503\,
            I => \TSn_c\
        );

    \I__781\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4493\
        );

    \I__780\ : InMux
    port map (
            O => \N__4497\,
            I => \N__4488\
        );

    \I__779\ : InMux
    port map (
            O => \N__4496\,
            I => \N__4488\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4493\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__4488\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__4483\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_cascade_\
        );

    \I__775\ : CEMux
    port map (
            O => \N__4480\,
            I => \N__4477\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4477\,
            I => \N__4474\
        );

    \I__773\ : Span4Mux_h
    port map (
            O => \N__4474\,
            I => \N__4471\
        );

    \I__772\ : Odrv4
    port map (
            O => \N__4471\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_0\
        );

    \I__771\ : IoInMux
    port map (
            O => \N__4468\,
            I => \N__4465\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4465\,
            I => \N__4462\
        );

    \I__769\ : IoSpan4Mux
    port map (
            O => \N__4462\,
            I => \N__4459\
        );

    \I__768\ : Span4Mux_s1_v
    port map (
            O => \N__4459\,
            I => \N__4456\
        );

    \I__767\ : Sp12to4
    port map (
            O => \N__4456\,
            I => \N__4453\
        );

    \I__766\ : Span12Mux_v
    port map (
            O => \N__4453\,
            I => \N__4450\
        );

    \I__765\ : Odrv12
    port map (
            O => \N__4450\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\
        );

    \I__764\ : InMux
    port map (
            O => \N__4447\,
            I => \N__4443\
        );

    \I__763\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4440\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4443\,
            I => \N__4432\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4440\,
            I => \N__4432\
        );

    \I__760\ : InMux
    port map (
            O => \N__4439\,
            I => \N__4429\
        );

    \I__759\ : InMux
    port map (
            O => \N__4438\,
            I => \N__4426\
        );

    \I__758\ : InMux
    port map (
            O => \N__4437\,
            I => \N__4420\
        );

    \I__757\ : Span4Mux_v
    port map (
            O => \N__4432\,
            I => \N__4417\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__4429\,
            I => \N__4412\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4426\,
            I => \N__4412\
        );

    \I__754\ : InMux
    port map (
            O => \N__4425\,
            I => \N__4409\
        );

    \I__753\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4406\
        );

    \I__752\ : InMux
    port map (
            O => \N__4423\,
            I => \N__4403\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4420\,
            I => \N__4400\
        );

    \I__750\ : Span4Mux_h
    port map (
            O => \N__4417\,
            I => \N__4395\
        );

    \I__749\ : Span4Mux_v
    port map (
            O => \N__4412\,
            I => \N__4395\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4409\,
            I => \N__4390\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__4406\,
            I => \N__4390\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4403\,
            I => \N__4386\
        );

    \I__745\ : Span4Mux_v
    port map (
            O => \N__4400\,
            I => \N__4383\
        );

    \I__744\ : Span4Mux_h
    port map (
            O => \N__4395\,
            I => \N__4378\
        );

    \I__743\ : Span4Mux_v
    port map (
            O => \N__4390\,
            I => \N__4378\
        );

    \I__742\ : InMux
    port map (
            O => \N__4389\,
            I => \N__4375\
        );

    \I__741\ : Span12Mux_v
    port map (
            O => \N__4386\,
            I => \N__4366\
        );

    \I__740\ : Sp12to4
    port map (
            O => \N__4383\,
            I => \N__4366\
        );

    \I__739\ : Sp12to4
    port map (
            O => \N__4378\,
            I => \N__4366\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4375\,
            I => \N__4366\
        );

    \I__737\ : Odrv12
    port map (
            O => \N__4366\,
            I => \A_c_21\
        );

    \I__736\ : InMux
    port map (
            O => \N__4363\,
            I => \N__4359\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__4362\,
            I => \N__4356\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__4359\,
            I => \N__4352\
        );

    \I__733\ : InMux
    port map (
            O => \N__4356\,
            I => \N__4349\
        );

    \I__732\ : InMux
    port map (
            O => \N__4355\,
            I => \N__4346\
        );

    \I__731\ : Span4Mux_v
    port map (
            O => \N__4352\,
            I => \N__4343\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4349\,
            I => \N__4338\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__4346\,
            I => \N__4338\
        );

    \I__728\ : Span4Mux_h
    port map (
            O => \N__4343\,
            I => \N__4333\
        );

    \I__727\ : Span4Mux_v
    port map (
            O => \N__4338\,
            I => \N__4333\
        );

    \I__726\ : Sp12to4
    port map (
            O => \N__4333\,
            I => \N__4330\
        );

    \I__725\ : Span12Mux_h
    port map (
            O => \N__4330\,
            I => \N__4327\
        );

    \I__724\ : Span12Mux_v
    port map (
            O => \N__4327\,
            I => \N__4324\
        );

    \I__723\ : Odrv12
    port map (
            O => \N__4324\,
            I => \OVL_c\
        );

    \I__722\ : InMux
    port map (
            O => \N__4321\,
            I => \N__4317\
        );

    \I__721\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4314\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4317\,
            I => \N__4309\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__4314\,
            I => \N__4309\
        );

    \I__718\ : Span4Mux_v
    port map (
            O => \N__4309\,
            I => \N__4305\
        );

    \I__717\ : InMux
    port map (
            O => \N__4308\,
            I => \N__4302\
        );

    \I__716\ : Span4Mux_h
    port map (
            O => \N__4305\,
            I => \N__4297\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4302\,
            I => \N__4297\
        );

    \I__714\ : Odrv4
    port map (
            O => \N__4297\,
            I => \U409_ADDRESS_DECODE_LOWROM_3\
        );

    \I__713\ : CascadeMux
    port map (
            O => \N__4294\,
            I => \N__4291\
        );

    \I__712\ : InMux
    port map (
            O => \N__4291\,
            I => \N__4287\
        );

    \I__711\ : InMux
    port map (
            O => \N__4290\,
            I => \N__4284\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4287\,
            I => \N__4281\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__4284\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__708\ : Odrv4
    port map (
            O => \N__4281\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__707\ : InMux
    port map (
            O => \N__4276\,
            I => \N__4273\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4273\,
            I => \N__4270\
        );

    \I__705\ : Odrv12
    port map (
            O => \N__4270\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__704\ : InMux
    port map (
            O => \N__4267\,
            I => \N__4264\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4264\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23\
        );

    \I__702\ : CascadeMux
    port map (
            O => \N__4261\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_cascade_\
        );

    \I__701\ : CascadeMux
    port map (
            O => \N__4258\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__700\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4252\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__4252\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__4249\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\
        );

    \I__697\ : CascadeMux
    port map (
            O => \N__4246\,
            I => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\
        );

    \I__696\ : IoInMux
    port map (
            O => \N__4243\,
            I => \N__4240\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4240\,
            I => \N__4235\
        );

    \I__694\ : IoInMux
    port map (
            O => \N__4239\,
            I => \N__4232\
        );

    \I__693\ : IoInMux
    port map (
            O => \N__4238\,
            I => \N__4229\
        );

    \I__692\ : Span4Mux_s3_v
    port map (
            O => \N__4235\,
            I => \N__4226\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__4232\,
            I => \N__4221\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4229\,
            I => \N__4221\
        );

    \I__689\ : Span4Mux_v
    port map (
            O => \N__4226\,
            I => \N__4218\
        );

    \I__688\ : Span12Mux_s7_v
    port map (
            O => \N__4221\,
            I => \N__4215\
        );

    \I__687\ : Sp12to4
    port map (
            O => \N__4218\,
            I => \N__4212\
        );

    \I__686\ : Span12Mux_v
    port map (
            O => \N__4215\,
            I => \N__4209\
        );

    \I__685\ : Span12Mux_s7_h
    port map (
            O => \N__4212\,
            I => \N__4206\
        );

    \I__684\ : Span12Mux_h
    port map (
            O => \N__4209\,
            I => \N__4201\
        );

    \I__683\ : Span12Mux_v
    port map (
            O => \N__4206\,
            I => \N__4198\
        );

    \I__682\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4195\
        );

    \I__681\ : InMux
    port map (
            O => \N__4204\,
            I => \N__4192\
        );

    \I__680\ : Odrv12
    port map (
            O => \N__4201\,
            I => \TACK_OUTn\
        );

    \I__679\ : Odrv12
    port map (
            O => \N__4198\,
            I => \TACK_OUTn\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__4195\,
            I => \TACK_OUTn\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4192\,
            I => \TACK_OUTn\
        );

    \I__676\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4177\
        );

    \I__675\ : InMux
    port map (
            O => \N__4182\,
            I => \N__4170\
        );

    \I__674\ : InMux
    port map (
            O => \N__4181\,
            I => \N__4170\
        );

    \I__673\ : InMux
    port map (
            O => \N__4180\,
            I => \N__4170\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4177\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4170\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__670\ : CascadeMux
    port map (
            O => \N__4165\,
            I => \N__4162\
        );

    \I__669\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4156\
        );

    \I__668\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4153\
        );

    \I__667\ : InMux
    port map (
            O => \N__4160\,
            I => \N__4148\
        );

    \I__666\ : InMux
    port map (
            O => \N__4159\,
            I => \N__4148\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4156\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4153\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4148\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__662\ : InMux
    port map (
            O => \N__4141\,
            I => \N__4137\
        );

    \I__661\ : InMux
    port map (
            O => \N__4140\,
            I => \N__4134\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4137\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__4134\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__658\ : InMux
    port map (
            O => \N__4129\,
            I => \N__4126\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__4126\,
            I => \U409_TRANSFER_ACK.N_35\
        );

    \I__656\ : IoInMux
    port map (
            O => \N__4123\,
            I => \N__4120\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__4120\,
            I => \N__4117\
        );

    \I__654\ : IoSpan4Mux
    port map (
            O => \N__4117\,
            I => \N__4114\
        );

    \I__653\ : Sp12to4
    port map (
            O => \N__4114\,
            I => \N__4111\
        );

    \I__652\ : Span12Mux_s6_v
    port map (
            O => \N__4111\,
            I => \N__4108\
        );

    \I__651\ : Span12Mux_v
    port map (
            O => \N__4108\,
            I => \N__4104\
        );

    \I__650\ : InMux
    port map (
            O => \N__4107\,
            I => \N__4101\
        );

    \I__649\ : Odrv12
    port map (
            O => \N__4104\,
            I => \ROMENn_c\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4101\,
            I => \ROMENn_c\
        );

    \I__647\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4092\
        );

    \I__646\ : InMux
    port map (
            O => \N__4095\,
            I => \N__4089\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4092\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4089\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__643\ : InMux
    port map (
            O => \N__4084\,
            I => \N__4078\
        );

    \I__642\ : InMux
    port map (
            O => \N__4083\,
            I => \N__4073\
        );

    \I__641\ : InMux
    port map (
            O => \N__4082\,
            I => \N__4073\
        );

    \I__640\ : InMux
    port map (
            O => \N__4081\,
            I => \N__4070\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4078\,
            I => \N__4063\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__4073\,
            I => \N__4063\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4070\,
            I => \N__4063\
        );

    \I__636\ : Span4Mux_v
    port map (
            O => \N__4063\,
            I => \N__4060\
        );

    \I__635\ : Sp12to4
    port map (
            O => \N__4060\,
            I => \N__4057\
        );

    \I__634\ : Span12Mux_h
    port map (
            O => \N__4057\,
            I => \N__4054\
        );

    \I__633\ : Odrv12
    port map (
            O => \N__4054\,
            I => \TM_c_1\
        );

    \I__632\ : InMux
    port map (
            O => \N__4051\,
            I => \N__4048\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4048\,
            I => \N__4042\
        );

    \I__630\ : InMux
    port map (
            O => \N__4047\,
            I => \N__4037\
        );

    \I__629\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4037\
        );

    \I__628\ : InMux
    port map (
            O => \N__4045\,
            I => \N__4034\
        );

    \I__627\ : Span4Mux_h
    port map (
            O => \N__4042\,
            I => \N__4027\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__4037\,
            I => \N__4027\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4034\,
            I => \N__4027\
        );

    \I__624\ : Span4Mux_v
    port map (
            O => \N__4027\,
            I => \N__4024\
        );

    \I__623\ : Sp12to4
    port map (
            O => \N__4024\,
            I => \N__4021\
        );

    \I__622\ : Span12Mux_h
    port map (
            O => \N__4021\,
            I => \N__4018\
        );

    \I__621\ : Odrv12
    port map (
            O => \N__4018\,
            I => \TM_c_0\
        );

    \I__620\ : InMux
    port map (
            O => \N__4015\,
            I => \N__4007\
        );

    \I__619\ : InMux
    port map (
            O => \N__4014\,
            I => \N__4007\
        );

    \I__618\ : InMux
    port map (
            O => \N__4013\,
            I => \N__4004\
        );

    \I__617\ : InMux
    port map (
            O => \N__4012\,
            I => \N__4001\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4007\,
            I => \N__3998\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__4004\,
            I => \N__3995\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__4001\,
            I => \N__3990\
        );

    \I__613\ : Span4Mux_v
    port map (
            O => \N__3998\,
            I => \N__3984\
        );

    \I__612\ : Span4Mux_v
    port map (
            O => \N__3995\,
            I => \N__3984\
        );

    \I__611\ : InMux
    port map (
            O => \N__3994\,
            I => \N__3981\
        );

    \I__610\ : InMux
    port map (
            O => \N__3993\,
            I => \N__3978\
        );

    \I__609\ : Span4Mux_v
    port map (
            O => \N__3990\,
            I => \N__3975\
        );

    \I__608\ : InMux
    port map (
            O => \N__3989\,
            I => \N__3972\
        );

    \I__607\ : Sp12to4
    port map (
            O => \N__3984\,
            I => \N__3965\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3981\,
            I => \N__3965\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3978\,
            I => \N__3965\
        );

    \I__604\ : Sp12to4
    port map (
            O => \N__3975\,
            I => \N__3960\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3972\,
            I => \N__3960\
        );

    \I__602\ : Odrv12
    port map (
            O => \N__3965\,
            I => \A_c_23\
        );

    \I__601\ : Odrv12
    port map (
            O => \N__3960\,
            I => \A_c_23\
        );

    \I__600\ : InMux
    port map (
            O => \N__3955\,
            I => \N__3950\
        );

    \I__599\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3947\
        );

    \I__598\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3944\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3950\,
            I => \N__3935\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3947\,
            I => \N__3935\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3944\,
            I => \N__3932\
        );

    \I__594\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3929\
        );

    \I__593\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3926\
        );

    \I__592\ : InMux
    port map (
            O => \N__3941\,
            I => \N__3921\
        );

    \I__591\ : InMux
    port map (
            O => \N__3940\,
            I => \N__3921\
        );

    \I__590\ : Span4Mux_h
    port map (
            O => \N__3935\,
            I => \N__3913\
        );

    \I__589\ : Span4Mux_v
    port map (
            O => \N__3932\,
            I => \N__3913\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3929\,
            I => \N__3913\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3926\,
            I => \N__3908\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__3921\,
            I => \N__3908\
        );

    \I__585\ : InMux
    port map (
            O => \N__3920\,
            I => \N__3905\
        );

    \I__584\ : Span4Mux_h
    port map (
            O => \N__3913\,
            I => \N__3902\
        );

    \I__583\ : Sp12to4
    port map (
            O => \N__3908\,
            I => \N__3897\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3905\,
            I => \N__3897\
        );

    \I__581\ : Span4Mux_v
    port map (
            O => \N__3902\,
            I => \N__3894\
        );

    \I__580\ : Span12Mux_v
    port map (
            O => \N__3897\,
            I => \N__3891\
        );

    \I__579\ : Span4Mux_v
    port map (
            O => \N__3894\,
            I => \N__3888\
        );

    \I__578\ : Odrv12
    port map (
            O => \N__3891\,
            I => \A_c_22\
        );

    \I__577\ : Odrv4
    port map (
            O => \N__3888\,
            I => \A_c_22\
        );

    \I__576\ : IoInMux
    port map (
            O => \N__3883\,
            I => \N__3880\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3880\,
            I => \N__3877\
        );

    \I__574\ : Span4Mux_s3_v
    port map (
            O => \N__3877\,
            I => \N__3874\
        );

    \I__573\ : Span4Mux_h
    port map (
            O => \N__3874\,
            I => \N__3871\
        );

    \I__572\ : Span4Mux_h
    port map (
            O => \N__3871\,
            I => \N__3868\
        );

    \I__571\ : Span4Mux_h
    port map (
            O => \N__3868\,
            I => \N__3865\
        );

    \I__570\ : Span4Mux_h
    port map (
            O => \N__3865\,
            I => \N__3862\
        );

    \I__569\ : Span4Mux_v
    port map (
            O => \N__3862\,
            I => \N__3859\
        );

    \I__568\ : Odrv4
    port map (
            O => \N__3859\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\
        );

    \I__567\ : InMux
    port map (
            O => \N__3856\,
            I => \N__3847\
        );

    \I__566\ : InMux
    port map (
            O => \N__3855\,
            I => \N__3847\
        );

    \I__565\ : InMux
    port map (
            O => \N__3854\,
            I => \N__3844\
        );

    \I__564\ : InMux
    port map (
            O => \N__3853\,
            I => \N__3839\
        );

    \I__563\ : InMux
    port map (
            O => \N__3852\,
            I => \N__3839\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3847\,
            I => \N__3836\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3844\,
            I => \N__3833\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3839\,
            I => \N__3830\
        );

    \I__559\ : Span4Mux_v
    port map (
            O => \N__3836\,
            I => \N__3827\
        );

    \I__558\ : Span4Mux_v
    port map (
            O => \N__3833\,
            I => \N__3822\
        );

    \I__557\ : Span4Mux_h
    port map (
            O => \N__3830\,
            I => \N__3822\
        );

    \I__556\ : Span4Mux_h
    port map (
            O => \N__3827\,
            I => \N__3819\
        );

    \I__555\ : Span4Mux_h
    port map (
            O => \N__3822\,
            I => \N__3816\
        );

    \I__554\ : Odrv4
    port map (
            O => \N__3819\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0\
        );

    \I__553\ : Odrv4
    port map (
            O => \N__3816\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0\
        );

    \I__552\ : CascadeMux
    port map (
            O => \N__3811\,
            I => \N__3808\
        );

    \I__551\ : InMux
    port map (
            O => \N__3808\,
            I => \N__3802\
        );

    \I__550\ : InMux
    port map (
            O => \N__3807\,
            I => \N__3802\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3802\,
            I => \N__3799\
        );

    \I__548\ : Span4Mux_v
    port map (
            O => \N__3799\,
            I => \N__3796\
        );

    \I__547\ : Odrv4
    port map (
            O => \N__3796\,
            I => \U409_ADDRESS_DECODE.un2_REGSPACEn_0_0\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__3793\,
            I => \N__3789\
        );

    \I__545\ : InMux
    port map (
            O => \N__3792\,
            I => \N__3784\
        );

    \I__544\ : InMux
    port map (
            O => \N__3789\,
            I => \N__3784\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3784\,
            I => \N__3781\
        );

    \I__542\ : Odrv4
    port map (
            O => \N__3781\,
            I => \U409_ADDRESS_DECODE.REG_SPACE_3_0\
        );

    \I__541\ : InMux
    port map (
            O => \N__3778\,
            I => \N__3772\
        );

    \I__540\ : InMux
    port map (
            O => \N__3777\,
            I => \N__3772\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3772\,
            I => \U409_ADDRESS_DECODE.REG_SPACEZ0Z_2\
        );

    \I__538\ : InMux
    port map (
            O => \N__3769\,
            I => \N__3766\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3766\,
            I => \N__3762\
        );

    \I__536\ : InMux
    port map (
            O => \N__3765\,
            I => \N__3759\
        );

    \I__535\ : Span4Mux_h
    port map (
            O => \N__3762\,
            I => \N__3754\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3759\,
            I => \N__3754\
        );

    \I__533\ : Odrv4
    port map (
            O => \N__3754\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn\
        );

    \I__532\ : IoInMux
    port map (
            O => \N__3751\,
            I => \N__3748\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3748\,
            I => \N__3745\
        );

    \I__530\ : Span12Mux_s10_v
    port map (
            O => \N__3745\,
            I => \N__3742\
        );

    \I__529\ : Odrv12
    port map (
            O => \N__3742\,
            I => \PORTSIZE_0_i\
        );

    \I__528\ : CascadeMux
    port map (
            O => \N__3739\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0_cascade_\
        );

    \I__527\ : CEMux
    port map (
            O => \N__3736\,
            I => \N__3733\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3733\,
            I => \N__3730\
        );

    \I__525\ : Span4Mux_v
    port map (
            O => \N__3730\,
            I => \N__3727\
        );

    \I__524\ : Odrv4
    port map (
            O => \N__3727\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_0\
        );

    \I__523\ : InMux
    port map (
            O => \N__3724\,
            I => \N__3721\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3721\,
            I => \N__3718\
        );

    \I__521\ : Span4Mux_v
    port map (
            O => \N__3718\,
            I => \N__3715\
        );

    \I__520\ : IoSpan4Mux
    port map (
            O => \N__3715\,
            I => \N__3712\
        );

    \I__519\ : Odrv4
    port map (
            O => \N__3712\,
            I => \TT_c_1\
        );

    \I__518\ : InMux
    port map (
            O => \N__3709\,
            I => \N__3706\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3706\,
            I => \N__3703\
        );

    \I__516\ : Span4Mux_h
    port map (
            O => \N__3703\,
            I => \N__3700\
        );

    \I__515\ : Span4Mux_v
    port map (
            O => \N__3700\,
            I => \N__3697\
        );

    \I__514\ : Odrv4
    port map (
            O => \N__3697\,
            I => \TT_c_0\
        );

    \I__513\ : InMux
    port map (
            O => \N__3694\,
            I => \N__3691\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3691\,
            I => \N__3688\
        );

    \I__511\ : Odrv12
    port map (
            O => \N__3688\,
            I => \U409_ADDRESS_DECODE_AUTOVECTOR_2\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__3685\,
            I => \U409_ADDRESS_DECODE_LOWROM_2_cascade_\
        );

    \I__509\ : InMux
    port map (
            O => \N__3682\,
            I => \N__3679\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3679\,
            I => \U409_TRANSFER_ACK.N_45\
        );

    \I__507\ : CascadeMux
    port map (
            O => \N__3676\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2Z0Z_1_cascade_\
        );

    \I__506\ : CascadeMux
    port map (
            O => \N__3673\,
            I => \N__3670\
        );

    \I__505\ : InMux
    port map (
            O => \N__3670\,
            I => \N__3667\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3667\,
            I => \N__3663\
        );

    \I__503\ : InMux
    port map (
            O => \N__3666\,
            I => \N__3660\
        );

    \I__502\ : Odrv4
    port map (
            O => \N__3663\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3660\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2\
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__3655\,
            I => \N__3651\
        );

    \I__499\ : InMux
    port map (
            O => \N__3654\,
            I => \N__3648\
        );

    \I__498\ : InMux
    port map (
            O => \N__3651\,
            I => \N__3642\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3648\,
            I => \N__3639\
        );

    \I__496\ : InMux
    port map (
            O => \N__3647\,
            I => \N__3634\
        );

    \I__495\ : InMux
    port map (
            O => \N__3646\,
            I => \N__3634\
        );

    \I__494\ : InMux
    port map (
            O => \N__3645\,
            I => \N__3631\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3642\,
            I => \N__3628\
        );

    \I__492\ : Span4Mux_v
    port map (
            O => \N__3639\,
            I => \N__3625\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3634\,
            I => \N__3620\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3631\,
            I => \N__3620\
        );

    \I__489\ : Span4Mux_v
    port map (
            O => \N__3628\,
            I => \N__3617\
        );

    \I__488\ : Span4Mux_h
    port map (
            O => \N__3625\,
            I => \N__3612\
        );

    \I__487\ : Span4Mux_v
    port map (
            O => \N__3620\,
            I => \N__3612\
        );

    \I__486\ : Sp12to4
    port map (
            O => \N__3617\,
            I => \N__3607\
        );

    \I__485\ : Sp12to4
    port map (
            O => \N__3612\,
            I => \N__3607\
        );

    \I__484\ : Span12Mux_h
    port map (
            O => \N__3607\,
            I => \N__3604\
        );

    \I__483\ : Span12Mux_v
    port map (
            O => \N__3604\,
            I => \N__3601\
        );

    \I__482\ : Odrv12
    port map (
            O => \N__3601\,
            I => \A_c_18\
        );

    \I__481\ : InMux
    port map (
            O => \N__3598\,
            I => \N__3590\
        );

    \I__480\ : InMux
    port map (
            O => \N__3597\,
            I => \N__3590\
        );

    \I__479\ : InMux
    port map (
            O => \N__3596\,
            I => \N__3585\
        );

    \I__478\ : InMux
    port map (
            O => \N__3595\,
            I => \N__3585\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3590\,
            I => \N__3580\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3585\,
            I => \N__3576\
        );

    \I__475\ : InMux
    port map (
            O => \N__3584\,
            I => \N__3573\
        );

    \I__474\ : InMux
    port map (
            O => \N__3583\,
            I => \N__3570\
        );

    \I__473\ : Span4Mux_v
    port map (
            O => \N__3580\,
            I => \N__3566\
        );

    \I__472\ : InMux
    port map (
            O => \N__3579\,
            I => \N__3563\
        );

    \I__471\ : Span4Mux_v
    port map (
            O => \N__3576\,
            I => \N__3560\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3573\,
            I => \N__3557\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3570\,
            I => \N__3554\
        );

    \I__468\ : InMux
    port map (
            O => \N__3569\,
            I => \N__3551\
        );

    \I__467\ : Sp12to4
    port map (
            O => \N__3566\,
            I => \N__3546\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3563\,
            I => \N__3546\
        );

    \I__465\ : Span4Mux_h
    port map (
            O => \N__3560\,
            I => \N__3539\
        );

    \I__464\ : Span4Mux_v
    port map (
            O => \N__3557\,
            I => \N__3539\
        );

    \I__463\ : Span4Mux_v
    port map (
            O => \N__3554\,
            I => \N__3539\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3551\,
            I => \N__3536\
        );

    \I__461\ : Span12Mux_h
    port map (
            O => \N__3546\,
            I => \N__3529\
        );

    \I__460\ : Sp12to4
    port map (
            O => \N__3539\,
            I => \N__3529\
        );

    \I__459\ : Span12Mux_v
    port map (
            O => \N__3536\,
            I => \N__3529\
        );

    \I__458\ : Odrv12
    port map (
            O => \N__3529\,
            I => \A_c_20\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__3526\,
            I => \N__3522\
        );

    \I__456\ : InMux
    port map (
            O => \N__3525\,
            I => \N__3518\
        );

    \I__455\ : InMux
    port map (
            O => \N__3522\,
            I => \N__3515\
        );

    \I__454\ : InMux
    port map (
            O => \N__3521\,
            I => \N__3512\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3518\,
            I => \N__3503\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3515\,
            I => \N__3503\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__3512\,
            I => \N__3503\
        );

    \I__450\ : InMux
    port map (
            O => \N__3511\,
            I => \N__3500\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__3510\,
            I => \N__3495\
        );

    \I__448\ : Span4Mux_v
    port map (
            O => \N__3503\,
            I => \N__3492\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3500\,
            I => \N__3489\
        );

    \I__446\ : InMux
    port map (
            O => \N__3499\,
            I => \N__3484\
        );

    \I__445\ : InMux
    port map (
            O => \N__3498\,
            I => \N__3484\
        );

    \I__444\ : InMux
    port map (
            O => \N__3495\,
            I => \N__3481\
        );

    \I__443\ : Span4Mux_v
    port map (
            O => \N__3492\,
            I => \N__3478\
        );

    \I__442\ : Span4Mux_h
    port map (
            O => \N__3489\,
            I => \N__3471\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3484\,
            I => \N__3471\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3481\,
            I => \N__3471\
        );

    \I__439\ : Span4Mux_v
    port map (
            O => \N__3478\,
            I => \N__3468\
        );

    \I__438\ : Span4Mux_h
    port map (
            O => \N__3471\,
            I => \N__3465\
        );

    \I__437\ : Sp12to4
    port map (
            O => \N__3468\,
            I => \N__3462\
        );

    \I__436\ : Sp12to4
    port map (
            O => \N__3465\,
            I => \N__3459\
        );

    \I__435\ : Span12Mux_h
    port map (
            O => \N__3462\,
            I => \N__3454\
        );

    \I__434\ : Span12Mux_v
    port map (
            O => \N__3459\,
            I => \N__3454\
        );

    \I__433\ : Odrv12
    port map (
            O => \N__3454\,
            I => \A_c_19\
        );

    \I__432\ : CascadeMux
    port map (
            O => \N__3451\,
            I => \N__3448\
        );

    \I__431\ : InMux
    port map (
            O => \N__3448\,
            I => \N__3442\
        );

    \I__430\ : InMux
    port map (
            O => \N__3447\,
            I => \N__3442\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3442\,
            I => \N__3438\
        );

    \I__428\ : InMux
    port map (
            O => \N__3441\,
            I => \N__3435\
        );

    \I__427\ : Span4Mux_v
    port map (
            O => \N__3438\,
            I => \N__3432\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__3435\,
            I => \N__3429\
        );

    \I__425\ : Span4Mux_h
    port map (
            O => \N__3432\,
            I => \N__3423\
        );

    \I__424\ : Span4Mux_v
    port map (
            O => \N__3429\,
            I => \N__3423\
        );

    \I__423\ : InMux
    port map (
            O => \N__3428\,
            I => \N__3420\
        );

    \I__422\ : Sp12to4
    port map (
            O => \N__3423\,
            I => \N__3417\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3420\,
            I => \N__3414\
        );

    \I__420\ : Span12Mux_s5_h
    port map (
            O => \N__3417\,
            I => \N__3409\
        );

    \I__419\ : Span12Mux_v
    port map (
            O => \N__3414\,
            I => \N__3409\
        );

    \I__418\ : Span12Mux_v
    port map (
            O => \N__3409\,
            I => \N__3406\
        );

    \I__417\ : Odrv12
    port map (
            O => \N__3406\,
            I => \A_c_17\
        );

    \I__416\ : InMux
    port map (
            O => \N__3403\,
            I => \N__3400\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3400\,
            I => \N__3397\
        );

    \I__414\ : Span4Mux_v
    port map (
            O => \N__3397\,
            I => \N__3393\
        );

    \I__413\ : InMux
    port map (
            O => \N__3396\,
            I => \N__3390\
        );

    \I__412\ : Odrv4
    port map (
            O => \N__3393\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__3390\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0\
        );

    \I__410\ : CascadeMux
    port map (
            O => \N__3385\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_\
        );

    \I__409\ : CascadeMux
    port map (
            O => \N__3382\,
            I => \N__3378\
        );

    \I__408\ : InMux
    port map (
            O => \N__3381\,
            I => \N__3373\
        );

    \I__407\ : InMux
    port map (
            O => \N__3378\,
            I => \N__3373\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3373\,
            I => \N__3370\
        );

    \I__405\ : Span4Mux_h
    port map (
            O => \N__3370\,
            I => \N__3367\
        );

    \I__404\ : Odrv4
    port map (
            O => \N__3367\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_4\
        );

    \I__403\ : InMux
    port map (
            O => \N__3364\,
            I => \N__3358\
        );

    \I__402\ : InMux
    port map (
            O => \N__3363\,
            I => \N__3358\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__3358\,
            I => \N__3355\
        );

    \I__400\ : Span4Mux_v
    port map (
            O => \N__3355\,
            I => \N__3352\
        );

    \I__399\ : Odrv4
    port map (
            O => \N__3352\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_5\
        );

    \I__398\ : CascadeMux
    port map (
            O => \N__3349\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_0_cascade_\
        );

    \I__397\ : InMux
    port map (
            O => \N__3346\,
            I => \N__3343\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3343\,
            I => \N__3340\
        );

    \I__395\ : Span4Mux_h
    port map (
            O => \N__3340\,
            I => \N__3337\
        );

    \I__394\ : Span4Mux_v
    port map (
            O => \N__3337\,
            I => \N__3334\
        );

    \I__393\ : Span4Mux_v
    port map (
            O => \N__3334\,
            I => \N__3331\
        );

    \I__392\ : Odrv4
    port map (
            O => \N__3331\,
            I => \RnW_c\
        );

    \I__391\ : IoInMux
    port map (
            O => \N__3328\,
            I => \N__3325\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3325\,
            I => \N__3319\
        );

    \I__389\ : IoInMux
    port map (
            O => \N__3324\,
            I => \N__3316\
        );

    \I__388\ : IoInMux
    port map (
            O => \N__3323\,
            I => \N__3313\
        );

    \I__387\ : IoInMux
    port map (
            O => \N__3322\,
            I => \N__3310\
        );

    \I__386\ : IoSpan4Mux
    port map (
            O => \N__3319\,
            I => \N__3300\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__3316\,
            I => \N__3300\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3313\,
            I => \N__3300\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3310\,
            I => \N__3297\
        );

    \I__382\ : IoInMux
    port map (
            O => \N__3309\,
            I => \N__3294\
        );

    \I__381\ : IoInMux
    port map (
            O => \N__3308\,
            I => \N__3291\
        );

    \I__380\ : IoInMux
    port map (
            O => \N__3307\,
            I => \N__3288\
        );

    \I__379\ : IoSpan4Mux
    port map (
            O => \N__3300\,
            I => \N__3281\
        );

    \I__378\ : IoSpan4Mux
    port map (
            O => \N__3297\,
            I => \N__3281\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__3294\,
            I => \N__3281\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__3291\,
            I => \N__3276\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__3288\,
            I => \N__3276\
        );

    \I__374\ : IoSpan4Mux
    port map (
            O => \N__3281\,
            I => \N__3270\
        );

    \I__373\ : IoSpan4Mux
    port map (
            O => \N__3276\,
            I => \N__3270\
        );

    \I__372\ : IoInMux
    port map (
            O => \N__3275\,
            I => \N__3267\
        );

    \I__371\ : Sp12to4
    port map (
            O => \N__3270\,
            I => \N__3262\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__3267\,
            I => \N__3262\
        );

    \I__369\ : Span12Mux_s3_v
    port map (
            O => \N__3262\,
            I => \N__3259\
        );

    \I__368\ : Span12Mux_v
    port map (
            O => \N__3259\,
            I => \N__3256\
        );

    \I__367\ : Odrv12
    port map (
            O => \N__3256\,
            I => \D_1_i\
        );

    \I__366\ : IoInMux
    port map (
            O => \N__3253\,
            I => \N__3250\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__3250\,
            I => \N__3247\
        );

    \I__364\ : IoSpan4Mux
    port map (
            O => \N__3247\,
            I => \N__3244\
        );

    \I__363\ : Span4Mux_s2_h
    port map (
            O => \N__3244\,
            I => \N__3241\
        );

    \I__362\ : Sp12to4
    port map (
            O => \N__3241\,
            I => \N__3238\
        );

    \I__361\ : Span12Mux_s11_h
    port map (
            O => \N__3238\,
            I => \N__3235\
        );

    \I__360\ : Span12Mux_h
    port map (
            O => \N__3235\,
            I => \N__3232\
        );

    \I__359\ : Span12Mux_v
    port map (
            O => \N__3232\,
            I => \N__3229\
        );

    \I__358\ : Odrv12
    port map (
            O => \N__3229\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn_i\
        );

    \I__357\ : InMux
    port map (
            O => \N__3226\,
            I => \N__3223\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__3223\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3\
        );

    \I__355\ : CascadeMux
    port map (
            O => \N__3220\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3_cascade_\
        );

    \I__354\ : InMux
    port map (
            O => \N__3217\,
            I => \N__3214\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__3214\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_0\
        );

    \I__352\ : InMux
    port map (
            O => \N__3211\,
            I => \N__3208\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__3208\,
            I => \N__3205\
        );

    \I__350\ : Span4Mux_v
    port map (
            O => \N__3205\,
            I => \N__3202\
        );

    \I__349\ : Odrv4
    port map (
            O => \N__3202\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5\
        );

    \I__348\ : CascadeMux
    port map (
            O => \N__3199\,
            I => \U409_ADDRESS_DECODE_LOWROM_3_cascade_\
        );

    \I__347\ : InMux
    port map (
            O => \N__3196\,
            I => \N__3193\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__3193\,
            I => \N__3190\
        );

    \I__345\ : Odrv4
    port map (
            O => \N__3190\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3\
        );

    \I__344\ : CascadeMux
    port map (
            O => \N__3187\,
            I => \N__3184\
        );

    \I__343\ : InMux
    port map (
            O => \N__3184\,
            I => \N__3181\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3181\,
            I => \N__3178\
        );

    \I__341\ : Span4Mux_v
    port map (
            O => \N__3178\,
            I => \N__3175\
        );

    \I__340\ : Odrv4
    port map (
            O => \N__3175\,
            I => \U409_ADDRESS_DECODE_AUTOVECTOR_3\
        );

    \I__339\ : InMux
    port map (
            O => \N__3172\,
            I => \N__3169\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__3169\,
            I => \N__3166\
        );

    \I__337\ : Odrv4
    port map (
            O => \N__3166\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\
        );

    \I__336\ : CascadeMux
    port map (
            O => \N__3163\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_\
        );

    \I__335\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3154\
        );

    \I__334\ : InMux
    port map (
            O => \N__3159\,
            I => \N__3154\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__3154\,
            I => \N__3151\
        );

    \I__332\ : Span4Mux_v
    port map (
            O => \N__3151\,
            I => \N__3148\
        );

    \I__331\ : Sp12to4
    port map (
            O => \N__3148\,
            I => \N__3145\
        );

    \I__330\ : Odrv12
    port map (
            O => \N__3145\,
            I => \A_c_31\
        );

    \I__329\ : InMux
    port map (
            O => \N__3142\,
            I => \N__3136\
        );

    \I__328\ : InMux
    port map (
            O => \N__3141\,
            I => \N__3136\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__3136\,
            I => \N__3133\
        );

    \I__326\ : Span4Mux_v
    port map (
            O => \N__3133\,
            I => \N__3130\
        );

    \I__325\ : Span4Mux_h
    port map (
            O => \N__3130\,
            I => \N__3127\
        );

    \I__324\ : Odrv4
    port map (
            O => \N__3127\,
            I => \A_c_30\
        );

    \I__323\ : CascadeMux
    port map (
            O => \N__3124\,
            I => \N__3120\
        );

    \I__322\ : InMux
    port map (
            O => \N__3123\,
            I => \N__3115\
        );

    \I__321\ : InMux
    port map (
            O => \N__3120\,
            I => \N__3115\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__3115\,
            I => \N__3112\
        );

    \I__319\ : Span4Mux_v
    port map (
            O => \N__3112\,
            I => \N__3109\
        );

    \I__318\ : Span4Mux_v
    port map (
            O => \N__3109\,
            I => \N__3106\
        );

    \I__317\ : Sp12to4
    port map (
            O => \N__3106\,
            I => \N__3103\
        );

    \I__316\ : Odrv12
    port map (
            O => \N__3103\,
            I => \A_c_28\
        );

    \I__315\ : InMux
    port map (
            O => \N__3100\,
            I => \N__3094\
        );

    \I__314\ : InMux
    port map (
            O => \N__3099\,
            I => \N__3094\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__3094\,
            I => \N__3091\
        );

    \I__312\ : Span4Mux_h
    port map (
            O => \N__3091\,
            I => \N__3088\
        );

    \I__311\ : Span4Mux_v
    port map (
            O => \N__3088\,
            I => \N__3085\
        );

    \I__310\ : Odrv4
    port map (
            O => \N__3085\,
            I => \A_c_29\
        );

    \I__309\ : CascadeMux
    port map (
            O => \N__3082\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_0Z0Z_1_cascade_\
        );

    \I__308\ : CascadeMux
    port map (
            O => \N__3079\,
            I => \N__3076\
        );

    \I__307\ : InMux
    port map (
            O => \N__3076\,
            I => \N__3072\
        );

    \I__306\ : InMux
    port map (
            O => \N__3075\,
            I => \N__3069\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__3072\,
            I => \N__3064\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__3069\,
            I => \N__3064\
        );

    \I__303\ : Span4Mux_h
    port map (
            O => \N__3064\,
            I => \N__3061\
        );

    \I__302\ : Span4Mux_v
    port map (
            O => \N__3061\,
            I => \N__3058\
        );

    \I__301\ : Sp12to4
    port map (
            O => \N__3058\,
            I => \N__3055\
        );

    \I__300\ : Span12Mux_v
    port map (
            O => \N__3055\,
            I => \N__3052\
        );

    \I__299\ : Odrv12
    port map (
            O => \N__3052\,
            I => \A_c_16\
        );

    \I__298\ : CascadeMux
    port map (
            O => \N__3049\,
            I => \U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0_cascade_\
        );

    \I__297\ : CascadeMux
    port map (
            O => \N__3046\,
            I => \N__3043\
        );

    \I__296\ : InMux
    port map (
            O => \N__3043\,
            I => \N__3037\
        );

    \I__295\ : InMux
    port map (
            O => \N__3042\,
            I => \N__3037\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__3037\,
            I => \N__3034\
        );

    \I__293\ : Span4Mux_v
    port map (
            O => \N__3034\,
            I => \N__3031\
        );

    \I__292\ : Span4Mux_h
    port map (
            O => \N__3031\,
            I => \N__3028\
        );

    \I__291\ : Odrv4
    port map (
            O => \N__3028\,
            I => \A_c_27\
        );

    \I__290\ : CascadeMux
    port map (
            O => \N__3025\,
            I => \N__3021\
        );

    \I__289\ : InMux
    port map (
            O => \N__3024\,
            I => \N__3016\
        );

    \I__288\ : InMux
    port map (
            O => \N__3021\,
            I => \N__3016\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__3016\,
            I => \N__3013\
        );

    \I__286\ : Span4Mux_v
    port map (
            O => \N__3013\,
            I => \N__3010\
        );

    \I__285\ : Span4Mux_v
    port map (
            O => \N__3010\,
            I => \N__3007\
        );

    \I__284\ : Sp12to4
    port map (
            O => \N__3007\,
            I => \N__3004\
        );

    \I__283\ : Odrv12
    port map (
            O => \N__3004\,
            I => \A_c_26\
        );

    \I__282\ : InMux
    port map (
            O => \N__3001\,
            I => \N__2995\
        );

    \I__281\ : InMux
    port map (
            O => \N__3000\,
            I => \N__2995\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__2995\,
            I => \N__2992\
        );

    \I__279\ : Span4Mux_v
    port map (
            O => \N__2992\,
            I => \N__2989\
        );

    \I__278\ : Sp12to4
    port map (
            O => \N__2989\,
            I => \N__2986\
        );

    \I__277\ : Odrv12
    port map (
            O => \N__2986\,
            I => \A_c_25\
        );

    \I__276\ : InMux
    port map (
            O => \N__2983\,
            I => \N__2980\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2980\,
            I => \N__2976\
        );

    \I__274\ : InMux
    port map (
            O => \N__2979\,
            I => \N__2973\
        );

    \I__273\ : Span4Mux_v
    port map (
            O => \N__2976\,
            I => \N__2968\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2973\,
            I => \N__2968\
        );

    \I__271\ : Span4Mux_h
    port map (
            O => \N__2968\,
            I => \N__2965\
        );

    \I__270\ : Span4Mux_v
    port map (
            O => \N__2965\,
            I => \N__2962\
        );

    \I__269\ : Odrv4
    port map (
            O => \N__2962\,
            I => \A_c_24\
        );

    \I__268\ : ClkMux
    port map (
            O => \N__2959\,
            I => \N__2920\
        );

    \I__267\ : ClkMux
    port map (
            O => \N__2958\,
            I => \N__2920\
        );

    \I__266\ : ClkMux
    port map (
            O => \N__2957\,
            I => \N__2920\
        );

    \I__265\ : ClkMux
    port map (
            O => \N__2956\,
            I => \N__2920\
        );

    \I__264\ : ClkMux
    port map (
            O => \N__2955\,
            I => \N__2920\
        );

    \I__263\ : ClkMux
    port map (
            O => \N__2954\,
            I => \N__2920\
        );

    \I__262\ : ClkMux
    port map (
            O => \N__2953\,
            I => \N__2920\
        );

    \I__261\ : ClkMux
    port map (
            O => \N__2952\,
            I => \N__2920\
        );

    \I__260\ : ClkMux
    port map (
            O => \N__2951\,
            I => \N__2920\
        );

    \I__259\ : ClkMux
    port map (
            O => \N__2950\,
            I => \N__2920\
        );

    \I__258\ : ClkMux
    port map (
            O => \N__2949\,
            I => \N__2920\
        );

    \I__257\ : ClkMux
    port map (
            O => \N__2948\,
            I => \N__2920\
        );

    \I__256\ : ClkMux
    port map (
            O => \N__2947\,
            I => \N__2920\
        );

    \I__255\ : GlobalMux
    port map (
            O => \N__2920\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            I => \N__2957\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            I => \N__2951\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            I => \N__2948\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            I => \N__2947\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            I => \N__2950\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            I => \N__2958\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            I => \N__2953\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            I => \N__2949\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC_net\,
            I => \N__2959\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\,
            I => \N__2956\
        );

    \INVU409_TRANSFER_ACK.TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            I => \N__2955\
        );

    \INVU409_TRANSFER_ACK.TACK_OUTnC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            I => \N__2954\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC_net\,
            I => \N__2952\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_11_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__3001\,
            in1 => \N__3024\,
            in2 => \N__3046\,
            in3 => \N__6207\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_4_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2983\,
            in1 => \N__3042\,
            in2 => \N__3025\,
            in3 => \N__3000\,
            lcout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__3160\,
            in1 => \N__3142\,
            in2 => \_gnd_net_\,
            in3 => \N__2979\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__3100\,
            in1 => \N__3172\,
            in2 => \N__3163\,
            in3 => \N__3123\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_5_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3159\,
            in1 => \N__3141\,
            in2 => \N__3124\,
            in3 => \N__3099\,
            lcout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_0_1_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4424\,
            in1 => \N__3569\,
            in2 => \N__3510\,
            in3 => \N__3645\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.CIA_SPACE_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_0_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__3075\,
            in1 => \_gnd_net_\,
            in2 => \N__3082\,
            in3 => \N__3428\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3498\,
            in1 => \N__3646\,
            in2 => \N__3079\,
            in3 => \N__3441\,
            lcout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__3953\,
            in1 => \N__4425\,
            in2 => \_gnd_net_\,
            in3 => \N__4012\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111001111"
        )
    port map (
            in0 => \N__3499\,
            in1 => \N__3583\,
            in2 => \N__3049\,
            in3 => \N__3647\,
            lcout => \U409_ADDRESS_DECODE.un2_REGSPACEn_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4389\,
            in1 => \N__3584\,
            in2 => \N__3382\,
            in3 => \N__3363\,
            lcout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_0_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3396\,
            in1 => \N__3989\,
            in2 => \_gnd_net_\,
            in3 => \N__3943\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_3_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3381\,
            in1 => \N__3364\,
            in2 => \N__3349\,
            in3 => \N__6242\,
            lcout => \U409_ADDRESS_DECODE_AUTOVECTOR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.D_1_i_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__3346\,
            in1 => \N__6326\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \D_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__3941\,
            in1 => \N__3598\,
            in2 => \N__3673\,
            in3 => \N__3226\,
            lcout => \U409_ADDRESS_DECODE_un1_RTC_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__3511\,
            in1 => \N__4437\,
            in2 => \N__3655\,
            in3 => \N__3854\,
            lcout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3\,
            ltout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3940\,
            in1 => \N__3597\,
            in2 => \N__3220\,
            in3 => \N__3666\,
            lcout => \U409_ADDRESS_DECODE_un1_RTC_ENn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__4045\,
            in1 => \N__4081\,
            in2 => \_gnd_net_\,
            in3 => \N__6243\,
            lcout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_9_0_a2_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3993\,
            in2 => \_gnd_net_\,
            in3 => \N__3954\,
            lcout => \U409_ADDRESS_DECODE_LOWROM_3\,
            ltout => \U409_ADDRESS_DECODE_LOWROM_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3217\,
            in1 => \N__3211\,
            in2 => \N__3199\,
            in3 => \N__3196\,
            lcout => \AUTOCONFIG_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__6244\,
            in1 => \N__3765\,
            in2 => \N__3187\,
            in3 => \N__3694\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_2_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3724\,
            in2 => \_gnd_net_\,
            in3 => \N__3709\,
            lcout => \U409_ADDRESS_DECODE_AUTOVECTOR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_8_0_a2_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4439\,
            in2 => \_gnd_net_\,
            in3 => \N__3579\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE_LOWROM_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__3521\,
            in1 => \N__4308\,
            in2 => \N__3685\,
            in3 => \N__4363\,
            lcout => \U409_TRANSFER_ACK.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2_1_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3596\,
            in1 => \N__4438\,
            in2 => \_gnd_net_\,
            in3 => \N__3942\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__3682\,
            in1 => \N__3525\,
            in2 => \N__3676\,
            in3 => \N__4015\,
            lcout => \U409_TRANSFER_ACK.N_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__4014\,
            in1 => \N__4084\,
            in2 => \N__3451\,
            in3 => \N__4051\,
            lcout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.REG_SPACE_3_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3654\,
            in1 => \N__3595\,
            in2 => \N__3526\,
            in3 => \N__3447\,
            lcout => \U409_ADDRESS_DECODE.REG_SPACE_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4046\,
            in1 => \N__4082\,
            in2 => \_gnd_net_\,
            in3 => \N__3994\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__3403\,
            in1 => \N__3855\,
            in2 => \N__3385\,
            in3 => \N__3955\,
            lcout => \CIA_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_1_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__4083\,
            in1 => \N__3856\,
            in2 => \_gnd_net_\,
            in3 => \N__4047\,
            lcout => \U409_ADDRESS_DECODE_ROMEN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.REG_SPACE_2_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__4423\,
            in1 => \N__4013\,
            in2 => \_gnd_net_\,
            in3 => \N__3920\,
            lcout => \U409_ADDRESS_DECODE.REG_SPACEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011111111"
        )
    port map (
            in0 => \N__3778\,
            in1 => \N__3792\,
            in2 => \N__3811\,
            in3 => \N__3853\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000100010"
        )
    port map (
            in0 => \N__3852\,
            in1 => \N__3807\,
            in2 => \N__3793\,
            in3 => \N__3777\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__3769\,
            in1 => \N__5402\,
            in2 => \_gnd_net_\,
            in3 => \N__6803\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4830\,
            in1 => \N__5251\,
            in2 => \N__4788\,
            in3 => \N__5150\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4668\,
            in1 => \N__5215\,
            in2 => \N__3739\,
            in3 => \N__5317\,
            lcout => \U409_TRANSFER_ACK.N_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4612\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC_net\,
            ce => \N__3736\,
            sr => \N__4747\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_sbtinv_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4267\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_RNIIFHQ_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4276\,
            in1 => \N__4255\,
            in2 => \N__4294\,
            in3 => \N__4095\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER6\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111011101"
        )
    port map (
            in0 => \N__4180\,
            in1 => \N__4159\,
            in2 => \N__4249\,
            in3 => \N__4204\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__6212\,
            in1 => \_gnd_net_\,
            in2 => \N__4246\,
            in3 => \N__4205\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001100"
        )
    port map (
            in0 => \N__4182\,
            in1 => \N__6208\,
            in2 => \N__4165\,
            in3 => \N__4140\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__4160\,
            in1 => \_gnd_net_\,
            in2 => \N__6225\,
            in3 => \N__4181\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111101110"
        )
    port map (
            in0 => \N__5163\,
            in1 => \N__5305\,
            in2 => \_gnd_net_\,
            in3 => \N__5269\,
            lcout => \U409_TRANSFER_ACK.N_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000001110001"
        )
    port map (
            in0 => \N__4183\,
            in1 => \N__4161\,
            in2 => \N__6353\,
            in3 => \N__4141\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            ce => 'H',
            sr => \N__6451\
        );

    \U409_TRANSFER_ACK.ROMENn_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__4107\,
            in1 => \N__5125\,
            in2 => \_gnd_net_\,
            in3 => \N__4129\,
            lcout => \ROMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            ce => 'H',
            sr => \N__6451\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010100100000"
        )
    port map (
            in0 => \N__4576\,
            in1 => \N__5629\,
            in2 => \N__5701\,
            in3 => \N__4096\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            ce => 'H',
            sr => \N__6451\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011010000"
        )
    port map (
            in0 => \N__5161\,
            in1 => \N__5219\,
            in2 => \N__5274\,
            in3 => \N__5319\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__6434\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111100000010"
        )
    port map (
            in0 => \N__4585\,
            in1 => \N__5320\,
            in2 => \N__5224\,
            in3 => \N__4290\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__6434\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101110100000"
        )
    port map (
            in0 => \N__5318\,
            in1 => \N__5264\,
            in2 => \N__5223\,
            in3 => \N__5160\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__6434\
        );

    \RESETn_ibuf_RNIM9SF_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6226\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4498\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC_net\,
            ce => \N__4480\,
            sr => \N__6446\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI8JGQ6_4_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4623\,
            in2 => \_gnd_net_\,
            in3 => \N__4642\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIEEVK7_0_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000010"
        )
    port map (
            in0 => \N__5541\,
            in1 => \N__4555\,
            in2 => \N__4261\,
            in3 => \N__4996\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4924\,
            in2 => \N__4258\,
            in3 => \N__4897\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__4746\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000110011"
        )
    port map (
            in0 => \N__4554\,
            in1 => \N__4997\,
            in2 => \N__5547\,
            in3 => \N__4624\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__4739\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5268\,
            in2 => \_gnd_net_\,
            in3 => \N__5162\,
            lcout => \U409_TRANSFER_ACK.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__5697\,
            in1 => \N__6475\,
            in2 => \N__5546\,
            in3 => \N__6505\,
            lcout => \U409_TRANSFER_ACK.N_142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__4532\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5496\,
            lcout => \U409_TRANSFER_ACK.N_35_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4497\,
            in1 => \N__4569\,
            in2 => \N__5542\,
            in3 => \N__4543\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNIBIO4C_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__4570\,
            in1 => \N__5527\,
            in2 => \N__4553\,
            in3 => \N__4496\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNO_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4483\,
            in3 => \N__6408\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__4321\,
            in1 => \N__4447\,
            in2 => \N__4829\,
            in3 => \N__4355\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__4811\,
            in1 => \N__4446\,
            in2 => \N__4362\,
            in3 => \N__4320\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CKM1_5_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4604\,
            in1 => \N__5026\,
            in2 => \N__5058\,
            in3 => \N__4890\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_4_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4994\,
            in1 => \N__4861\,
            in2 => \N__4645\,
            in3 => \N__4636\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__4961\,
            in1 => \N__4942\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_5_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5027\,
            in1 => \N__4603\,
            in2 => \N__5059\,
            in3 => \N__4860\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4635\,
            in1 => \N__4993\,
            in2 => \N__4627\,
            in3 => \N__4891\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__5057\,
            in1 => \N__4608\,
            in2 => \N__5089\,
            in3 => \N__5008\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__4721\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4840\,
            in1 => \N__5029\,
            in2 => \_gnd_net_\,
            in3 => \N__5073\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__4721\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__4998\,
            in1 => \_gnd_net_\,
            in2 => \N__5087\,
            in3 => \N__4945\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__4721\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__4944\,
            in1 => \N__4999\,
            in2 => \_gnd_net_\,
            in3 => \N__4963\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__4721\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__4922\,
            in1 => \N__4898\,
            in2 => \N__5088\,
            in3 => \N__4864\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__4721\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5007\,
            in2 => \N__5086\,
            in3 => \N__5056\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__4721\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4899\,
            in1 => \N__5028\,
            in2 => \N__4923\,
            in3 => \N__4862\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4995\,
            in1 => \N__4962\,
            in2 => \_gnd_net_\,
            in3 => \N__4943\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__4900\,
            in1 => \_gnd_net_\,
            in2 => \N__4867\,
            in3 => \N__4863\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5214\,
            in1 => \N__4834\,
            in2 => \N__4792\,
            in3 => \N__5273\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__5409\,
            in1 => \N__5427\,
            in2 => \N__6232\,
            in3 => \N__4765\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__5202\,
            in1 => \N__4684\,
            in2 => \N__4675\,
            in3 => \N__4654\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__6442\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5201\,
            in2 => \_gnd_net_\,
            in3 => \N__5304\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__6442\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5111\,
            in1 => \N__5962\,
            in2 => \_gnd_net_\,
            in3 => \N__5362\,
            lcout => \U409_TICK.TICK603_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5112\,
            in2 => \_gnd_net_\,
            in3 => \N__6038\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6878\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__5840\,
            in1 => \N__5801\,
            in2 => \N__5116\,
            in3 => \N__5767\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6878\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__5303\,
            in1 => \N__5275\,
            in2 => \N__5213\,
            in3 => \N__5167\,
            lcout => \U409_TRANSFER_ACK.N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5766\,
            in1 => \N__5841\,
            in2 => \N__5808\,
            in3 => \N__5341\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6878\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5110\,
            in2 => \N__6039\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6051\,
            in2 => \_gnd_net_\,
            in3 => \N__5095\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__6881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5982\,
            in2 => \_gnd_net_\,
            in3 => \N__5092\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__6881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5961\,
            in2 => \_gnd_net_\,
            in3 => \N__5365\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5361\,
            in2 => \_gnd_net_\,
            in3 => \N__5350\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__6881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5934\,
            in2 => \_gnd_net_\,
            in3 => \N__5347\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5874\,
            in2 => \_gnd_net_\,
            in3 => \N__5344\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__6881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5949\,
            in2 => \_gnd_net_\,
            in3 => \N__5335\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5712\,
            in2 => \_gnd_net_\,
            in3 => \N__5332\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5889\,
            in2 => \_gnd_net_\,
            in3 => \N__5329\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__6884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6003\,
            in2 => \_gnd_net_\,
            in3 => \N__5326\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__6884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6063\,
            in2 => \_gnd_net_\,
            in3 => \N__5323\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__6884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5902\,
            in2 => \_gnd_net_\,
            in3 => \N__5440\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__6884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5913\,
            in2 => \_gnd_net_\,
            in3 => \N__5437\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5853\,
            in2 => \_gnd_net_\,
            in3 => \N__5434\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6016\,
            in2 => \_gnd_net_\,
            in3 => \N__5431\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_DATA_BUFFERS.un1_BUFENn_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5428\,
            in1 => \N__6333\,
            in2 => \_gnd_net_\,
            in3 => \N__5410\,
            lcout => \BUFENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5577\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            ce => 'H',
            sr => \N__6450\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6775\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6186\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            ce => 'H',
            sr => \N__6450\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000011111"
        )
    port map (
            in0 => \N__5575\,
            in1 => \N__5598\,
            in2 => \N__5696\,
            in3 => \N__5635\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.i6_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110000001000"
        )
    port map (
            in0 => \N__5621\,
            in1 => \N__6188\,
            in2 => \N__5368\,
            in3 => \N__5689\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000011111"
        )
    port map (
            in0 => \N__5599\,
            in1 => \N__5576\,
            in2 => \N__5625\,
            in3 => \N__5452\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110000001000"
        )
    port map (
            in0 => \N__5688\,
            in1 => \N__6187\,
            in2 => \N__5665\,
            in3 => \N__5554\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__5765\,
            in1 => \N__5646\,
            in2 => \N__5809\,
            in3 => \N__5842\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6580\,
            in2 => \_gnd_net_\,
            in3 => \N__6558\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6470\,
            in2 => \_gnd_net_\,
            in3 => \N__6500\,
            lcout => \U409_TRANSFER_ACK.N_4\,
            ltout => \U409_TRANSFER_ACK.N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m4_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111000001010"
        )
    port map (
            in0 => \N__5617\,
            in1 => \N__5597\,
            in2 => \N__5581\,
            in3 => \N__5578\,
            lcout => \U409_TRANSFER_ACK.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_1_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5534\,
            in1 => \N__6471\,
            in2 => \_gnd_net_\,
            in3 => \N__6501\,
            lcout => \U409_TRANSFER_ACK.m8_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5837\,
            in1 => \N__5798\,
            in2 => \N__5769\,
            in3 => \N__5446\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6877\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6941\,
            in1 => \N__6982\,
            in2 => \N__7033\,
            in3 => \N__6619\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6877\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6064\,
            in1 => \N__6052\,
            in2 => \N__6040\,
            in3 => \N__6015\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6004\,
            in1 => \N__5992\,
            in2 => \N__5986\,
            in3 => \N__5983\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5836\,
            in1 => \N__5770\,
            in2 => \N__5971\,
            in3 => \N__5968\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6877\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5713\,
            in1 => \N__5950\,
            in2 => \N__5938\,
            in3 => \N__5914\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5758\,
            in1 => \N__5797\,
            in2 => \N__5923\,
            in3 => \N__5920\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6877\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__5901\,
            in1 => \N__5890\,
            in2 => \N__5878\,
            in3 => \N__5854\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => \U409_TICK.TICK603_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5838\,
            in1 => \N__5799\,
            in2 => \N__5863\,
            in3 => \N__5860\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5839\,
            in1 => \N__5800\,
            in2 => \N__5768\,
            in3 => \N__5719\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7166\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__6441\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6499\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__6441\
        );

    \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__6360\,
            in1 => \N__6334\,
            in2 => \_gnd_net_\,
            in3 => \N__6810\,
            lcout => \TCIn_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__6280\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6115\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS1n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNI692L_0_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6185\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6774\,
            lcout => \CIA_ENABLE\,
            ltout => \CIA_ENABLE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__6109\,
            in1 => \_gnd_net_\,
            in2 => \N__6091\,
            in3 => \_gnd_net_\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS0n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6975\,
            in1 => \N__6946\,
            in2 => \N__7030\,
            in3 => \N__6661\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6835\,
            in1 => \N__6538\,
            in2 => \N__6697\,
            in3 => \N__6557\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6610\,
            in1 => \N__6589\,
            in2 => \N__6067\,
            in3 => \N__6649\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__6736\,
            in1 => \N__6976\,
            in2 => \N__6592\,
            in3 => \N__7018\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__6748\,
            in1 => \N__6523\,
            in2 => \_gnd_net_\,
            in3 => \N__6578\,
            lcout => \U409_TICK.TICK503_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6631\,
            in1 => \N__6724\,
            in2 => \N__6679\,
            in3 => \N__7092\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__7014\,
            in1 => \N__6945\,
            in2 => \N__6583\,
            in3 => \N__6579\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__6944\,
            in1 => \N__6977\,
            in2 => \N__6712\,
            in3 => \N__7019\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6577\,
            in2 => \N__6559\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6537\,
            in2 => \_gnd_net_\,
            in3 => \N__6526\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__6882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6522\,
            in2 => \_gnd_net_\,
            in3 => \N__6511\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__6882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7059\,
            in2 => \_gnd_net_\,
            in3 => \N__6508\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__6882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6747\,
            in2 => \_gnd_net_\,
            in3 => \N__6727\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6723\,
            in2 => \_gnd_net_\,
            in3 => \N__6703\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7044\,
            in2 => \_gnd_net_\,
            in3 => \N__6700\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__6882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6693\,
            in2 => \_gnd_net_\,
            in3 => \N__6682\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__6882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6678\,
            in2 => \_gnd_net_\,
            in3 => \N__6652\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6645\,
            in2 => \_gnd_net_\,
            in3 => \N__6634\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__6885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6630\,
            in2 => \_gnd_net_\,
            in3 => \N__6613\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6606\,
            in2 => \_gnd_net_\,
            in3 => \N__6595\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__6885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7096\,
            in3 => \N__6847\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7071\,
            in2 => \_gnd_net_\,
            in3 => \N__6844\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6897\,
            in2 => \_gnd_net_\,
            in3 => \N__6841\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6834\,
            in2 => \_gnd_net_\,
            in3 => \N__6838\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_0_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7455\,
            in1 => \N__7414\,
            in2 => \N__7330\,
            in3 => \N__7431\,
            lcout => OPEN,
            ltout => \U409_CIA.CLK_CIA6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001101010101010"
        )
    port map (
            in0 => \N__7165\,
            in1 => \N__7213\,
            in2 => \N__6820\,
            in3 => \N__7144\,
            lcout => \CLK_CIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_1_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__7271\,
            in1 => \N__7295\,
            in2 => \N__7218\,
            in3 => \N__7413\,
            lcout => OPEN,
            ltout => \U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__7325\,
            in1 => \N__7346\,
            in2 => \N__6817\,
            in3 => \N__7242\,
            lcout => OPEN,
            ltout => \U409_CIA.VMA_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__6814\,
            in1 => \N__6764\,
            in2 => \N__6778\,
            in3 => \N__7326\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7430\,
            in2 => \_gnd_net_\,
            in3 => \N__7454\,
            lcout => \U409_CIA.CLK_CIA6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_1_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000010000"
        )
    port map (
            in0 => \N__7296\,
            in1 => \N__7243\,
            in2 => \N__7170\,
            in3 => \N__7272\,
            lcout => \U409_CIA.CLK_CIA_r_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__6939\,
            in1 => \N__6979\,
            in2 => \N__7031\,
            in3 => \N__7122\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__6978\,
            in1 => \N__6940\,
            in2 => \N__7111\,
            in3 => \N__7023\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6980\,
            in1 => \N__6942\,
            in2 => \N__7032\,
            in3 => \N__7078\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7072\,
            in1 => \N__7060\,
            in2 => \N__7048\,
            in3 => \N__6898\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6981\,
            in1 => \N__6943\,
            in2 => \N__6907\,
            in3 => \N__6904\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__7348\,
            in1 => \N__7369\,
            in2 => \N__7363\,
            in3 => \N__7192\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7273\,
            in1 => \N__7297\,
            in2 => \N__7219\,
            in3 => \N__7415\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__7324\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7416\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7241\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7323\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_2\,
            ltout => \U409_CIA.CIA_CLK_COUNT11_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__7359\,
            in1 => \N__7347\,
            in2 => \N__7333\,
            in3 => \N__7252\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7322\,
            in2 => \N__7417\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7294\,
            in2 => \_gnd_net_\,
            in3 => \N__7276\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__7382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7270\,
            in2 => \_gnd_net_\,
            in3 => \N__7246\,
            lcout => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7240\,
            in2 => \_gnd_net_\,
            in3 => \N__7222\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__7382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7214\,
            in2 => \_gnd_net_\,
            in3 => \N__7186\,
            lcout => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_6_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7456\,
            in2 => \_gnd_net_\,
            in3 => \N__7438\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\,
            clk => \N__7382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_7_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7432\,
            in2 => \_gnd_net_\,
            in3 => \N__7435\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7412\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7382\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 19 2024 10:38:08

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RAMENn : out std_logic;
    RASn : out std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__9952\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_OUT_i_i\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \N_888_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_451_cascade_\ : std_logic;
signal \N_48_i\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \U712_BYTE_ENABLE.N_352_cascade_\ : std_logic;
signal \N_49_i\ : std_logic;
signal \CLK40_OUT_i_i\ : std_logic;
signal \A_c_1\ : std_logic;
signal \U712_BYTE_ENABLE.N_457\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\ : std_logic;
signal \CLK40_OUT_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_BYTE_ENABLE.N_455\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_459_cascade_\ : std_logic;
signal \U712_BYTE_ENABLE.N_352\ : std_logic;
signal \N_47_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.N_362_i_0_en_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_362_i_0_en_0\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_7_cascade_\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_ac0_7_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \DRDDIR_i_0\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \U712_REG_SM.N_343_cascade_\ : std_logic;
signal \U712_REG_SM.N_358_cascade_\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_CHIP_RAM.N_563_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_215_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_565\ : std_logic;
signal \U712_CHIP_RAM.N_565_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_563\ : std_logic;
signal \U712_CHIP_RAM.N_445_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_a3_2_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_333_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_564\ : std_logic;
signal \U712_CHIP_RAM.N_471_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0_cascade_\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.N_447_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_333\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_330_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CHIP_RAM.N_554_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.N_332_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_493\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_351\ : std_logic;
signal \U712_CHIP_RAM.N_351_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_o2_1\ : std_logic;
signal \U712_CHIP_RAM.N_402\ : std_logic;
signal \U712_CHIP_RAM.N_341\ : std_logic;
signal \U712_CHIP_RAM.N_341_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_560\ : std_logic;
signal \U712_CHIP_RAM.N_450_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_326_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_326\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_CHIP_RAM.N_450\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_450_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_7\ : std_logic;
signal \U712_REG_SM.N_338\ : std_logic;
signal \U712_REG_SM.N_338_cascade_\ : std_logic;
signal \U712_REG_SM.N_354_cascade_\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \U712_REG_SM.N_431\ : std_logic;
signal \U712_REG_SM.N_358\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_71\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.N_369\ : std_logic;
signal \U712_CHIP_RAM.N_445\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_492\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_tz_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_331\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\ : std_logic;
signal \U712_CHIP_RAM.N_222\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_332\ : std_logic;
signal \U712_CHIP_RAM.N_346\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_0_i_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_4_0\ : std_logic;
signal \U712_CHIP_RAM.N_330\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_5_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_0_i_a3_0_1_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_2_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_2\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_3\ : std_logic;
signal \U712_CHIP_RAM.N_52\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.N_361\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_0\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_1\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_347_cascade_\ : std_logic;
signal \U712_REG_SM.N_559\ : std_logic;
signal \U712_REG_SM.N_559_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_GOZ0\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1\ : std_logic;
signal \U712_REG_SM.N_186_0\ : std_logic;
signal \U712_REG_SM.N_348_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.N_364_cascade_\ : std_logic;
signal \U712_REG_SM.N_343\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_2\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_370\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_368\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_2\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.N_374\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_2\ : std_logic;
signal \U712_BYTE_ENABLE.N_453\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_451\ : std_logic;
signal \N_50_i\ : std_logic;
signal \U712_REG_SM.N_354\ : std_logic;
signal \U712_REG_SM.N_394\ : std_logic;
signal \U712_REG_SM.N_364\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_5\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \A_c_0\ : std_logic;
signal \U712_REG_SM.N_395\ : std_logic;
signal \U712_REG_SM.LDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_LDSn_i\ : std_logic;
signal \U712_REG_SM.N_348\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_347\ : std_logic;
signal \U712_REG_SM.N_433\ : std_logic;
signal \U712_REG_SM.UDS_OUTZ0\ : std_logic;
signal \U712_REG_SM.DS_ENZ0\ : std_logic;
signal \U712_REG_SM_un1_UDSn_i\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \RnW_c\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U712_REG_SM.LDS_OUT_2_0_a3_0_a3Z0Z_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_8\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.N_367_cascade_\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \A_c_14\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.N_371\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_6\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\ : std_logic;
signal \CASn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.N_373\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.N_372\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i_0\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    CLK_EN <= \CLK_EN_wire\;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    LDSn <= \LDSn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_OUT_i\,
            REFERENCECLK => \N__3540\,
            RESETB => \N__5061\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_OUT\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9952\,
            DIN => \N__9951\,
            DOUT => \N__9950\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9952\,
            PADOUT => \N__9951\,
            PADIN => \N__9950\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4740\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9943\,
            DIN => \N__9942\,
            DOUT => \N__9941\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9943\,
            PADOUT => \N__9942\,
            PADIN => \N__9941\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9934\,
            DIN => \N__9933\,
            DOUT => \N__9932\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9934\,
            PADOUT => \N__9933\,
            PADIN => \N__9932\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7890\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9925\,
            DIN => \N__9924\,
            DOUT => \N__9923\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9925\,
            PADOUT => \N__9924\,
            PADIN => \N__9923\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4074\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9916\,
            DIN => \N__9915\,
            DOUT => \N__9914\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9916\,
            PADOUT => \N__9915\,
            PADIN => \N__9914\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9907\,
            DIN => \N__9906\,
            DOUT => \N__9905\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9907\,
            PADOUT => \N__9906\,
            PADIN => \N__9905\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9898\,
            DIN => \N__9897\,
            DOUT => \N__9896\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9898\,
            PADOUT => \N__9897\,
            PADIN => \N__9896\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9889\,
            DIN => \N__9888\,
            DOUT => \N__9887\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9889\,
            PADOUT => \N__9888\,
            PADIN => \N__9887\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9880\,
            DIN => \N__9879\,
            DOUT => \N__9878\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9880\,
            PADOUT => \N__9879\,
            PADIN => \N__9878\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9871\,
            DIN => \N__9870\,
            DOUT => \N__9869\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9871\,
            PADOUT => \N__9870\,
            PADIN => \N__9869\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9862\,
            DIN => \N__9861\,
            DOUT => \N__9860\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9862\,
            PADOUT => \N__9861\,
            PADIN => \N__9860\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6594\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9853\,
            DIN => \N__9852\,
            DOUT => \N__9851\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9853\,
            PADOUT => \N__9852\,
            PADIN => \N__9851\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5330\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9844\,
            DIN => \N__9843\,
            DOUT => \N__9842\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9844\,
            PADOUT => \N__9843\,
            PADIN => \N__9842\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9835\,
            DIN => \N__9834\,
            DOUT => \N__9833\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9835\,
            PADOUT => \N__9834\,
            PADIN => \N__9833\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9826\,
            DIN => \N__9825\,
            DOUT => \N__9824\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9826\,
            PADOUT => \N__9825\,
            PADIN => \N__9824\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3948\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9817\,
            DIN => \N__9816\,
            DOUT => \N__9815\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9817\,
            PADOUT => \N__9816\,
            PADIN => \N__9815\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9808\,
            DIN => \N__9807\,
            DOUT => \N__9806\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9808\,
            PADOUT => \N__9807\,
            PADIN => \N__9806\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9799\,
            DIN => \N__9798\,
            DOUT => \N__9797\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9799\,
            PADOUT => \N__9798\,
            PADIN => \N__9797\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7173\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9790\,
            DIN => \N__9789\,
            DOUT => \N__9788\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9790\,
            PADOUT => \N__9789\,
            PADIN => \N__9788\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9781\,
            DIN => \N__9780\,
            DOUT => \N__9779\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9781\,
            PADOUT => \N__9780\,
            PADIN => \N__9779\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7812\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9772\,
            DIN => \N__9771\,
            DOUT => \N__9770\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9772\,
            PADOUT => \N__9771\,
            PADIN => \N__9770\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9763\,
            DIN => \N__9762\,
            DOUT => \N__9761\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9763\,
            PADOUT => \N__9762\,
            PADIN => \N__9761\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9754\,
            DIN => \N__9753\,
            DOUT => \N__9752\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9754\,
            PADOUT => \N__9753\,
            PADIN => \N__9752\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9745\,
            DIN => \N__9744\,
            DOUT => \N__9743\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9745\,
            PADOUT => \N__9744\,
            PADIN => \N__9743\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9736\,
            DIN => \N__9735\,
            DOUT => \N__9734\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9736\,
            PADOUT => \N__9735\,
            PADIN => \N__9734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9727\,
            DIN => \N__9726\,
            DOUT => \N__9725\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9727\,
            PADOUT => \N__9726\,
            PADIN => \N__9725\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4446\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9718\,
            DIN => \N__9717\,
            DOUT => \N__9716\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9718\,
            PADOUT => \N__9717\,
            PADIN => \N__9716\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9709\,
            DIN => \N__9708\,
            DOUT => \N__9707\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9709\,
            PADOUT => \N__9708\,
            PADIN => \N__9707\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9700\,
            DIN => \N__9699\,
            DOUT => \N__9698\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9700\,
            PADOUT => \N__9699\,
            PADIN => \N__9698\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9691\,
            DIN => \N__9690\,
            DOUT => \N__9689\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9691\,
            PADOUT => \N__9690\,
            PADIN => \N__9689\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9682\,
            DIN => \N__9681\,
            DOUT => \N__9680\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9682\,
            PADOUT => \N__9681\,
            PADIN => \N__9680\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9673\,
            DIN => \N__9672\,
            DOUT => \N__9671\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9673\,
            PADOUT => \N__9672\,
            PADIN => \N__9671\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7773\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9664\,
            DIN => \N__9663\,
            DOUT => \N__9662\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9664\,
            PADOUT => \N__9663\,
            PADIN => \N__9662\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9655\,
            DIN => \N__9654\,
            DOUT => \N__9653\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9655\,
            PADOUT => \N__9654\,
            PADIN => \N__9653\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9646\,
            DIN => \N__9645\,
            DOUT => \N__9644\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9646\,
            PADOUT => \N__9645\,
            PADIN => \N__9644\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9637\,
            DIN => \N__9636\,
            DOUT => \N__9635\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9637\,
            PADOUT => \N__9636\,
            PADIN => \N__9635\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9628\,
            DIN => \N__9627\,
            DOUT => \N__9626\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9628\,
            PADOUT => \N__9627\,
            PADIN => \N__9626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3675\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9619\,
            DIN => \N__9618\,
            DOUT => \N__9617\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9619\,
            PADOUT => \N__9618\,
            PADIN => \N__9617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6825\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9610\,
            DIN => \N__9609\,
            DOUT => \N__9608\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9610\,
            PADOUT => \N__9609\,
            PADIN => \N__9608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9601\,
            DIN => \N__9600\,
            DOUT => \N__9599\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9601\,
            PADOUT => \N__9600\,
            PADIN => \N__9599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7797\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9592\,
            DIN => \N__9591\,
            DOUT => \N__9590\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9592\,
            PADOUT => \N__9591\,
            PADIN => \N__9590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9583\,
            DIN => \N__9582\,
            DOUT => \N__9581\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9583\,
            PADOUT => \N__9582\,
            PADIN => \N__9581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9574\,
            DIN => \N__9573\,
            DOUT => \N__9572\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9574\,
            PADOUT => \N__9573\,
            PADIN => \N__9572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3564\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9565\,
            DIN => \N__9564\,
            DOUT => \N__9563\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9565\,
            PADOUT => \N__9564\,
            PADIN => \N__9563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9556\,
            DIN => \N__9555\,
            DOUT => \N__9554\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9556\,
            PADOUT => \N__9555\,
            PADIN => \N__9554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6213\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9547\,
            DIN => \N__9546\,
            DOUT => \N__9545\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9547\,
            PADOUT => \N__9546\,
            PADIN => \N__9545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6360\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9538\,
            DIN => \N__9537\,
            DOUT => \N__9536\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9538\,
            PADOUT => \N__9537\,
            PADIN => \N__9536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9529\,
            DIN => \N__9528\,
            DOUT => \N__9527\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9529\,
            PADOUT => \N__9528\,
            PADIN => \N__9527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9520\,
            DIN => \N__9519\,
            DOUT => \N__9518\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9520\,
            PADOUT => \N__9519\,
            PADIN => \N__9518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9511\,
            DIN => \N__9510\,
            DOUT => \N__9509\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9511\,
            PADOUT => \N__9510\,
            PADIN => \N__9509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7323\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9502\,
            DIN => \N__9501\,
            DOUT => \N__9500\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9502\,
            PADOUT => \N__9501\,
            PADIN => \N__9500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9493\,
            DIN => \N__9492\,
            DOUT => \N__9491\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9493\,
            PADOUT => \N__9492\,
            PADIN => \N__9491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7302\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9484\,
            DIN => \N__9483\,
            DOUT => \N__9482\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9484\,
            PADOUT => \N__9483\,
            PADIN => \N__9482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4245\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9475\,
            DIN => \N__9474\,
            DOUT => \N__9473\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9475\,
            PADOUT => \N__9474\,
            PADIN => \N__9473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4029\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9466\,
            DIN => \N__9465\,
            DOUT => \N__9464\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9466\,
            PADOUT => \N__9465\,
            PADIN => \N__9464\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6624\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9457\,
            DIN => \N__9456\,
            DOUT => \N__9455\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9457\,
            PADOUT => \N__9456\,
            PADIN => \N__9455\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6212\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9448\,
            DIN => \N__9447\,
            DOUT => \N__9446\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9448\,
            PADOUT => \N__9447\,
            PADIN => \N__9446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9439\,
            DIN => \N__9438\,
            DOUT => \N__9437\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9439\,
            PADOUT => \N__9438\,
            PADIN => \N__9437\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9430\,
            DIN => \N__9429\,
            DOUT => \N__9428\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9430\,
            PADOUT => \N__9429\,
            PADIN => \N__9428\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3588\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9421\,
            DIN => \N__9420\,
            DOUT => \N__9419\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9421\,
            PADOUT => \N__9420\,
            PADIN => \N__9419\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7872\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9412\,
            DIN => \N__9411\,
            DOUT => \N__9410\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9412\,
            PADOUT => \N__9411\,
            PADIN => \N__9410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4107\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9403\,
            DIN => \N__9402\,
            DOUT => \N__9401\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9403\,
            PADOUT => \N__9402\,
            PADIN => \N__9401\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3699\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9394\,
            DIN => \N__9393\,
            DOUT => \N__9392\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9394\,
            PADOUT => \N__9393\,
            PADIN => \N__9392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9385\,
            DIN => \N__9384\,
            DOUT => \N__9383\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9385\,
            PADOUT => \N__9384\,
            PADIN => \N__9383\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9376\,
            DIN => \N__9375\,
            DOUT => \N__9374\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9376\,
            PADOUT => \N__9375\,
            PADIN => \N__9374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9367\,
            DIN => \N__9366\,
            DOUT => \N__9365\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9367\,
            PADOUT => \N__9366\,
            PADIN => \N__9365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9358\,
            DIN => \N__9357\,
            DOUT => \N__9356\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9358\,
            PADOUT => \N__9357\,
            PADIN => \N__9356\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6336\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9349\,
            DIN => \N__9348\,
            DOUT => \N__9347\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9349\,
            PADOUT => \N__9348\,
            PADIN => \N__9347\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9340\,
            DIN => \N__9339\,
            DOUT => \N__9338\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9340\,
            PADOUT => \N__9339\,
            PADIN => \N__9338\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7023\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9331\,
            DIN => \N__9330\,
            DOUT => \N__9329\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9331\,
            PADOUT => \N__9330\,
            PADIN => \N__9329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3606\,
            DIN0 => OPEN,
            DOUT0 => \N__3837\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9322\,
            DIN => \N__9321\,
            DOUT => \N__9320\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9322\,
            PADOUT => \N__9321\,
            PADIN => \N__9320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5070\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9313\,
            DIN => \N__9312\,
            DOUT => \N__9311\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9313\,
            PADOUT => \N__9312\,
            PADIN => \N__9311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9304\,
            DIN => \N__9303\,
            DOUT => \N__9302\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9304\,
            PADOUT => \N__9303\,
            PADIN => \N__9302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9295\,
            DIN => \N__9294\,
            DOUT => \N__9293\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9295\,
            PADOUT => \N__9294\,
            PADIN => \N__9293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7245\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9286\,
            DIN => \N__9285\,
            DOUT => \N__9284\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9286\,
            PADOUT => \N__9285\,
            PADIN => \N__9284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9277\,
            DIN => \N__9276\,
            DOUT => \N__9275\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9277\,
            PADOUT => \N__9276\,
            PADIN => \N__9275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9268\,
            DIN => \N__9267\,
            DOUT => \N__9266\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9268\,
            PADOUT => \N__9267\,
            PADIN => \N__9266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9259\,
            DIN => \N__9258\,
            DOUT => \N__9257\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9259\,
            PADOUT => \N__9258\,
            PADIN => \N__9257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9250\,
            DIN => \N__9249\,
            DOUT => \N__9248\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9250\,
            PADOUT => \N__9249\,
            PADIN => \N__9248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8490\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9241\,
            DIN => \N__9240\,
            DOUT => \N__9239\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9241\,
            PADOUT => \N__9240\,
            PADIN => \N__9239\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7548\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2198\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9218\
        );

    \I__2197\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9215\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__9218\,
            I => \N__9212\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__9215\,
            I => \N__9209\
        );

    \I__2194\ : Span4Mux_v
    port map (
            O => \N__9212\,
            I => \N__9206\
        );

    \I__2193\ : Span12Mux_v
    port map (
            O => \N__9209\,
            I => \N__9203\
        );

    \I__2192\ : Span4Mux_h
    port map (
            O => \N__9206\,
            I => \N__9200\
        );

    \I__2191\ : Span12Mux_h
    port map (
            O => \N__9203\,
            I => \N__9197\
        );

    \I__2190\ : Span4Mux_h
    port map (
            O => \N__9200\,
            I => \N__9194\
        );

    \I__2189\ : Odrv12
    port map (
            O => \N__9197\,
            I => \RAS0n_c\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__9194\,
            I => \RAS0n_c\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9189\,
            I => \N__9186\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9186\,
            I => \N__9183\
        );

    \I__2185\ : Span4Mux_v
    port map (
            O => \N__9183\,
            I => \N__9180\
        );

    \I__2184\ : Sp12to4
    port map (
            O => \N__9180\,
            I => \N__9177\
        );

    \I__2183\ : Odrv12
    port map (
            O => \N__9177\,
            I => \RAS1n_c\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9174\,
            I => \N__9170\
        );

    \I__2181\ : InMux
    port map (
            O => \N__9173\,
            I => \N__9167\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__9170\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9167\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2178\ : InMux
    port map (
            O => \N__9162\,
            I => \N__9159\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__9159\,
            I => \N__9142\
        );

    \I__2176\ : ClkMux
    port map (
            O => \N__9158\,
            I => \N__9030\
        );

    \I__2175\ : ClkMux
    port map (
            O => \N__9157\,
            I => \N__9030\
        );

    \I__2174\ : ClkMux
    port map (
            O => \N__9156\,
            I => \N__9030\
        );

    \I__2173\ : ClkMux
    port map (
            O => \N__9155\,
            I => \N__9030\
        );

    \I__2172\ : ClkMux
    port map (
            O => \N__9154\,
            I => \N__9030\
        );

    \I__2171\ : ClkMux
    port map (
            O => \N__9153\,
            I => \N__9030\
        );

    \I__2170\ : ClkMux
    port map (
            O => \N__9152\,
            I => \N__9030\
        );

    \I__2169\ : ClkMux
    port map (
            O => \N__9151\,
            I => \N__9030\
        );

    \I__2168\ : ClkMux
    port map (
            O => \N__9150\,
            I => \N__9030\
        );

    \I__2167\ : ClkMux
    port map (
            O => \N__9149\,
            I => \N__9030\
        );

    \I__2166\ : ClkMux
    port map (
            O => \N__9148\,
            I => \N__9030\
        );

    \I__2165\ : ClkMux
    port map (
            O => \N__9147\,
            I => \N__9030\
        );

    \I__2164\ : ClkMux
    port map (
            O => \N__9146\,
            I => \N__9030\
        );

    \I__2163\ : ClkMux
    port map (
            O => \N__9145\,
            I => \N__9030\
        );

    \I__2162\ : Glb2LocalMux
    port map (
            O => \N__9142\,
            I => \N__9030\
        );

    \I__2161\ : ClkMux
    port map (
            O => \N__9141\,
            I => \N__9030\
        );

    \I__2160\ : ClkMux
    port map (
            O => \N__9140\,
            I => \N__9030\
        );

    \I__2159\ : ClkMux
    port map (
            O => \N__9139\,
            I => \N__9030\
        );

    \I__2158\ : ClkMux
    port map (
            O => \N__9138\,
            I => \N__9030\
        );

    \I__2157\ : ClkMux
    port map (
            O => \N__9137\,
            I => \N__9030\
        );

    \I__2156\ : ClkMux
    port map (
            O => \N__9136\,
            I => \N__9030\
        );

    \I__2155\ : ClkMux
    port map (
            O => \N__9135\,
            I => \N__9030\
        );

    \I__2154\ : ClkMux
    port map (
            O => \N__9134\,
            I => \N__9030\
        );

    \I__2153\ : ClkMux
    port map (
            O => \N__9133\,
            I => \N__9030\
        );

    \I__2152\ : ClkMux
    port map (
            O => \N__9132\,
            I => \N__9030\
        );

    \I__2151\ : ClkMux
    port map (
            O => \N__9131\,
            I => \N__9030\
        );

    \I__2150\ : ClkMux
    port map (
            O => \N__9130\,
            I => \N__9030\
        );

    \I__2149\ : ClkMux
    port map (
            O => \N__9129\,
            I => \N__9030\
        );

    \I__2148\ : ClkMux
    port map (
            O => \N__9128\,
            I => \N__9030\
        );

    \I__2147\ : ClkMux
    port map (
            O => \N__9127\,
            I => \N__9030\
        );

    \I__2146\ : ClkMux
    port map (
            O => \N__9126\,
            I => \N__9030\
        );

    \I__2145\ : ClkMux
    port map (
            O => \N__9125\,
            I => \N__9030\
        );

    \I__2144\ : ClkMux
    port map (
            O => \N__9124\,
            I => \N__9030\
        );

    \I__2143\ : ClkMux
    port map (
            O => \N__9123\,
            I => \N__9030\
        );

    \I__2142\ : ClkMux
    port map (
            O => \N__9122\,
            I => \N__9030\
        );

    \I__2141\ : ClkMux
    port map (
            O => \N__9121\,
            I => \N__9030\
        );

    \I__2140\ : ClkMux
    port map (
            O => \N__9120\,
            I => \N__9030\
        );

    \I__2139\ : ClkMux
    port map (
            O => \N__9119\,
            I => \N__9030\
        );

    \I__2138\ : ClkMux
    port map (
            O => \N__9118\,
            I => \N__9030\
        );

    \I__2137\ : ClkMux
    port map (
            O => \N__9117\,
            I => \N__9030\
        );

    \I__2136\ : ClkMux
    port map (
            O => \N__9116\,
            I => \N__9030\
        );

    \I__2135\ : ClkMux
    port map (
            O => \N__9115\,
            I => \N__9030\
        );

    \I__2134\ : GlobalMux
    port map (
            O => \N__9030\,
            I => \CLK80_OUT\
        );

    \I__2133\ : InMux
    port map (
            O => \N__9027\,
            I => \N__9013\
        );

    \I__2132\ : InMux
    port map (
            O => \N__9026\,
            I => \N__9010\
        );

    \I__2131\ : InMux
    port map (
            O => \N__9025\,
            I => \N__9007\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9024\,
            I => \N__9000\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9023\,
            I => \N__9000\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9022\,
            I => \N__9000\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9021\,
            I => \N__8997\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9020\,
            I => \N__8994\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9019\,
            I => \N__8991\
        );

    \I__2124\ : InMux
    port map (
            O => \N__9018\,
            I => \N__8988\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9017\,
            I => \N__8983\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9016\,
            I => \N__8983\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__9013\,
            I => \N__8975\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9010\,
            I => \N__8969\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__9007\,
            I => \N__8961\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9000\,
            I => \N__8958\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__8997\,
            I => \N__8955\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__8994\,
            I => \N__8948\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__8991\,
            I => \N__8945\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__8988\,
            I => \N__8939\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__8983\,
            I => \N__8924\
        );

    \I__2112\ : SRMux
    port map (
            O => \N__8982\,
            I => \N__8832\
        );

    \I__2111\ : SRMux
    port map (
            O => \N__8981\,
            I => \N__8832\
        );

    \I__2110\ : SRMux
    port map (
            O => \N__8980\,
            I => \N__8832\
        );

    \I__2109\ : SRMux
    port map (
            O => \N__8979\,
            I => \N__8832\
        );

    \I__2108\ : SRMux
    port map (
            O => \N__8978\,
            I => \N__8832\
        );

    \I__2107\ : Glb2LocalMux
    port map (
            O => \N__8975\,
            I => \N__8832\
        );

    \I__2106\ : SRMux
    port map (
            O => \N__8974\,
            I => \N__8832\
        );

    \I__2105\ : SRMux
    port map (
            O => \N__8973\,
            I => \N__8832\
        );

    \I__2104\ : SRMux
    port map (
            O => \N__8972\,
            I => \N__8832\
        );

    \I__2103\ : Glb2LocalMux
    port map (
            O => \N__8969\,
            I => \N__8832\
        );

    \I__2102\ : SRMux
    port map (
            O => \N__8968\,
            I => \N__8832\
        );

    \I__2101\ : SRMux
    port map (
            O => \N__8967\,
            I => \N__8832\
        );

    \I__2100\ : SRMux
    port map (
            O => \N__8966\,
            I => \N__8832\
        );

    \I__2099\ : SRMux
    port map (
            O => \N__8965\,
            I => \N__8832\
        );

    \I__2098\ : SRMux
    port map (
            O => \N__8964\,
            I => \N__8832\
        );

    \I__2097\ : Glb2LocalMux
    port map (
            O => \N__8961\,
            I => \N__8832\
        );

    \I__2096\ : Glb2LocalMux
    port map (
            O => \N__8958\,
            I => \N__8832\
        );

    \I__2095\ : Glb2LocalMux
    port map (
            O => \N__8955\,
            I => \N__8832\
        );

    \I__2094\ : SRMux
    port map (
            O => \N__8954\,
            I => \N__8832\
        );

    \I__2093\ : SRMux
    port map (
            O => \N__8953\,
            I => \N__8832\
        );

    \I__2092\ : SRMux
    port map (
            O => \N__8952\,
            I => \N__8832\
        );

    \I__2091\ : SRMux
    port map (
            O => \N__8951\,
            I => \N__8832\
        );

    \I__2090\ : Glb2LocalMux
    port map (
            O => \N__8948\,
            I => \N__8832\
        );

    \I__2089\ : Glb2LocalMux
    port map (
            O => \N__8945\,
            I => \N__8832\
        );

    \I__2088\ : SRMux
    port map (
            O => \N__8944\,
            I => \N__8832\
        );

    \I__2087\ : SRMux
    port map (
            O => \N__8943\,
            I => \N__8832\
        );

    \I__2086\ : SRMux
    port map (
            O => \N__8942\,
            I => \N__8832\
        );

    \I__2085\ : Glb2LocalMux
    port map (
            O => \N__8939\,
            I => \N__8832\
        );

    \I__2084\ : SRMux
    port map (
            O => \N__8938\,
            I => \N__8832\
        );

    \I__2083\ : SRMux
    port map (
            O => \N__8937\,
            I => \N__8832\
        );

    \I__2082\ : SRMux
    port map (
            O => \N__8936\,
            I => \N__8832\
        );

    \I__2081\ : SRMux
    port map (
            O => \N__8935\,
            I => \N__8832\
        );

    \I__2080\ : SRMux
    port map (
            O => \N__8934\,
            I => \N__8832\
        );

    \I__2079\ : SRMux
    port map (
            O => \N__8933\,
            I => \N__8832\
        );

    \I__2078\ : SRMux
    port map (
            O => \N__8932\,
            I => \N__8832\
        );

    \I__2077\ : SRMux
    port map (
            O => \N__8931\,
            I => \N__8832\
        );

    \I__2076\ : SRMux
    port map (
            O => \N__8930\,
            I => \N__8832\
        );

    \I__2075\ : SRMux
    port map (
            O => \N__8929\,
            I => \N__8832\
        );

    \I__2074\ : SRMux
    port map (
            O => \N__8928\,
            I => \N__8832\
        );

    \I__2073\ : SRMux
    port map (
            O => \N__8927\,
            I => \N__8832\
        );

    \I__2072\ : Glb2LocalMux
    port map (
            O => \N__8924\,
            I => \N__8832\
        );

    \I__2071\ : SRMux
    port map (
            O => \N__8923\,
            I => \N__8832\
        );

    \I__2070\ : SRMux
    port map (
            O => \N__8922\,
            I => \N__8832\
        );

    \I__2069\ : SRMux
    port map (
            O => \N__8921\,
            I => \N__8832\
        );

    \I__2068\ : GlobalMux
    port map (
            O => \N__8832\,
            I => \N__8829\
        );

    \I__2067\ : gio2CtrlBuf
    port map (
            O => \N__8829\,
            I => \RESETn_c_i_g\
        );

    \I__2066\ : InMux
    port map (
            O => \N__8826\,
            I => \N__8823\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__8823\,
            I => \U712_CHIP_RAM.N_372\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__8820\,
            I => \N__8814\
        );

    \I__2063\ : InMux
    port map (
            O => \N__8819\,
            I => \N__8809\
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__8818\,
            I => \N__8806\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__8817\,
            I => \N__8803\
        );

    \I__2060\ : InMux
    port map (
            O => \N__8814\,
            I => \N__8797\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__8813\,
            I => \N__8794\
        );

    \I__2058\ : InMux
    port map (
            O => \N__8812\,
            I => \N__8791\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__8809\,
            I => \N__8785\
        );

    \I__2056\ : InMux
    port map (
            O => \N__8806\,
            I => \N__8782\
        );

    \I__2055\ : InMux
    port map (
            O => \N__8803\,
            I => \N__8779\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__8802\,
            I => \N__8776\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__8801\,
            I => \N__8773\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__8800\,
            I => \N__8770\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__8797\,
            I => \N__8765\
        );

    \I__2050\ : InMux
    port map (
            O => \N__8794\,
            I => \N__8762\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__8791\,
            I => \N__8759\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__8790\,
            I => \N__8755\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__8789\,
            I => \N__8752\
        );

    \I__2046\ : InMux
    port map (
            O => \N__8788\,
            I => \N__8749\
        );

    \I__2045\ : Span4Mux_v
    port map (
            O => \N__8785\,
            I => \N__8744\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__8782\,
            I => \N__8744\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__8779\,
            I => \N__8741\
        );

    \I__2042\ : InMux
    port map (
            O => \N__8776\,
            I => \N__8734\
        );

    \I__2041\ : InMux
    port map (
            O => \N__8773\,
            I => \N__8734\
        );

    \I__2040\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8734\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__8769\,
            I => \N__8730\
        );

    \I__2038\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8727\
        );

    \I__2037\ : Span4Mux_v
    port map (
            O => \N__8765\,
            I => \N__8724\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__8762\,
            I => \N__8719\
        );

    \I__2035\ : Span4Mux_h
    port map (
            O => \N__8759\,
            I => \N__8719\
        );

    \I__2034\ : InMux
    port map (
            O => \N__8758\,
            I => \N__8714\
        );

    \I__2033\ : InMux
    port map (
            O => \N__8755\,
            I => \N__8714\
        );

    \I__2032\ : InMux
    port map (
            O => \N__8752\,
            I => \N__8711\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__8749\,
            I => \N__8704\
        );

    \I__2030\ : Span4Mux_h
    port map (
            O => \N__8744\,
            I => \N__8704\
        );

    \I__2029\ : Span4Mux_h
    port map (
            O => \N__8741\,
            I => \N__8704\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__8734\,
            I => \N__8701\
        );

    \I__2027\ : InMux
    port map (
            O => \N__8733\,
            I => \N__8696\
        );

    \I__2026\ : InMux
    port map (
            O => \N__8730\,
            I => \N__8696\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__8727\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2024\ : Odrv4
    port map (
            O => \N__8724\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__8719\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__8714\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__8711\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__8704\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2019\ : Odrv12
    port map (
            O => \N__8701\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__8696\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2017\ : InMux
    port map (
            O => \N__8679\,
            I => \N__8666\
        );

    \I__2016\ : InMux
    port map (
            O => \N__8678\,
            I => \N__8666\
        );

    \I__2015\ : InMux
    port map (
            O => \N__8677\,
            I => \N__8661\
        );

    \I__2014\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8661\
        );

    \I__2013\ : CascadeMux
    port map (
            O => \N__8675\,
            I => \N__8658\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__8674\,
            I => \N__8655\
        );

    \I__2011\ : InMux
    port map (
            O => \N__8673\,
            I => \N__8651\
        );

    \I__2010\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8647\
        );

    \I__2009\ : InMux
    port map (
            O => \N__8671\,
            I => \N__8644\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__8666\,
            I => \N__8639\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__8661\,
            I => \N__8639\
        );

    \I__2006\ : InMux
    port map (
            O => \N__8658\,
            I => \N__8634\
        );

    \I__2005\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8634\
        );

    \I__2004\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8631\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__8651\,
            I => \N__8628\
        );

    \I__2002\ : InMux
    port map (
            O => \N__8650\,
            I => \N__8625\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__8647\,
            I => \N__8620\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__8644\,
            I => \N__8620\
        );

    \I__1999\ : Span4Mux_v
    port map (
            O => \N__8639\,
            I => \N__8615\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__8634\,
            I => \N__8615\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__8631\,
            I => \N__8610\
        );

    \I__1996\ : Span12Mux_s9_v
    port map (
            O => \N__8628\,
            I => \N__8607\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__8625\,
            I => \N__8600\
        );

    \I__1994\ : Span4Mux_v
    port map (
            O => \N__8620\,
            I => \N__8600\
        );

    \I__1993\ : Span4Mux_h
    port map (
            O => \N__8615\,
            I => \N__8600\
        );

    \I__1992\ : InMux
    port map (
            O => \N__8614\,
            I => \N__8597\
        );

    \I__1991\ : InMux
    port map (
            O => \N__8613\,
            I => \N__8594\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__8610\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__1989\ : Odrv12
    port map (
            O => \N__8607\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__8600\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__8597\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__8594\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__1985\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8573\
        );

    \I__1984\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8568\
        );

    \I__1983\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8568\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8580\,
            I => \N__8565\
        );

    \I__1981\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8560\
        );

    \I__1980\ : InMux
    port map (
            O => \N__8578\,
            I => \N__8560\
        );

    \I__1979\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8555\
        );

    \I__1978\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8552\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__8573\,
            I => \N__8549\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__8568\,
            I => \N__8546\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__8565\,
            I => \N__8543\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__8560\,
            I => \N__8540\
        );

    \I__1973\ : InMux
    port map (
            O => \N__8559\,
            I => \N__8531\
        );

    \I__1972\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8531\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__8555\,
            I => \N__8528\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__8552\,
            I => \N__8523\
        );

    \I__1969\ : Span4Mux_h
    port map (
            O => \N__8549\,
            I => \N__8523\
        );

    \I__1968\ : Span4Mux_h
    port map (
            O => \N__8546\,
            I => \N__8516\
        );

    \I__1967\ : Span4Mux_v
    port map (
            O => \N__8543\,
            I => \N__8516\
        );

    \I__1966\ : Span4Mux_v
    port map (
            O => \N__8540\,
            I => \N__8516\
        );

    \I__1965\ : InMux
    port map (
            O => \N__8539\,
            I => \N__8513\
        );

    \I__1964\ : InMux
    port map (
            O => \N__8538\,
            I => \N__8508\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8537\,
            I => \N__8508\
        );

    \I__1962\ : InMux
    port map (
            O => \N__8536\,
            I => \N__8505\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__8531\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1960\ : Odrv4
    port map (
            O => \N__8528\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__8523\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__8516\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__8513\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__8508\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__8505\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1954\ : IoInMux
    port map (
            O => \N__8490\,
            I => \N__8487\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__8487\,
            I => \N__8484\
        );

    \I__1952\ : Span12Mux_s1_h
    port map (
            O => \N__8484\,
            I => \N__8481\
        );

    \I__1951\ : Span12Mux_h
    port map (
            O => \N__8481\,
            I => \N__8478\
        );

    \I__1950\ : Odrv12
    port map (
            O => \N__8478\,
            I => \CMA_c_5\
        );

    \I__1949\ : CEMux
    port map (
            O => \N__8475\,
            I => \N__8471\
        );

    \I__1948\ : CEMux
    port map (
            O => \N__8474\,
            I => \N__8468\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__8471\,
            I => \N__8461\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__8468\,
            I => \N__8458\
        );

    \I__1945\ : CEMux
    port map (
            O => \N__8467\,
            I => \N__8455\
        );

    \I__1944\ : CEMux
    port map (
            O => \N__8466\,
            I => \N__8452\
        );

    \I__1943\ : CEMux
    port map (
            O => \N__8465\,
            I => \N__8449\
        );

    \I__1942\ : CEMux
    port map (
            O => \N__8464\,
            I => \N__8446\
        );

    \I__1941\ : Span4Mux_v
    port map (
            O => \N__8461\,
            I => \N__8441\
        );

    \I__1940\ : Span4Mux_h
    port map (
            O => \N__8458\,
            I => \N__8441\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__8455\,
            I => \N__8438\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__8452\,
            I => \N__8431\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__8449\,
            I => \N__8431\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8446\,
            I => \N__8431\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__8441\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1934\ : Odrv12
    port map (
            O => \N__8438\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1933\ : Odrv4
    port map (
            O => \N__8431\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8424\,
            I => \N__8420\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8417\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__8420\,
            I => \N__8414\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__8417\,
            I => \N__8411\
        );

    \I__1928\ : Sp12to4
    port map (
            O => \N__8414\,
            I => \N__8408\
        );

    \I__1927\ : Span12Mux_v
    port map (
            O => \N__8411\,
            I => \N__8405\
        );

    \I__1926\ : Span12Mux_v
    port map (
            O => \N__8408\,
            I => \N__8402\
        );

    \I__1925\ : Span12Mux_h
    port map (
            O => \N__8405\,
            I => \N__8399\
        );

    \I__1924\ : Span12Mux_h
    port map (
            O => \N__8402\,
            I => \N__8396\
        );

    \I__1923\ : Odrv12
    port map (
            O => \N__8399\,
            I => \DRA_c_4\
        );

    \I__1922\ : Odrv12
    port map (
            O => \N__8396\,
            I => \DRA_c_4\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8391\,
            I => \N__8388\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__8388\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8385\,
            I => \N__8382\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__8382\,
            I => \N__8378\
        );

    \I__1917\ : InMux
    port map (
            O => \N__8381\,
            I => \N__8375\
        );

    \I__1916\ : Span4Mux_h
    port map (
            O => \N__8378\,
            I => \N__8370\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__8375\,
            I => \N__8370\
        );

    \I__1914\ : Span4Mux_v
    port map (
            O => \N__8370\,
            I => \N__8367\
        );

    \I__1913\ : Sp12to4
    port map (
            O => \N__8367\,
            I => \N__8364\
        );

    \I__1912\ : Span12Mux_h
    port map (
            O => \N__8364\,
            I => \N__8361\
        );

    \I__1911\ : Odrv12
    port map (
            O => \N__8361\,
            I => \DRA_c_8\
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__8358\,
            I => \N__8355\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8352\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8352\,
            I => \N__8349\
        );

    \I__1907\ : Span4Mux_v
    port map (
            O => \N__8349\,
            I => \N__8346\
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__8346\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1905\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8340\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8340\,
            I => \N__8336\
        );

    \I__1903\ : InMux
    port map (
            O => \N__8339\,
            I => \N__8333\
        );

    \I__1902\ : Span4Mux_v
    port map (
            O => \N__8336\,
            I => \N__8330\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__8333\,
            I => \N__8327\
        );

    \I__1900\ : Sp12to4
    port map (
            O => \N__8330\,
            I => \N__8324\
        );

    \I__1899\ : Span12Mux_v
    port map (
            O => \N__8327\,
            I => \N__8321\
        );

    \I__1898\ : Span12Mux_h
    port map (
            O => \N__8324\,
            I => \N__8318\
        );

    \I__1897\ : Span12Mux_h
    port map (
            O => \N__8321\,
            I => \N__8313\
        );

    \I__1896\ : Span12Mux_v
    port map (
            O => \N__8318\,
            I => \N__8313\
        );

    \I__1895\ : Odrv12
    port map (
            O => \N__8313\,
            I => \DRA_c_5\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8310\,
            I => \N__8307\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__8307\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1892\ : InMux
    port map (
            O => \N__8304\,
            I => \N__8300\
        );

    \I__1891\ : InMux
    port map (
            O => \N__8303\,
            I => \N__8297\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__8300\,
            I => \N__8292\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__8297\,
            I => \N__8292\
        );

    \I__1888\ : Span4Mux_h
    port map (
            O => \N__8292\,
            I => \N__8289\
        );

    \I__1887\ : Sp12to4
    port map (
            O => \N__8289\,
            I => \N__8286\
        );

    \I__1886\ : Span12Mux_v
    port map (
            O => \N__8286\,
            I => \N__8283\
        );

    \I__1885\ : Odrv12
    port map (
            O => \N__8283\,
            I => \DRA_c_6\
        );

    \I__1884\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8277\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__8277\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8274\,
            I => \N__8271\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__8271\,
            I => \N__8267\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8270\,
            I => \N__8264\
        );

    \I__1879\ : Span4Mux_h
    port map (
            O => \N__8267\,
            I => \N__8261\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8264\,
            I => \N__8258\
        );

    \I__1877\ : Span4Mux_v
    port map (
            O => \N__8261\,
            I => \N__8255\
        );

    \I__1876\ : Sp12to4
    port map (
            O => \N__8258\,
            I => \N__8252\
        );

    \I__1875\ : Sp12to4
    port map (
            O => \N__8255\,
            I => \N__8247\
        );

    \I__1874\ : Span12Mux_v
    port map (
            O => \N__8252\,
            I => \N__8247\
        );

    \I__1873\ : Span12Mux_h
    port map (
            O => \N__8247\,
            I => \N__8244\
        );

    \I__1872\ : Odrv12
    port map (
            O => \N__8244\,
            I => \DRA_c_7\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8241\,
            I => \N__8238\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8238\,
            I => \N__8235\
        );

    \I__1869\ : Odrv12
    port map (
            O => \N__8235\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8232\,
            I => \N__8228\
        );

    \I__1867\ : InMux
    port map (
            O => \N__8231\,
            I => \N__8225\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__8228\,
            I => \N__8222\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8225\,
            I => \N__8219\
        );

    \I__1864\ : Span4Mux_v
    port map (
            O => \N__8222\,
            I => \N__8214\
        );

    \I__1863\ : Span4Mux_h
    port map (
            O => \N__8219\,
            I => \N__8214\
        );

    \I__1862\ : Sp12to4
    port map (
            O => \N__8214\,
            I => \N__8211\
        );

    \I__1861\ : Span12Mux_v
    port map (
            O => \N__8211\,
            I => \N__8208\
        );

    \I__1860\ : Span12Mux_h
    port map (
            O => \N__8208\,
            I => \N__8205\
        );

    \I__1859\ : Odrv12
    port map (
            O => \N__8205\,
            I => \DRA_c_0\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8202\,
            I => \N__8199\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__8199\,
            I => \N__8196\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__8196\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1855\ : CEMux
    port map (
            O => \N__8193\,
            I => \N__8190\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8190\,
            I => \N__8187\
        );

    \I__1853\ : Span4Mux_h
    port map (
            O => \N__8187\,
            I => \N__8182\
        );

    \I__1852\ : CEMux
    port map (
            O => \N__8186\,
            I => \N__8179\
        );

    \I__1851\ : CEMux
    port map (
            O => \N__8185\,
            I => \N__8176\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__8182\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8179\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8176\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8169\,
            I => \N__8166\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__8166\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__8163\,
            I => \N__8148\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8162\,
            I => \N__8145\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8161\,
            I => \N__8139\
        );

    \I__1842\ : InMux
    port map (
            O => \N__8160\,
            I => \N__8132\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8159\,
            I => \N__8132\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8158\,
            I => \N__8132\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8157\,
            I => \N__8125\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8156\,
            I => \N__8125\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8122\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8154\,
            I => \N__8119\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8153\,
            I => \N__8112\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8105\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8151\,
            I => \N__8105\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8148\,
            I => \N__8105\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__8145\,
            I => \N__8101\
        );

    \I__1830\ : InMux
    port map (
            O => \N__8144\,
            I => \N__8098\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8143\,
            I => \N__8095\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8142\,
            I => \N__8092\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8139\,
            I => \N__8087\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__8132\,
            I => \N__8087\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8082\
        );

    \I__1824\ : InMux
    port map (
            O => \N__8130\,
            I => \N__8082\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8125\,
            I => \N__8077\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__8122\,
            I => \N__8077\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8119\,
            I => \N__8071\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8118\,
            I => \N__8068\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8117\,
            I => \N__8065\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8116\,
            I => \N__8060\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8115\,
            I => \N__8060\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8112\,
            I => \N__8057\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__8105\,
            I => \N__8054\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8104\,
            I => \N__8051\
        );

    \I__1813\ : Span4Mux_v
    port map (
            O => \N__8101\,
            I => \N__8044\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8098\,
            I => \N__8044\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8095\,
            I => \N__8044\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8092\,
            I => \N__8037\
        );

    \I__1809\ : Span4Mux_h
    port map (
            O => \N__8087\,
            I => \N__8037\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8082\,
            I => \N__8037\
        );

    \I__1807\ : Span4Mux_v
    port map (
            O => \N__8077\,
            I => \N__8034\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8076\,
            I => \N__8031\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8075\,
            I => \N__8026\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8074\,
            I => \N__8026\
        );

    \I__1803\ : Span4Mux_h
    port map (
            O => \N__8071\,
            I => \N__8023\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8068\,
            I => \N__8016\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8065\,
            I => \N__8016\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__8060\,
            I => \N__8016\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__8057\,
            I => \N__8009\
        );

    \I__1798\ : Span4Mux_h
    port map (
            O => \N__8054\,
            I => \N__8009\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8051\,
            I => \N__8009\
        );

    \I__1796\ : Span4Mux_v
    port map (
            O => \N__8044\,
            I => \N__8004\
        );

    \I__1795\ : Span4Mux_v
    port map (
            O => \N__8037\,
            I => \N__8004\
        );

    \I__1794\ : Odrv4
    port map (
            O => \N__8034\,
            I => \CPU_CYCLEm\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8031\,
            I => \CPU_CYCLEm\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__8026\,
            I => \CPU_CYCLEm\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__8023\,
            I => \CPU_CYCLEm\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__8016\,
            I => \CPU_CYCLEm\
        );

    \I__1789\ : Odrv4
    port map (
            O => \N__8009\,
            I => \CPU_CYCLEm\
        );

    \I__1788\ : Odrv4
    port map (
            O => \N__8004\,
            I => \CPU_CYCLEm\
        );

    \I__1787\ : InMux
    port map (
            O => \N__7989\,
            I => \N__7986\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__7986\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_6\
        );

    \I__1785\ : InMux
    port map (
            O => \N__7983\,
            I => \N__7980\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__7980\,
            I => \N__7977\
        );

    \I__1783\ : Span4Mux_h
    port map (
            O => \N__7977\,
            I => \N__7973\
        );

    \I__1782\ : InMux
    port map (
            O => \N__7976\,
            I => \N__7970\
        );

    \I__1781\ : Span4Mux_v
    port map (
            O => \N__7973\,
            I => \N__7967\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__7970\,
            I => \N__7964\
        );

    \I__1779\ : Sp12to4
    port map (
            O => \N__7967\,
            I => \N__7959\
        );

    \I__1778\ : Span12Mux_v
    port map (
            O => \N__7964\,
            I => \N__7959\
        );

    \I__1777\ : Span12Mux_h
    port map (
            O => \N__7959\,
            I => \N__7956\
        );

    \I__1776\ : Span12Mux_v
    port map (
            O => \N__7956\,
            I => \N__7953\
        );

    \I__1775\ : Odrv12
    port map (
            O => \N__7953\,
            I => \DRA_c_1\
        );

    \I__1774\ : InMux
    port map (
            O => \N__7950\,
            I => \N__7947\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__7947\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1772\ : InMux
    port map (
            O => \N__7944\,
            I => \N__7941\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__7941\,
            I => \N__7938\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__7938\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1769\ : CEMux
    port map (
            O => \N__7935\,
            I => \N__7932\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__7932\,
            I => \N__7928\
        );

    \I__1767\ : CEMux
    port map (
            O => \N__7931\,
            I => \N__7925\
        );

    \I__1766\ : Span4Mux_v
    port map (
            O => \N__7928\,
            I => \N__7920\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__7925\,
            I => \N__7917\
        );

    \I__1764\ : CEMux
    port map (
            O => \N__7924\,
            I => \N__7914\
        );

    \I__1763\ : CEMux
    port map (
            O => \N__7923\,
            I => \N__7911\
        );

    \I__1762\ : Span4Mux_h
    port map (
            O => \N__7920\,
            I => \N__7904\
        );

    \I__1761\ : Span4Mux_v
    port map (
            O => \N__7917\,
            I => \N__7904\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__7914\,
            I => \N__7904\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__7911\,
            I => \N__7901\
        );

    \I__1758\ : Span4Mux_h
    port map (
            O => \N__7904\,
            I => \N__7898\
        );

    \I__1757\ : Span4Mux_h
    port map (
            O => \N__7901\,
            I => \N__7895\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__7898\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1755\ : Odrv4
    port map (
            O => \N__7895\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1754\ : IoInMux
    port map (
            O => \N__7890\,
            I => \N__7887\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__7887\,
            I => \N__7884\
        );

    \I__1752\ : Span4Mux_s2_v
    port map (
            O => \N__7884\,
            I => \N__7881\
        );

    \I__1751\ : Span4Mux_v
    port map (
            O => \N__7881\,
            I => \N__7878\
        );

    \I__1750\ : Sp12to4
    port map (
            O => \N__7878\,
            I => \N__7875\
        );

    \I__1749\ : Odrv12
    port map (
            O => \N__7875\,
            I => \CASn_c\
        );

    \I__1748\ : IoInMux
    port map (
            O => \N__7872\,
            I => \N__7869\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__7869\,
            I => \N__7866\
        );

    \I__1746\ : Span12Mux_s1_h
    port map (
            O => \N__7866\,
            I => \N__7863\
        );

    \I__1745\ : Span12Mux_h
    port map (
            O => \N__7863\,
            I => \N__7860\
        );

    \I__1744\ : Odrv12
    port map (
            O => \N__7860\,
            I => \WEn_c\
        );

    \I__1743\ : InMux
    port map (
            O => \N__7857\,
            I => \N__7854\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__7854\,
            I => \N__7850\
        );

    \I__1741\ : InMux
    port map (
            O => \N__7853\,
            I => \N__7847\
        );

    \I__1740\ : Span4Mux_h
    port map (
            O => \N__7850\,
            I => \N__7843\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__7847\,
            I => \N__7840\
        );

    \I__1738\ : InMux
    port map (
            O => \N__7846\,
            I => \N__7835\
        );

    \I__1737\ : Span4Mux_h
    port map (
            O => \N__7843\,
            I => \N__7832\
        );

    \I__1736\ : Span4Mux_h
    port map (
            O => \N__7840\,
            I => \N__7829\
        );

    \I__1735\ : InMux
    port map (
            O => \N__7839\,
            I => \N__7826\
        );

    \I__1734\ : InMux
    port map (
            O => \N__7838\,
            I => \N__7823\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__7835\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__7832\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__7829\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__7826\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__7823\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1728\ : IoInMux
    port map (
            O => \N__7812\,
            I => \N__7809\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__7809\,
            I => \N__7806\
        );

    \I__1726\ : Span4Mux_s3_v
    port map (
            O => \N__7806\,
            I => \N__7803\
        );

    \I__1725\ : Span4Mux_h
    port map (
            O => \N__7803\,
            I => \N__7800\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__7800\,
            I => \CRCSn_c\
        );

    \I__1723\ : IoInMux
    port map (
            O => \N__7797\,
            I => \N__7794\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__7794\,
            I => \N__7791\
        );

    \I__1721\ : Span4Mux_s3_v
    port map (
            O => \N__7791\,
            I => \N__7788\
        );

    \I__1720\ : Span4Mux_v
    port map (
            O => \N__7788\,
            I => \N__7785\
        );

    \I__1719\ : Span4Mux_h
    port map (
            O => \N__7785\,
            I => \N__7782\
        );

    \I__1718\ : Odrv4
    port map (
            O => \N__7782\,
            I => \RASn_c\
        );

    \I__1717\ : InMux
    port map (
            O => \N__7779\,
            I => \N__7776\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__7776\,
            I => \U712_CHIP_RAM.N_373\
        );

    \I__1715\ : IoInMux
    port map (
            O => \N__7773\,
            I => \N__7770\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__7770\,
            I => \N__7767\
        );

    \I__1713\ : Span4Mux_s2_h
    port map (
            O => \N__7767\,
            I => \N__7764\
        );

    \I__1712\ : Span4Mux_v
    port map (
            O => \N__7764\,
            I => \N__7761\
        );

    \I__1711\ : Sp12to4
    port map (
            O => \N__7761\,
            I => \N__7758\
        );

    \I__1710\ : Span12Mux_h
    port map (
            O => \N__7758\,
            I => \N__7755\
        );

    \I__1709\ : Odrv12
    port map (
            O => \N__7755\,
            I => \CMA_c_6\
        );

    \I__1708\ : InMux
    port map (
            O => \N__7752\,
            I => \N__7749\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__7749\,
            I => \N__7746\
        );

    \I__1706\ : Odrv12
    port map (
            O => \N__7746\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1705\ : InMux
    port map (
            O => \N__7743\,
            I => \N__7740\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__7740\,
            I => \N__7737\
        );

    \I__1703\ : Span4Mux_h
    port map (
            O => \N__7737\,
            I => \N__7734\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__7734\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1701\ : InMux
    port map (
            O => \N__7731\,
            I => \N__7728\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__7728\,
            I => \N__7725\
        );

    \I__1699\ : Span12Mux_v
    port map (
            O => \N__7725\,
            I => \N__7722\
        );

    \I__1698\ : Span12Mux_h
    port map (
            O => \N__7722\,
            I => \N__7719\
        );

    \I__1697\ : Odrv12
    port map (
            O => \N__7719\,
            I => \A_c_14\
        );

    \I__1696\ : InMux
    port map (
            O => \N__7716\,
            I => \N__7713\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__7713\,
            I => \N__7710\
        );

    \I__1694\ : Span4Mux_h
    port map (
            O => \N__7710\,
            I => \N__7707\
        );

    \I__1693\ : Sp12to4
    port map (
            O => \N__7707\,
            I => \N__7704\
        );

    \I__1692\ : Span12Mux_v
    port map (
            O => \N__7704\,
            I => \N__7701\
        );

    \I__1691\ : Span12Mux_h
    port map (
            O => \N__7701\,
            I => \N__7698\
        );

    \I__1690\ : Odrv12
    port map (
            O => \N__7698\,
            I => \A_c_7\
        );

    \I__1689\ : InMux
    port map (
            O => \N__7695\,
            I => \N__7692\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__7692\,
            I => \N__7689\
        );

    \I__1687\ : Span4Mux_v
    port map (
            O => \N__7689\,
            I => \N__7686\
        );

    \I__1686\ : Sp12to4
    port map (
            O => \N__7686\,
            I => \N__7683\
        );

    \I__1685\ : Span12Mux_h
    port map (
            O => \N__7683\,
            I => \N__7680\
        );

    \I__1684\ : Odrv12
    port map (
            O => \N__7680\,
            I => \A_c_13\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__7677\,
            I => \N__7674\
        );

    \I__1682\ : InMux
    port map (
            O => \N__7674\,
            I => \N__7671\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__7671\,
            I => \N__7668\
        );

    \I__1680\ : Span4Mux_v
    port map (
            O => \N__7668\,
            I => \N__7665\
        );

    \I__1679\ : Sp12to4
    port map (
            O => \N__7665\,
            I => \N__7662\
        );

    \I__1678\ : Span12Mux_h
    port map (
            O => \N__7662\,
            I => \N__7659\
        );

    \I__1677\ : Span12Mux_v
    port map (
            O => \N__7659\,
            I => \N__7656\
        );

    \I__1676\ : Odrv12
    port map (
            O => \N__7656\,
            I => \A_c_6\
        );

    \I__1675\ : InMux
    port map (
            O => \N__7653\,
            I => \N__7650\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__7650\,
            I => \U712_CHIP_RAM.N_371\
        );

    \I__1673\ : InMux
    port map (
            O => \N__7647\,
            I => \N__7644\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__7644\,
            I => \N__7641\
        );

    \I__1671\ : Span4Mux_v
    port map (
            O => \N__7641\,
            I => \N__7638\
        );

    \I__1670\ : Sp12to4
    port map (
            O => \N__7638\,
            I => \N__7635\
        );

    \I__1669\ : Span12Mux_h
    port map (
            O => \N__7635\,
            I => \N__7632\
        );

    \I__1668\ : Odrv12
    port map (
            O => \N__7632\,
            I => \A_c_15\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__7629\,
            I => \N__7626\
        );

    \I__1666\ : InMux
    port map (
            O => \N__7626\,
            I => \N__7623\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__7623\,
            I => \N__7620\
        );

    \I__1664\ : Span12Mux_v
    port map (
            O => \N__7620\,
            I => \N__7617\
        );

    \I__1663\ : Span12Mux_h
    port map (
            O => \N__7617\,
            I => \N__7614\
        );

    \I__1662\ : Odrv12
    port map (
            O => \N__7614\,
            I => \A_c_8\
        );

    \I__1661\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7608\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7608\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_5\
        );

    \I__1659\ : InMux
    port map (
            O => \N__7605\,
            I => \N__7602\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__7602\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1657\ : InMux
    port map (
            O => \N__7599\,
            I => \N__7596\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__7596\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_4\
        );

    \I__1655\ : InMux
    port map (
            O => \N__7593\,
            I => \N__7590\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__7590\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1653\ : InMux
    port map (
            O => \N__7587\,
            I => \N__7584\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__7584\,
            I => \N__7580\
        );

    \I__1651\ : InMux
    port map (
            O => \N__7583\,
            I => \N__7577\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__7580\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__7577\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7572\,
            I => \N__7568\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7565\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__7568\,
            I => \N__7560\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__7565\,
            I => \N__7560\
        );

    \I__1644\ : Span4Mux_v
    port map (
            O => \N__7560\,
            I => \N__7556\
        );

    \I__1643\ : InMux
    port map (
            O => \N__7559\,
            I => \N__7553\
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__7556\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7553\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1640\ : IoInMux
    port map (
            O => \N__7548\,
            I => \N__7545\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__7545\,
            I => \N__7542\
        );

    \I__1638\ : Span4Mux_s2_v
    port map (
            O => \N__7542\,
            I => \N__7539\
        );

    \I__1637\ : Span4Mux_v
    port map (
            O => \N__7539\,
            I => \N__7536\
        );

    \I__1636\ : Sp12to4
    port map (
            O => \N__7536\,
            I => \N__7533\
        );

    \I__1635\ : Span12Mux_h
    port map (
            O => \N__7533\,
            I => \N__7530\
        );

    \I__1634\ : Odrv12
    port map (
            O => \N__7530\,
            I => \U712_REG_SM_un1_UDSn_i\
        );

    \I__1633\ : CascadeMux
    port map (
            O => \N__7527\,
            I => \N__7524\
        );

    \I__1632\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7513\
        );

    \I__1631\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7513\
        );

    \I__1630\ : InMux
    port map (
            O => \N__7522\,
            I => \N__7510\
        );

    \I__1629\ : InMux
    port map (
            O => \N__7521\,
            I => \N__7507\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7520\,
            I => \N__7504\
        );

    \I__1627\ : InMux
    port map (
            O => \N__7519\,
            I => \N__7498\
        );

    \I__1626\ : InMux
    port map (
            O => \N__7518\,
            I => \N__7498\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__7513\,
            I => \N__7491\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7510\,
            I => \N__7491\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7507\,
            I => \N__7491\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__7504\,
            I => \N__7488\
        );

    \I__1621\ : InMux
    port map (
            O => \N__7503\,
            I => \N__7485\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__7498\,
            I => \N__7482\
        );

    \I__1619\ : Span4Mux_h
    port map (
            O => \N__7491\,
            I => \N__7479\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__7488\,
            I => \N__7474\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__7485\,
            I => \N__7474\
        );

    \I__1616\ : Span4Mux_v
    port map (
            O => \N__7482\,
            I => \N__7470\
        );

    \I__1615\ : Span4Mux_v
    port map (
            O => \N__7479\,
            I => \N__7465\
        );

    \I__1614\ : Span4Mux_h
    port map (
            O => \N__7474\,
            I => \N__7465\
        );

    \I__1613\ : InMux
    port map (
            O => \N__7473\,
            I => \N__7462\
        );

    \I__1612\ : Span4Mux_v
    port map (
            O => \N__7470\,
            I => \N__7459\
        );

    \I__1611\ : Sp12to4
    port map (
            O => \N__7465\,
            I => \N__7454\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__7462\,
            I => \N__7454\
        );

    \I__1609\ : Sp12to4
    port map (
            O => \N__7459\,
            I => \N__7451\
        );

    \I__1608\ : Span12Mux_v
    port map (
            O => \N__7454\,
            I => \N__7448\
        );

    \I__1607\ : Span12Mux_h
    port map (
            O => \N__7451\,
            I => \N__7445\
        );

    \I__1606\ : Span12Mux_h
    port map (
            O => \N__7448\,
            I => \N__7442\
        );

    \I__1605\ : Odrv12
    port map (
            O => \N__7445\,
            I => \RESETn_c\
        );

    \I__1604\ : Odrv12
    port map (
            O => \N__7442\,
            I => \RESETn_c\
        );

    \I__1603\ : IoInMux
    port map (
            O => \N__7437\,
            I => \N__7434\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__7434\,
            I => \N__7431\
        );

    \I__1601\ : Span12Mux_s5_v
    port map (
            O => \N__7431\,
            I => \N__7428\
        );

    \I__1600\ : Odrv12
    port map (
            O => \N__7428\,
            I => \RESETn_c_i\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7425\,
            I => \N__7421\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__7424\,
            I => \N__7417\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__7421\,
            I => \N__7414\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7420\,
            I => \N__7410\
        );

    \I__1595\ : InMux
    port map (
            O => \N__7417\,
            I => \N__7407\
        );

    \I__1594\ : Span4Mux_v
    port map (
            O => \N__7414\,
            I => \N__7404\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7413\,
            I => \N__7401\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__7410\,
            I => \N__7398\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__7407\,
            I => \N__7391\
        );

    \I__1590\ : Sp12to4
    port map (
            O => \N__7404\,
            I => \N__7391\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7401\,
            I => \N__7391\
        );

    \I__1588\ : Sp12to4
    port map (
            O => \N__7398\,
            I => \N__7388\
        );

    \I__1587\ : Span12Mux_h
    port map (
            O => \N__7391\,
            I => \N__7385\
        );

    \I__1586\ : Span12Mux_v
    port map (
            O => \N__7388\,
            I => \N__7382\
        );

    \I__1585\ : Span12Mux_v
    port map (
            O => \N__7385\,
            I => \N__7377\
        );

    \I__1584\ : Span12Mux_h
    port map (
            O => \N__7382\,
            I => \N__7377\
        );

    \I__1583\ : Odrv12
    port map (
            O => \N__7377\,
            I => \RnW_c\
        );

    \I__1582\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7370\
        );

    \I__1581\ : InMux
    port map (
            O => \N__7373\,
            I => \N__7367\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__7370\,
            I => \N__7364\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__7367\,
            I => \N__7361\
        );

    \I__1578\ : Span4Mux_v
    port map (
            O => \N__7364\,
            I => \N__7358\
        );

    \I__1577\ : Span12Mux_h
    port map (
            O => \N__7361\,
            I => \N__7355\
        );

    \I__1576\ : Sp12to4
    port map (
            O => \N__7358\,
            I => \N__7352\
        );

    \I__1575\ : Span12Mux_v
    port map (
            O => \N__7355\,
            I => \N__7349\
        );

    \I__1574\ : Span12Mux_v
    port map (
            O => \N__7352\,
            I => \N__7346\
        );

    \I__1573\ : Odrv12
    port map (
            O => \N__7349\,
            I => \SIZ_c_0\
        );

    \I__1572\ : Odrv12
    port map (
            O => \N__7346\,
            I => \SIZ_c_0\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__7341\,
            I => \N__7337\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__7340\,
            I => \N__7334\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7337\,
            I => \N__7329\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7334\,
            I => \N__7329\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__7329\,
            I => \N__7326\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__7326\,
            I => \U712_REG_SM.LDS_OUT_2_0_a3_0_a3Z0Z_0\
        );

    \I__1565\ : IoInMux
    port map (
            O => \N__7323\,
            I => \N__7320\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__7320\,
            I => \N__7317\
        );

    \I__1563\ : Span4Mux_s0_v
    port map (
            O => \N__7317\,
            I => \N__7314\
        );

    \I__1562\ : Span4Mux_v
    port map (
            O => \N__7314\,
            I => \N__7311\
        );

    \I__1561\ : Span4Mux_v
    port map (
            O => \N__7311\,
            I => \N__7308\
        );

    \I__1560\ : Span4Mux_h
    port map (
            O => \N__7308\,
            I => \N__7305\
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__7305\,
            I => \CMA_c_10\
        );

    \I__1558\ : IoInMux
    port map (
            O => \N__7302\,
            I => \N__7299\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7299\,
            I => \N__7296\
        );

    \I__1556\ : IoSpan4Mux
    port map (
            O => \N__7296\,
            I => \N__7293\
        );

    \I__1555\ : IoSpan4Mux
    port map (
            O => \N__7293\,
            I => \N__7290\
        );

    \I__1554\ : Span4Mux_s2_h
    port map (
            O => \N__7290\,
            I => \N__7287\
        );

    \I__1553\ : Sp12to4
    port map (
            O => \N__7287\,
            I => \N__7284\
        );

    \I__1552\ : Odrv12
    port map (
            O => \N__7284\,
            I => \CMA_c_4\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7281\,
            I => \N__7277\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7280\,
            I => \N__7274\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7277\,
            I => \N__7271\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7274\,
            I => \N__7268\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__7271\,
            I => \U712_CHIP_RAM.CMA_5_i_0_8\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__7268\,
            I => \U712_CHIP_RAM.CMA_5_i_0_8\
        );

    \I__1545\ : InMux
    port map (
            O => \N__7263\,
            I => \N__7260\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7260\,
            I => \N__7257\
        );

    \I__1543\ : Span4Mux_v
    port map (
            O => \N__7257\,
            I => \N__7254\
        );

    \I__1542\ : Sp12to4
    port map (
            O => \N__7254\,
            I => \N__7251\
        );

    \I__1541\ : Span12Mux_h
    port map (
            O => \N__7251\,
            I => \N__7248\
        );

    \I__1540\ : Odrv12
    port map (
            O => \N__7248\,
            I => \A_c_17\
        );

    \I__1539\ : IoInMux
    port map (
            O => \N__7245\,
            I => \N__7242\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7242\,
            I => \N__7239\
        );

    \I__1537\ : Span4Mux_s2_h
    port map (
            O => \N__7239\,
            I => \N__7236\
        );

    \I__1536\ : Span4Mux_v
    port map (
            O => \N__7236\,
            I => \N__7233\
        );

    \I__1535\ : Span4Mux_h
    port map (
            O => \N__7233\,
            I => \N__7230\
        );

    \I__1534\ : Sp12to4
    port map (
            O => \N__7230\,
            I => \N__7227\
        );

    \I__1533\ : Odrv12
    port map (
            O => \N__7227\,
            I => \CMA_c_8\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7224\,
            I => \N__7221\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__7221\,
            I => \N__7218\
        );

    \I__1530\ : Span4Mux_v
    port map (
            O => \N__7218\,
            I => \N__7215\
        );

    \I__1529\ : Span4Mux_v
    port map (
            O => \N__7215\,
            I => \N__7212\
        );

    \I__1528\ : Sp12to4
    port map (
            O => \N__7212\,
            I => \N__7209\
        );

    \I__1527\ : Span12Mux_h
    port map (
            O => \N__7209\,
            I => \N__7206\
        );

    \I__1526\ : Odrv12
    port map (
            O => \N__7206\,
            I => \A_c_9\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__7203\,
            I => \N__7200\
        );

    \I__1524\ : InMux
    port map (
            O => \N__7200\,
            I => \N__7197\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7197\,
            I => \N__7194\
        );

    \I__1522\ : Span4Mux_h
    port map (
            O => \N__7194\,
            I => \N__7191\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__7191\,
            I => \N__7188\
        );

    \I__1520\ : Sp12to4
    port map (
            O => \N__7188\,
            I => \N__7185\
        );

    \I__1519\ : Span12Mux_h
    port map (
            O => \N__7185\,
            I => \N__7182\
        );

    \I__1518\ : Span12Mux_v
    port map (
            O => \N__7182\,
            I => \N__7179\
        );

    \I__1517\ : Odrv12
    port map (
            O => \N__7179\,
            I => \A_c_2\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__7176\,
            I => \U712_CHIP_RAM.N_367_cascade_\
        );

    \I__1515\ : IoInMux
    port map (
            O => \N__7173\,
            I => \N__7170\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__7170\,
            I => \N__7167\
        );

    \I__1513\ : Span4Mux_s3_v
    port map (
            O => \N__7167\,
            I => \N__7164\
        );

    \I__1512\ : Span4Mux_v
    port map (
            O => \N__7164\,
            I => \N__7161\
        );

    \I__1511\ : Span4Mux_h
    port map (
            O => \N__7161\,
            I => \N__7158\
        );

    \I__1510\ : Odrv4
    port map (
            O => \N__7158\,
            I => \CMA_c_0\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7155\,
            I => \N__7152\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7152\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_0\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7149\,
            I => \N__7143\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7148\,
            I => \N__7138\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7147\,
            I => \N__7133\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7146\,
            I => \N__7133\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7143\,
            I => \N__7130\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7142\,
            I => \N__7125\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7141\,
            I => \N__7125\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7138\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__7133\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__7130\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7125\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7116\,
            I => \N__7109\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7115\,
            I => \N__7109\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7114\,
            I => \N__7106\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__7109\,
            I => \N__7101\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7106\,
            I => \N__7101\
        );

    \I__1491\ : Span4Mux_h
    port map (
            O => \N__7101\,
            I => \N__7096\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7093\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7099\,
            I => \N__7090\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__7096\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7093\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7090\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7083\,
            I => \N__7080\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7080\,
            I => \N__7077\
        );

    \I__1483\ : Span4Mux_v
    port map (
            O => \N__7077\,
            I => \N__7074\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__7074\,
            I => \U712_BYTE_ENABLE.N_453\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__7071\,
            I => \N__7068\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7068\,
            I => \N__7065\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7065\,
            I => \N__7062\
        );

    \I__1478\ : Span4Mux_h
    port map (
            O => \N__7062\,
            I => \N__7059\
        );

    \I__1477\ : Span4Mux_h
    port map (
            O => \N__7059\,
            I => \N__7055\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7058\,
            I => \N__7052\
        );

    \I__1475\ : Odrv4
    port map (
            O => \N__7055\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3Z0Z_0\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7052\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3Z0Z_0\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7047\,
            I => \N__7043\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7046\,
            I => \N__7040\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7043\,
            I => \N__7036\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7040\,
            I => \N__7033\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7039\,
            I => \N__7030\
        );

    \I__1468\ : Odrv12
    port map (
            O => \N__7036\,
            I => \U712_BYTE_ENABLE.N_451\
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__7033\,
            I => \U712_BYTE_ENABLE.N_451\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7030\,
            I => \U712_BYTE_ENABLE.N_451\
        );

    \I__1465\ : IoInMux
    port map (
            O => \N__7023\,
            I => \N__7020\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7020\,
            I => \N__7017\
        );

    \I__1463\ : IoSpan4Mux
    port map (
            O => \N__7017\,
            I => \N__7014\
        );

    \I__1462\ : IoSpan4Mux
    port map (
            O => \N__7014\,
            I => \N__7011\
        );

    \I__1461\ : Span4Mux_s3_h
    port map (
            O => \N__7011\,
            I => \N__7008\
        );

    \I__1460\ : Sp12to4
    port map (
            O => \N__7008\,
            I => \N__7005\
        );

    \I__1459\ : Odrv12
    port map (
            O => \N__7005\,
            I => \N_50_i\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7002\,
            I => \N__6998\
        );

    \I__1457\ : InMux
    port map (
            O => \N__7001\,
            I => \N__6995\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__6998\,
            I => \N__6992\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__6995\,
            I => \N__6989\
        );

    \I__1454\ : Odrv4
    port map (
            O => \N__6992\,
            I => \U712_REG_SM.N_354\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__6989\,
            I => \U712_REG_SM.N_354\
        );

    \I__1452\ : InMux
    port map (
            O => \N__6984\,
            I => \N__6980\
        );

    \I__1451\ : InMux
    port map (
            O => \N__6983\,
            I => \N__6977\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__6980\,
            I => \U712_REG_SM.N_394\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__6977\,
            I => \U712_REG_SM.N_394\
        );

    \I__1448\ : InMux
    port map (
            O => \N__6972\,
            I => \N__6969\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__6969\,
            I => \U712_REG_SM.N_364\
        );

    \I__1446\ : InMux
    port map (
            O => \N__6966\,
            I => \N__6962\
        );

    \I__1445\ : InMux
    port map (
            O => \N__6965\,
            I => \N__6959\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__6962\,
            I => \N__6956\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__6959\,
            I => \N__6953\
        );

    \I__1442\ : Span4Mux_h
    port map (
            O => \N__6956\,
            I => \N__6948\
        );

    \I__1441\ : Span4Mux_h
    port map (
            O => \N__6953\,
            I => \N__6945\
        );

    \I__1440\ : InMux
    port map (
            O => \N__6952\,
            I => \N__6942\
        );

    \I__1439\ : InMux
    port map (
            O => \N__6951\,
            I => \N__6939\
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__6948\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1437\ : Odrv4
    port map (
            O => \N__6945\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__6942\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__6939\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1434\ : CascadeMux
    port map (
            O => \N__6930\,
            I => \N__6927\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6927\,
            I => \N__6922\
        );

    \I__1432\ : InMux
    port map (
            O => \N__6926\,
            I => \N__6919\
        );

    \I__1431\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6916\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6922\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__6919\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__6916\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6909\,
            I => \N__6904\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6908\,
            I => \N__6899\
        );

    \I__1425\ : InMux
    port map (
            O => \N__6907\,
            I => \N__6899\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__6904\,
            I => \N__6894\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__6899\,
            I => \N__6894\
        );

    \I__1422\ : Span4Mux_v
    port map (
            O => \N__6894\,
            I => \N__6889\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6884\
        );

    \I__1420\ : InMux
    port map (
            O => \N__6892\,
            I => \N__6884\
        );

    \I__1419\ : Span4Mux_h
    port map (
            O => \N__6889\,
            I => \N__6879\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__6884\,
            I => \N__6879\
        );

    \I__1417\ : Sp12to4
    port map (
            O => \N__6879\,
            I => \N__6876\
        );

    \I__1416\ : Span12Mux_v
    port map (
            O => \N__6876\,
            I => \N__6873\
        );

    \I__1415\ : Odrv12
    port map (
            O => \N__6873\,
            I => \A_c_0\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__6870\,
            I => \N__6867\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6867\,
            I => \N__6864\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6864\,
            I => \N__6857\
        );

    \I__1411\ : InMux
    port map (
            O => \N__6863\,
            I => \N__6852\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6862\,
            I => \N__6852\
        );

    \I__1409\ : InMux
    port map (
            O => \N__6861\,
            I => \N__6849\
        );

    \I__1408\ : InMux
    port map (
            O => \N__6860\,
            I => \N__6846\
        );

    \I__1407\ : Odrv4
    port map (
            O => \N__6857\,
            I => \U712_REG_SM.N_395\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__6852\,
            I => \U712_REG_SM.N_395\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__6849\,
            I => \U712_REG_SM.N_395\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__6846\,
            I => \U712_REG_SM.N_395\
        );

    \I__1403\ : InMux
    port map (
            O => \N__6837\,
            I => \N__6833\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6836\,
            I => \N__6830\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__6833\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__6830\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__1399\ : IoInMux
    port map (
            O => \N__6825\,
            I => \N__6822\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6822\,
            I => \N__6819\
        );

    \I__1397\ : Span12Mux_s5_v
    port map (
            O => \N__6819\,
            I => \N__6816\
        );

    \I__1396\ : Span12Mux_h
    port map (
            O => \N__6816\,
            I => \N__6813\
        );

    \I__1395\ : Odrv12
    port map (
            O => \N__6813\,
            I => \U712_REG_SM_un1_LDSn_i\
        );

    \I__1394\ : InMux
    port map (
            O => \N__6810\,
            I => \N__6804\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6809\,
            I => \N__6801\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6808\,
            I => \N__6798\
        );

    \I__1391\ : InMux
    port map (
            O => \N__6807\,
            I => \N__6795\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6804\,
            I => \N__6792\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__6801\,
            I => \N__6787\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__6798\,
            I => \N__6787\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__6795\,
            I => \U712_REG_SM.N_348\
        );

    \I__1386\ : Odrv4
    port map (
            O => \N__6792\,
            I => \U712_REG_SM.N_348\
        );

    \I__1385\ : Odrv4
    port map (
            O => \N__6787\,
            I => \U712_REG_SM.N_348\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6780\,
            I => \N__6775\
        );

    \I__1383\ : InMux
    port map (
            O => \N__6779\,
            I => \N__6772\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6778\,
            I => \N__6769\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__6775\,
            I => \N__6759\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__6772\,
            I => \N__6759\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6769\,
            I => \N__6759\
        );

    \I__1378\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6756\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6767\,
            I => \N__6751\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6766\,
            I => \N__6751\
        );

    \I__1375\ : Odrv4
    port map (
            O => \N__6759\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__6756\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__6751\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__6744\,
            I => \N__6740\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__6743\,
            I => \N__6737\
        );

    \I__1370\ : InMux
    port map (
            O => \N__6740\,
            I => \N__6734\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6729\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__6734\,
            I => \N__6726\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6733\,
            I => \N__6723\
        );

    \I__1366\ : InMux
    port map (
            O => \N__6732\,
            I => \N__6717\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__6729\,
            I => \N__6710\
        );

    \I__1364\ : Span4Mux_h
    port map (
            O => \N__6726\,
            I => \N__6710\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__6723\,
            I => \N__6710\
        );

    \I__1362\ : InMux
    port map (
            O => \N__6722\,
            I => \N__6705\
        );

    \I__1361\ : InMux
    port map (
            O => \N__6721\,
            I => \N__6705\
        );

    \I__1360\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6702\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__6717\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__6710\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__6705\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__6702\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6693\,
            I => \N__6688\
        );

    \I__1354\ : InMux
    port map (
            O => \N__6692\,
            I => \N__6685\
        );

    \I__1353\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6682\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__6688\,
            I => \N__6677\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6685\,
            I => \N__6677\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6682\,
            I => \U712_REG_SM.N_347\
        );

    \I__1349\ : Odrv4
    port map (
            O => \N__6677\,
            I => \U712_REG_SM.N_347\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6672\,
            I => \N__6669\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__6669\,
            I => \U712_REG_SM.N_433\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6666\,
            I => \N__6663\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__6663\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i\
        );

    \I__1344\ : InMux
    port map (
            O => \N__6660\,
            I => \N__6657\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__6657\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1342\ : InMux
    port map (
            O => \N__6654\,
            I => \N__6651\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__6651\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6648\,
            I => \N__6645\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__6645\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1338\ : CascadeMux
    port map (
            O => \N__6642\,
            I => \N__6639\
        );

    \I__1337\ : InMux
    port map (
            O => \N__6639\,
            I => \N__6636\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__6636\,
            I => \N__6633\
        );

    \I__1335\ : Span12Mux_v
    port map (
            O => \N__6633\,
            I => \N__6630\
        );

    \I__1334\ : Span12Mux_h
    port map (
            O => \N__6630\,
            I => \N__6627\
        );

    \I__1333\ : Odrv12
    port map (
            O => \N__6627\,
            I => \A_c_19\
        );

    \I__1332\ : IoInMux
    port map (
            O => \N__6624\,
            I => \N__6621\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__6621\,
            I => \N__6618\
        );

    \I__1330\ : Span4Mux_s3_h
    port map (
            O => \N__6618\,
            I => \N__6615\
        );

    \I__1329\ : Span4Mux_v
    port map (
            O => \N__6615\,
            I => \N__6612\
        );

    \I__1328\ : Sp12to4
    port map (
            O => \N__6612\,
            I => \N__6609\
        );

    \I__1327\ : Span12Mux_h
    port map (
            O => \N__6609\,
            I => \N__6606\
        );

    \I__1326\ : Odrv12
    port map (
            O => \N__6606\,
            I => \CMA_c_9\
        );

    \I__1325\ : InMux
    port map (
            O => \N__6603\,
            I => \N__6600\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6600\,
            I => \N__6597\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__6597\,
            I => \U712_CHIP_RAM.N_374\
        );

    \I__1322\ : IoInMux
    port map (
            O => \N__6594\,
            I => \N__6591\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6591\,
            I => \N__6588\
        );

    \I__1320\ : IoSpan4Mux
    port map (
            O => \N__6588\,
            I => \N__6585\
        );

    \I__1319\ : IoSpan4Mux
    port map (
            O => \N__6585\,
            I => \N__6582\
        );

    \I__1318\ : Sp12to4
    port map (
            O => \N__6582\,
            I => \N__6579\
        );

    \I__1317\ : Span12Mux_s7_h
    port map (
            O => \N__6579\,
            I => \N__6576\
        );

    \I__1316\ : Odrv12
    port map (
            O => \N__6576\,
            I => \CMA_c_7\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6573\,
            I => \N__6570\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__6570\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6567\,
            I => \N__6563\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6566\,
            I => \N__6560\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__6563\,
            I => \N__6555\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__6560\,
            I => \N__6555\
        );

    \I__1309\ : Span4Mux_v
    port map (
            O => \N__6555\,
            I => \N__6552\
        );

    \I__1308\ : Sp12to4
    port map (
            O => \N__6552\,
            I => \N__6549\
        );

    \I__1307\ : Span12Mux_h
    port map (
            O => \N__6549\,
            I => \N__6546\
        );

    \I__1306\ : Span12Mux_v
    port map (
            O => \N__6546\,
            I => \N__6543\
        );

    \I__1305\ : Odrv12
    port map (
            O => \N__6543\,
            I => \DRA_c_3\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6540\,
            I => \N__6537\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6537\,
            I => \N__6534\
        );

    \I__1302\ : Odrv12
    port map (
            O => \N__6534\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6531\,
            I => \N__6528\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6528\,
            I => \N__6524\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6527\,
            I => \N__6521\
        );

    \I__1298\ : Span4Mux_v
    port map (
            O => \N__6524\,
            I => \N__6518\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6521\,
            I => \N__6515\
        );

    \I__1296\ : Sp12to4
    port map (
            O => \N__6518\,
            I => \N__6512\
        );

    \I__1295\ : Span12Mux_h
    port map (
            O => \N__6515\,
            I => \N__6509\
        );

    \I__1294\ : Span12Mux_h
    port map (
            O => \N__6512\,
            I => \N__6506\
        );

    \I__1293\ : Span12Mux_v
    port map (
            O => \N__6509\,
            I => \N__6503\
        );

    \I__1292\ : Span12Mux_v
    port map (
            O => \N__6506\,
            I => \N__6500\
        );

    \I__1291\ : Odrv12
    port map (
            O => \N__6503\,
            I => \DRA_c_2\
        );

    \I__1290\ : Odrv12
    port map (
            O => \N__6500\,
            I => \DRA_c_2\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__6495\,
            I => \N__6492\
        );

    \I__1288\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6489\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__6489\,
            I => \N__6486\
        );

    \I__1286\ : Odrv12
    port map (
            O => \N__6486\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6483\,
            I => \N__6480\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__6480\,
            I => \N__6477\
        );

    \I__1283\ : Span4Mux_h
    port map (
            O => \N__6477\,
            I => \N__6472\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6476\,
            I => \N__6467\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6467\
        );

    \I__1280\ : Odrv4
    port map (
            O => \N__6472\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6467\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1278\ : CascadeMux
    port map (
            O => \N__6462\,
            I => \U712_REG_SM.N_364_cascade_\
        );

    \I__1277\ : InMux
    port map (
            O => \N__6459\,
            I => \N__6455\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__6458\,
            I => \N__6451\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6455\,
            I => \N__6448\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6454\,
            I => \N__6443\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6451\,
            I => \N__6443\
        );

    \I__1272\ : Span4Mux_h
    port map (
            O => \N__6448\,
            I => \N__6440\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__6443\,
            I => \U712_REG_SM.N_343\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__6440\,
            I => \U712_REG_SM.N_343\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6435\,
            I => \N__6432\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6432\,
            I => \N__6429\
        );

    \I__1267\ : Span4Mux_h
    port map (
            O => \N__6429\,
            I => \N__6425\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6428\,
            I => \N__6422\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__6425\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6422\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6417\,
            I => \N__6414\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__6414\,
            I => \N__6411\
        );

    \I__1261\ : Span12Mux_h
    port map (
            O => \N__6411\,
            I => \N__6408\
        );

    \I__1260\ : Span12Mux_v
    port map (
            O => \N__6408\,
            I => \N__6405\
        );

    \I__1259\ : Odrv12
    port map (
            O => \N__6405\,
            I => \C3_c\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__6402\,
            I => \N__6399\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6399\,
            I => \N__6395\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6398\,
            I => \N__6392\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__6395\,
            I => \N__6388\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6392\,
            I => \N__6384\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6391\,
            I => \N__6381\
        );

    \I__1252\ : Span4Mux_v
    port map (
            O => \N__6388\,
            I => \N__6378\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6387\,
            I => \N__6375\
        );

    \I__1250\ : Odrv12
    port map (
            O => \N__6384\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__6381\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__6378\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6375\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6366\,
            I => \N__6363\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6363\,
            I => \U712_CHIP_RAM.N_370\
        );

    \I__1244\ : IoInMux
    port map (
            O => \N__6360\,
            I => \N__6357\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__6357\,
            I => \N__6354\
        );

    \I__1242\ : Span4Mux_s3_h
    port map (
            O => \N__6354\,
            I => \N__6351\
        );

    \I__1241\ : Span4Mux_v
    port map (
            O => \N__6351\,
            I => \N__6348\
        );

    \I__1240\ : Span4Mux_h
    port map (
            O => \N__6348\,
            I => \N__6345\
        );

    \I__1239\ : Span4Mux_h
    port map (
            O => \N__6345\,
            I => \N__6342\
        );

    \I__1238\ : Span4Mux_h
    port map (
            O => \N__6342\,
            I => \N__6339\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__6339\,
            I => \CMA_c_3\
        );

    \I__1236\ : IoInMux
    port map (
            O => \N__6336\,
            I => \N__6333\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6333\,
            I => \N__6330\
        );

    \I__1234\ : Odrv12
    port map (
            O => \N__6330\,
            I => \CMA_c_1\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6324\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6324\,
            I => \N__6321\
        );

    \I__1231\ : Span4Mux_v
    port map (
            O => \N__6321\,
            I => \N__6318\
        );

    \I__1230\ : Sp12to4
    port map (
            O => \N__6318\,
            I => \N__6315\
        );

    \I__1229\ : Span12Mux_h
    port map (
            O => \N__6315\,
            I => \N__6312\
        );

    \I__1228\ : Span12Mux_v
    port map (
            O => \N__6312\,
            I => \N__6309\
        );

    \I__1227\ : Odrv12
    port map (
            O => \N__6309\,
            I => \A_c_3\
        );

    \I__1226\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6303\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6303\,
            I => \N__6300\
        );

    \I__1224\ : Span4Mux_v
    port map (
            O => \N__6300\,
            I => \N__6297\
        );

    \I__1223\ : Sp12to4
    port map (
            O => \N__6297\,
            I => \N__6294\
        );

    \I__1222\ : Span12Mux_h
    port map (
            O => \N__6294\,
            I => \N__6291\
        );

    \I__1221\ : Odrv12
    port map (
            O => \N__6291\,
            I => \A_c_10\
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__6288\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_1_cascade_\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6285\,
            I => \N__6282\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6282\,
            I => \U712_CHIP_RAM.N_368\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6279\,
            I => \N__6276\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__6276\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_2\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__6273\,
            I => \U712_REG_SM.N_347_cascade_\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6267\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__6267\,
            I => \U712_REG_SM.N_559\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__6264\,
            I => \U712_REG_SM.N_559_cascade_\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6261\,
            I => \N__6255\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6252\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6259\,
            I => \N__6247\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6258\,
            I => \N__6247\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6255\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__6252\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6247\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1204\ : CascadeMux
    port map (
            O => \N__6240\,
            I => \N__6237\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6237\,
            I => \N__6228\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6236\,
            I => \N__6228\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6235\,
            I => \N__6228\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6228\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6221\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6224\,
            I => \N__6218\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6221\,
            I => \U712_REG_SM.REG_CYCLE_GOZ0\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__6218\,
            I => \U712_REG_SM.REG_CYCLE_GOZ0\
        );

    \I__1195\ : IoInMux
    port map (
            O => \N__6213\,
            I => \N__6209\
        );

    \I__1194\ : IoInMux
    port map (
            O => \N__6212\,
            I => \N__6206\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6209\,
            I => \N__6203\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6206\,
            I => \N__6200\
        );

    \I__1191\ : IoSpan4Mux
    port map (
            O => \N__6203\,
            I => \N__6197\
        );

    \I__1190\ : IoSpan4Mux
    port map (
            O => \N__6200\,
            I => \N__6194\
        );

    \I__1189\ : Span4Mux_s2_v
    port map (
            O => \N__6197\,
            I => \N__6191\
        );

    \I__1188\ : Span4Mux_s2_v
    port map (
            O => \N__6194\,
            I => \N__6188\
        );

    \I__1187\ : Sp12to4
    port map (
            O => \N__6191\,
            I => \N__6185\
        );

    \I__1186\ : Sp12to4
    port map (
            O => \N__6188\,
            I => \N__6182\
        );

    \I__1185\ : Span12Mux_s8_v
    port map (
            O => \N__6185\,
            I => \N__6179\
        );

    \I__1184\ : Span12Mux_s8_v
    port map (
            O => \N__6182\,
            I => \N__6176\
        );

    \I__1183\ : Span12Mux_h
    port map (
            O => \N__6179\,
            I => \N__6171\
        );

    \I__1182\ : Span12Mux_h
    port map (
            O => \N__6176\,
            I => \N__6171\
        );

    \I__1181\ : Odrv12
    port map (
            O => \N__6171\,
            I => \ASn_c\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6168\,
            I => \N__6165\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6165\,
            I => \N__6161\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6164\,
            I => \N__6158\
        );

    \I__1177\ : Odrv4
    port map (
            O => \N__6161\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__6158\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1175\ : InMux
    port map (
            O => \N__6153\,
            I => \N__6150\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6150\,
            I => \N__6145\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6149\,
            I => \N__6142\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6148\,
            I => \N__6139\
        );

    \I__1171\ : Odrv4
    port map (
            O => \N__6145\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6142\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6139\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6132\,
            I => \N__6128\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6131\,
            I => \N__6125\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6128\,
            I => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6125\,
            I => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1\
        );

    \I__1164\ : CEMux
    port map (
            O => \N__6120\,
            I => \N__6117\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6117\,
            I => \U712_REG_SM.N_186_0\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__6114\,
            I => \U712_REG_SM.N_348_cascade_\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6111\,
            I => \N__6103\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6103\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6109\,
            I => \N__6098\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6108\,
            I => \N__6098\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6103\,
            I => \N__6094\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6098\,
            I => \N__6091\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__6097\,
            I => \N__6087\
        );

    \I__1154\ : Span4Mux_v
    port map (
            O => \N__6094\,
            I => \N__6079\
        );

    \I__1153\ : Span4Mux_v
    port map (
            O => \N__6091\,
            I => \N__6079\
        );

    \I__1152\ : InMux
    port map (
            O => \N__6090\,
            I => \N__6074\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6087\,
            I => \N__6074\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6086\,
            I => \N__6071\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6068\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6084\,
            I => \N__6065\
        );

    \I__1147\ : Odrv4
    port map (
            O => \N__6079\,
            I => \DMA_CYCLEm\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6074\,
            I => \DMA_CYCLEm\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6071\,
            I => \DMA_CYCLEm\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6068\,
            I => \DMA_CYCLEm\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6065\,
            I => \DMA_CYCLEm\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__6054\,
            I => \N__6047\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6053\,
            I => \N__6042\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6042\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__6051\,
            I => \N__6039\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__6050\,
            I => \N__6034\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6047\,
            I => \N__6031\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6042\,
            I => \N__6028\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6039\,
            I => \N__6023\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6023\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6018\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6034\,
            I => \N__6018\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6031\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1130\ : Odrv4
    port map (
            O => \N__6028\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6023\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6018\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6009\,
            I => \N__6005\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6008\,
            I => \N__6002\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6005\,
            I => \U712_REG_SM.N_361\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6002\,
            I => \U712_REG_SM.N_361\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__5997\,
            I => \N__5994\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5994\,
            I => \N__5990\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5993\,
            I => \N__5986\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__5990\,
            I => \N__5983\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5989\,
            I => \N__5980\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5986\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__5983\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5980\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5973\,
            I => \N__5970\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__5970\,
            I => \N__5967\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__5967\,
            I => \N__5964\
        );

    \I__1112\ : Sp12to4
    port map (
            O => \N__5964\,
            I => \N__5961\
        );

    \I__1111\ : Span12Mux_h
    port map (
            O => \N__5961\,
            I => \N__5958\
        );

    \I__1110\ : Span12Mux_v
    port map (
            O => \N__5958\,
            I => \N__5955\
        );

    \I__1109\ : Odrv12
    port map (
            O => \N__5955\,
            I => \DBRn_c\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5952\,
            I => \N__5949\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__5949\,
            I => \N__5943\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5948\,
            I => \N__5938\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5947\,
            I => \N__5938\
        );

    \I__1104\ : InMux
    port map (
            O => \N__5946\,
            I => \N__5934\
        );

    \I__1103\ : Span4Mux_h
    port map (
            O => \N__5943\,
            I => \N__5931\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5938\,
            I => \N__5928\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5937\,
            I => \N__5925\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5934\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1099\ : Odrv4
    port map (
            O => \N__5931\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1098\ : Odrv4
    port map (
            O => \N__5928\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5925\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5916\,
            I => \N__5913\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5913\,
            I => \N__5908\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5912\,
            I => \N__5903\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5903\
        );

    \I__1092\ : Span4Mux_h
    port map (
            O => \N__5908\,
            I => \N__5897\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5903\,
            I => \N__5897\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5894\
        );

    \I__1089\ : Odrv4
    port map (
            O => \N__5897\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5894\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5889\,
            I => \N__5885\
        );

    \I__1086\ : IoInMux
    port map (
            O => \N__5888\,
            I => \N__5882\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5885\,
            I => \N__5879\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__5882\,
            I => \N__5876\
        );

    \I__1083\ : Sp12to4
    port map (
            O => \N__5879\,
            I => \N__5873\
        );

    \I__1082\ : Span4Mux_s3_h
    port map (
            O => \N__5876\,
            I => \N__5870\
        );

    \I__1081\ : Span12Mux_v
    port map (
            O => \N__5873\,
            I => \N__5867\
        );

    \I__1080\ : Sp12to4
    port map (
            O => \N__5870\,
            I => \N__5864\
        );

    \I__1079\ : Span12Mux_h
    port map (
            O => \N__5867\,
            I => \N__5861\
        );

    \I__1078\ : Span12Mux_v
    port map (
            O => \N__5864\,
            I => \N__5858\
        );

    \I__1077\ : Odrv12
    port map (
            O => \N__5861\,
            I => \C1_c\
        );

    \I__1076\ : Odrv12
    port map (
            O => \N__5858\,
            I => \C1_c\
        );

    \I__1075\ : InMux
    port map (
            O => \N__5853\,
            I => \N__5849\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5846\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__5849\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5846\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__5841\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_2_1_cascade_\
        );

    \I__1070\ : CascadeMux
    port map (
            O => \N__5838\,
            I => \N__5835\
        );

    \I__1069\ : InMux
    port map (
            O => \N__5835\,
            I => \N__5832\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__5832\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_2\
        );

    \I__1067\ : InMux
    port map (
            O => \N__5829\,
            I => \N__5822\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5828\,
            I => \N__5822\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5827\,
            I => \N__5819\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__5822\,
            I => \N__5816\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__5819\,
            I => \N__5813\
        );

    \I__1062\ : Span4Mux_h
    port map (
            O => \N__5816\,
            I => \N__5810\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__5813\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3\
        );

    \I__1060\ : Odrv4
    port map (
            O => \N__5810\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__5805\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3_cascade_\
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__5802\,
            I => \N__5799\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5799\,
            I => \N__5792\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5786\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5786\
        );

    \I__1054\ : CascadeMux
    port map (
            O => \N__5796\,
            I => \N__5779\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5795\,
            I => \N__5775\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5792\,
            I => \N__5772\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5791\,
            I => \N__5769\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__5786\,
            I => \N__5766\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5785\,
            I => \N__5757\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5757\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5757\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5782\,
            I => \N__5757\
        );

    \I__1045\ : InMux
    port map (
            O => \N__5779\,
            I => \N__5752\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5778\,
            I => \N__5752\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5775\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1042\ : Odrv4
    port map (
            O => \N__5772\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5769\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1040\ : Odrv4
    port map (
            O => \N__5766\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__5757\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__5752\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__5739\,
            I => \N__5736\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5736\,
            I => \N__5733\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5733\,
            I => \N__5730\
        );

    \I__1034\ : Odrv4
    port map (
            O => \N__5730\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_3\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5727\,
            I => \N__5718\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5726\,
            I => \N__5718\
        );

    \I__1031\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5718\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5718\,
            I => \U712_CHIP_RAM.N_52\
        );

    \I__1029\ : InMux
    port map (
            O => \N__5715\,
            I => \N__5712\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__5712\,
            I => \N__5704\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5711\,
            I => \N__5701\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5710\,
            I => \N__5696\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5709\,
            I => \N__5691\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5708\,
            I => \N__5691\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5707\,
            I => \N__5688\
        );

    \I__1022\ : Span4Mux_h
    port map (
            O => \N__5704\,
            I => \N__5683\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__5701\,
            I => \N__5683\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5700\,
            I => \N__5680\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5699\,
            I => \N__5666\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5696\,
            I => \N__5661\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5691\,
            I => \N__5661\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5688\,
            I => \N__5654\
        );

    \I__1015\ : Span4Mux_v
    port map (
            O => \N__5683\,
            I => \N__5654\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5680\,
            I => \N__5654\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5679\,
            I => \N__5647\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5647\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5677\,
            I => \N__5647\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5638\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5675\,
            I => \N__5638\
        );

    \I__1008\ : InMux
    port map (
            O => \N__5674\,
            I => \N__5638\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5673\,
            I => \N__5638\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5672\,
            I => \N__5631\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5631\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5631\
        );

    \I__1003\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5628\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__5666\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1001\ : Odrv4
    port map (
            O => \N__5661\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1000\ : Odrv4
    port map (
            O => \N__5654\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5647\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__5638\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5631\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5628\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__5613\,
            I => \N__5610\
        );

    \I__994\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5604\
        );

    \I__993\ : InMux
    port map (
            O => \N__5609\,
            I => \N__5600\
        );

    \I__992\ : InMux
    port map (
            O => \N__5608\,
            I => \N__5594\
        );

    \I__991\ : InMux
    port map (
            O => \N__5607\,
            I => \N__5594\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__5604\,
            I => \N__5591\
        );

    \I__989\ : CascadeMux
    port map (
            O => \N__5603\,
            I => \N__5587\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5600\,
            I => \N__5583\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__5599\,
            I => \N__5579\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5594\,
            I => \N__5568\
        );

    \I__985\ : Span4Mux_h
    port map (
            O => \N__5591\,
            I => \N__5568\
        );

    \I__984\ : InMux
    port map (
            O => \N__5590\,
            I => \N__5565\
        );

    \I__983\ : InMux
    port map (
            O => \N__5587\,
            I => \N__5560\
        );

    \I__982\ : InMux
    port map (
            O => \N__5586\,
            I => \N__5560\
        );

    \I__981\ : Span4Mux_h
    port map (
            O => \N__5583\,
            I => \N__5557\
        );

    \I__980\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5548\
        );

    \I__979\ : InMux
    port map (
            O => \N__5579\,
            I => \N__5548\
        );

    \I__978\ : InMux
    port map (
            O => \N__5578\,
            I => \N__5548\
        );

    \I__977\ : InMux
    port map (
            O => \N__5577\,
            I => \N__5548\
        );

    \I__976\ : InMux
    port map (
            O => \N__5576\,
            I => \N__5543\
        );

    \I__975\ : InMux
    port map (
            O => \N__5575\,
            I => \N__5543\
        );

    \I__974\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5540\
        );

    \I__973\ : InMux
    port map (
            O => \N__5573\,
            I => \N__5537\
        );

    \I__972\ : Odrv4
    port map (
            O => \N__5568\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__5565\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5560\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__969\ : Odrv4
    port map (
            O => \N__5557\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5548\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__5543\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5540\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__5537\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__964\ : CascadeMux
    port map (
            O => \N__5520\,
            I => \N__5515\
        );

    \I__963\ : CascadeMux
    port map (
            O => \N__5519\,
            I => \N__5511\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__5518\,
            I => \N__5506\
        );

    \I__961\ : InMux
    port map (
            O => \N__5515\,
            I => \N__5498\
        );

    \I__960\ : InMux
    port map (
            O => \N__5514\,
            I => \N__5495\
        );

    \I__959\ : InMux
    port map (
            O => \N__5511\,
            I => \N__5488\
        );

    \I__958\ : InMux
    port map (
            O => \N__5510\,
            I => \N__5488\
        );

    \I__957\ : InMux
    port map (
            O => \N__5509\,
            I => \N__5488\
        );

    \I__956\ : InMux
    port map (
            O => \N__5506\,
            I => \N__5485\
        );

    \I__955\ : InMux
    port map (
            O => \N__5505\,
            I => \N__5480\
        );

    \I__954\ : InMux
    port map (
            O => \N__5504\,
            I => \N__5480\
        );

    \I__953\ : InMux
    port map (
            O => \N__5503\,
            I => \N__5473\
        );

    \I__952\ : InMux
    port map (
            O => \N__5502\,
            I => \N__5473\
        );

    \I__951\ : InMux
    port map (
            O => \N__5501\,
            I => \N__5473\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5498\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5495\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5488\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__5485\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__5480\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__5473\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__944\ : InMux
    port map (
            O => \N__5460\,
            I => \N__5456\
        );

    \I__943\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5453\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5456\,
            I => \N__5450\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5453\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__940\ : Odrv12
    port map (
            O => \N__5450\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__939\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5442\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5442\,
            I => \N__5439\
        );

    \I__937\ : Odrv12
    port map (
            O => \N__5439\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__5436\,
            I => \N__5433\
        );

    \I__935\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5430\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5430\,
            I => \N__5426\
        );

    \I__933\ : InMux
    port map (
            O => \N__5429\,
            I => \N__5423\
        );

    \I__932\ : Span4Mux_h
    port map (
            O => \N__5426\,
            I => \N__5420\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5423\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__930\ : Odrv4
    port map (
            O => \N__5420\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__929\ : InMux
    port map (
            O => \N__5415\,
            I => \N__5412\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5412\,
            I => \N__5409\
        );

    \I__927\ : Odrv12
    port map (
            O => \N__5409\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__926\ : InMux
    port map (
            O => \N__5406\,
            I => \N__5403\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__5403\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__924\ : InMux
    port map (
            O => \N__5400\,
            I => \N__5397\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5397\,
            I => \N__5394\
        );

    \I__922\ : Span4Mux_h
    port map (
            O => \N__5394\,
            I => \N__5389\
        );

    \I__921\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5384\
        );

    \I__920\ : InMux
    port map (
            O => \N__5392\,
            I => \N__5384\
        );

    \I__919\ : Odrv4
    port map (
            O => \N__5389\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5384\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__917\ : InMux
    port map (
            O => \N__5379\,
            I => \N__5376\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5376\,
            I => \N__5372\
        );

    \I__915\ : InMux
    port map (
            O => \N__5375\,
            I => \N__5369\
        );

    \I__914\ : Span4Mux_v
    port map (
            O => \N__5372\,
            I => \N__5366\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5369\,
            I => \N__5363\
        );

    \I__912\ : Span4Mux_v
    port map (
            O => \N__5366\,
            I => \N__5360\
        );

    \I__911\ : Span4Mux_v
    port map (
            O => \N__5363\,
            I => \N__5357\
        );

    \I__910\ : Sp12to4
    port map (
            O => \N__5360\,
            I => \N__5352\
        );

    \I__909\ : Sp12to4
    port map (
            O => \N__5357\,
            I => \N__5352\
        );

    \I__908\ : Span12Mux_h
    port map (
            O => \N__5352\,
            I => \N__5349\
        );

    \I__907\ : Span12Mux_v
    port map (
            O => \N__5349\,
            I => \N__5346\
        );

    \I__906\ : Odrv12
    port map (
            O => \N__5346\,
            I => \TSn_c\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__5343\,
            I => \N__5340\
        );

    \I__904\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5337\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5337\,
            I => \N__5334\
        );

    \I__902\ : Span4Mux_v
    port map (
            O => \N__5334\,
            I => \N__5331\
        );

    \I__901\ : Span4Mux_h
    port map (
            O => \N__5331\,
            I => \N__5327\
        );

    \I__900\ : IoInMux
    port map (
            O => \N__5330\,
            I => \N__5324\
        );

    \I__899\ : Sp12to4
    port map (
            O => \N__5327\,
            I => \N__5321\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__5324\,
            I => \N__5318\
        );

    \I__897\ : Span12Mux_v
    port map (
            O => \N__5321\,
            I => \N__5315\
        );

    \I__896\ : IoSpan4Mux
    port map (
            O => \N__5318\,
            I => \N__5312\
        );

    \I__895\ : Odrv12
    port map (
            O => \N__5315\,
            I => \RAMENn_c\
        );

    \I__894\ : Odrv4
    port map (
            O => \N__5312\,
            I => \RAMENn_c\
        );

    \I__893\ : InMux
    port map (
            O => \N__5307\,
            I => \N__5303\
        );

    \I__892\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5297\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__5303\,
            I => \N__5294\
        );

    \I__890\ : InMux
    port map (
            O => \N__5302\,
            I => \N__5289\
        );

    \I__889\ : InMux
    port map (
            O => \N__5301\,
            I => \N__5289\
        );

    \I__888\ : InMux
    port map (
            O => \N__5300\,
            I => \N__5286\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5297\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__886\ : Odrv4
    port map (
            O => \N__5294\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5289\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5286\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__883\ : InMux
    port map (
            O => \N__5277\,
            I => \N__5274\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__5274\,
            I => \N__5270\
        );

    \I__881\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5267\
        );

    \I__880\ : Odrv4
    port map (
            O => \N__5270\,
            I => \U712_CHIP_RAM.N_492\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5267\,
            I => \U712_CHIP_RAM.N_492\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__5262\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_tz_cascade_\
        );

    \I__877\ : InMux
    port map (
            O => \N__5259\,
            I => \N__5256\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5256\,
            I => \N__5252\
        );

    \I__875\ : InMux
    port map (
            O => \N__5255\,
            I => \N__5249\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__5252\,
            I => \U712_CHIP_RAM.N_331\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5249\,
            I => \U712_CHIP_RAM.N_331\
        );

    \I__872\ : InMux
    port map (
            O => \N__5244\,
            I => \N__5237\
        );

    \I__871\ : InMux
    port map (
            O => \N__5243\,
            I => \N__5237\
        );

    \I__870\ : InMux
    port map (
            O => \N__5242\,
            I => \N__5234\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5237\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5234\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__867\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5226\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5226\,
            I => \U712_CHIP_RAM.N_222\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__5223\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_\
        );

    \I__864\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5214\
        );

    \I__863\ : InMux
    port map (
            O => \N__5219\,
            I => \N__5209\
        );

    \I__862\ : InMux
    port map (
            O => \N__5218\,
            I => \N__5209\
        );

    \I__861\ : InMux
    port map (
            O => \N__5217\,
            I => \N__5204\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__5214\,
            I => \N__5199\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5209\,
            I => \N__5199\
        );

    \I__858\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5194\
        );

    \I__857\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5194\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__5204\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__855\ : Odrv4
    port map (
            O => \N__5199\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__5194\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__853\ : CascadeMux
    port map (
            O => \N__5187\,
            I => \N__5182\
        );

    \I__852\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5175\
        );

    \I__851\ : InMux
    port map (
            O => \N__5185\,
            I => \N__5172\
        );

    \I__850\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5169\
        );

    \I__849\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5166\
        );

    \I__848\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5163\
        );

    \I__847\ : InMux
    port map (
            O => \N__5179\,
            I => \N__5158\
        );

    \I__846\ : InMux
    port map (
            O => \N__5178\,
            I => \N__5158\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5175\,
            I => \N__5153\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5172\,
            I => \N__5153\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__5169\,
            I => \U712_CHIP_RAM.N_346\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5166\,
            I => \U712_CHIP_RAM.N_346\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5163\,
            I => \U712_CHIP_RAM.N_346\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5158\,
            I => \U712_CHIP_RAM.N_346\
        );

    \I__839\ : Odrv4
    port map (
            O => \N__5153\,
            I => \U712_CHIP_RAM.N_346\
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__5142\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_0_i_0_0_cascade_\
        );

    \I__837\ : InMux
    port map (
            O => \N__5139\,
            I => \N__5136\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__5136\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_4_0\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__5133\,
            I => \N__5127\
        );

    \I__834\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5124\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__5131\,
            I => \N__5120\
        );

    \I__832\ : InMux
    port map (
            O => \N__5130\,
            I => \N__5116\
        );

    \I__831\ : InMux
    port map (
            O => \N__5127\,
            I => \N__5113\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5124\,
            I => \N__5110\
        );

    \I__829\ : InMux
    port map (
            O => \N__5123\,
            I => \N__5105\
        );

    \I__828\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5105\
        );

    \I__827\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5102\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5116\,
            I => \U712_CHIP_RAM.N_330\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5113\,
            I => \U712_CHIP_RAM.N_330\
        );

    \I__824\ : Odrv4
    port map (
            O => \N__5110\,
            I => \U712_CHIP_RAM.N_330\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__5105\,
            I => \U712_CHIP_RAM.N_330\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5102\,
            I => \U712_CHIP_RAM.N_330\
        );

    \I__821\ : InMux
    port map (
            O => \N__5091\,
            I => \N__5088\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5088\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_5_0\
        );

    \I__819\ : InMux
    port map (
            O => \N__5085\,
            I => \N__5082\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5082\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_0_i_a3_0_1_0_0\
        );

    \I__817\ : CascadeMux
    port map (
            O => \N__5079\,
            I => \N__5076\
        );

    \I__816\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5073\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__5073\,
            I => \U712_REG_SM.N_71\
        );

    \I__814\ : IoInMux
    port map (
            O => \N__5070\,
            I => \N__5067\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5067\,
            I => \N__5064\
        );

    \I__812\ : Odrv12
    port map (
            O => \N__5064\,
            I => \CMA_c_2\
        );

    \I__811\ : IoInMux
    port map (
            O => \N__5061\,
            I => \N__5058\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__5058\,
            I => \N__5055\
        );

    \I__809\ : Span4Mux_s3_v
    port map (
            O => \N__5055\,
            I => \N__5052\
        );

    \I__808\ : Span4Mux_v
    port map (
            O => \N__5052\,
            I => \N__5049\
        );

    \I__807\ : Span4Mux_h
    port map (
            O => \N__5049\,
            I => \N__5046\
        );

    \I__806\ : Odrv4
    port map (
            O => \N__5046\,
            I => \CONSTANT_ONE_NET\
        );

    \I__805\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5040\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5040\,
            I => \N__5037\
        );

    \I__803\ : Span4Mux_v
    port map (
            O => \N__5037\,
            I => \N__5034\
        );

    \I__802\ : Sp12to4
    port map (
            O => \N__5034\,
            I => \N__5031\
        );

    \I__801\ : Span12Mux_h
    port map (
            O => \N__5031\,
            I => \N__5028\
        );

    \I__800\ : Odrv12
    port map (
            O => \N__5028\,
            I => \A_c_11\
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__5025\,
            I => \N__5022\
        );

    \I__798\ : InMux
    port map (
            O => \N__5022\,
            I => \N__5019\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5019\,
            I => \N__5016\
        );

    \I__796\ : Span4Mux_v
    port map (
            O => \N__5016\,
            I => \N__5013\
        );

    \I__795\ : Sp12to4
    port map (
            O => \N__5013\,
            I => \N__5010\
        );

    \I__794\ : Span12Mux_h
    port map (
            O => \N__5010\,
            I => \N__5007\
        );

    \I__793\ : Span12Mux_v
    port map (
            O => \N__5007\,
            I => \N__5004\
        );

    \I__792\ : Odrv12
    port map (
            O => \N__5004\,
            I => \A_c_4\
        );

    \I__791\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4998\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4998\,
            I => \U712_CHIP_RAM.N_369\
        );

    \I__789\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4992\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4992\,
            I => \U712_CHIP_RAM.N_445\
        );

    \I__787\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4986\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4986\,
            I => \N__4983\
        );

    \I__785\ : Span4Mux_v
    port map (
            O => \N__4983\,
            I => \N__4980\
        );

    \I__784\ : Sp12to4
    port map (
            O => \N__4980\,
            I => \N__4977\
        );

    \I__783\ : Span12Mux_h
    port map (
            O => \N__4977\,
            I => \N__4974\
        );

    \I__782\ : Odrv12
    port map (
            O => \N__4974\,
            I => \A_c_12\
        );

    \I__781\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4968\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4968\,
            I => \N__4965\
        );

    \I__779\ : Sp12to4
    port map (
            O => \N__4965\,
            I => \N__4962\
        );

    \I__778\ : Span12Mux_v
    port map (
            O => \N__4962\,
            I => \N__4959\
        );

    \I__777\ : Span12Mux_h
    port map (
            O => \N__4959\,
            I => \N__4956\
        );

    \I__776\ : Odrv12
    port map (
            O => \N__4956\,
            I => \A_c_5\
        );

    \I__775\ : SRMux
    port map (
            O => \N__4953\,
            I => \N__4950\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4950\,
            I => \N__4947\
        );

    \I__773\ : Span4Mux_h
    port map (
            O => \N__4947\,
            I => \N__4944\
        );

    \I__772\ : Span4Mux_h
    port map (
            O => \N__4944\,
            I => \N__4941\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__4941\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__770\ : CascadeMux
    port map (
            O => \N__4938\,
            I => \U712_CHIP_RAM.REFRESH_RST_cascade_\
        );

    \I__769\ : InMux
    port map (
            O => \N__4935\,
            I => \N__4931\
        );

    \I__768\ : InMux
    port map (
            O => \N__4934\,
            I => \N__4928\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4931\,
            I => \U712_REG_SM.N_338\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4928\,
            I => \U712_REG_SM.N_338\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__4923\,
            I => \U712_REG_SM.N_338_cascade_\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__4920\,
            I => \U712_REG_SM.N_354_cascade_\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__4917\,
            I => \N__4914\
        );

    \I__762\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4911\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4911\,
            I => \N__4908\
        );

    \I__760\ : Span4Mux_v
    port map (
            O => \N__4908\,
            I => \N__4905\
        );

    \I__759\ : Sp12to4
    port map (
            O => \N__4905\,
            I => \N__4902\
        );

    \I__758\ : Span12Mux_h
    port map (
            O => \N__4902\,
            I => \N__4899\
        );

    \I__757\ : Span12Mux_v
    port map (
            O => \N__4899\,
            I => \N__4896\
        );

    \I__756\ : Odrv12
    port map (
            O => \N__4896\,
            I => \REGSPACEn_c\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__4893\,
            I => \N__4889\
        );

    \I__754\ : InMux
    port map (
            O => \N__4892\,
            I => \N__4885\
        );

    \I__753\ : InMux
    port map (
            O => \N__4889\,
            I => \N__4880\
        );

    \I__752\ : InMux
    port map (
            O => \N__4888\,
            I => \N__4880\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4885\,
            I => \N__4877\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__4880\,
            I => \N__4874\
        );

    \I__749\ : Span4Mux_v
    port map (
            O => \N__4877\,
            I => \N__4871\
        );

    \I__748\ : Span12Mux_v
    port map (
            O => \N__4874\,
            I => \N__4868\
        );

    \I__747\ : Sp12to4
    port map (
            O => \N__4871\,
            I => \N__4865\
        );

    \I__746\ : Span12Mux_h
    port map (
            O => \N__4868\,
            I => \N__4862\
        );

    \I__745\ : Span12Mux_h
    port map (
            O => \N__4865\,
            I => \N__4859\
        );

    \I__744\ : Span12Mux_v
    port map (
            O => \N__4862\,
            I => \N__4856\
        );

    \I__743\ : Span12Mux_v
    port map (
            O => \N__4859\,
            I => \N__4853\
        );

    \I__742\ : Odrv12
    port map (
            O => \N__4856\,
            I => \CASUn_c\
        );

    \I__741\ : Odrv12
    port map (
            O => \N__4853\,
            I => \CASUn_c\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__4848\,
            I => \N__4845\
        );

    \I__739\ : InMux
    port map (
            O => \N__4845\,
            I => \N__4839\
        );

    \I__738\ : InMux
    port map (
            O => \N__4844\,
            I => \N__4839\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__4839\,
            I => \N__4835\
        );

    \I__736\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4832\
        );

    \I__735\ : Span4Mux_v
    port map (
            O => \N__4835\,
            I => \N__4829\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__4832\,
            I => \N__4826\
        );

    \I__733\ : Sp12to4
    port map (
            O => \N__4829\,
            I => \N__4823\
        );

    \I__732\ : Sp12to4
    port map (
            O => \N__4826\,
            I => \N__4820\
        );

    \I__731\ : Span12Mux_h
    port map (
            O => \N__4823\,
            I => \N__4817\
        );

    \I__730\ : Span12Mux_v
    port map (
            O => \N__4820\,
            I => \N__4814\
        );

    \I__729\ : Span12Mux_v
    port map (
            O => \N__4817\,
            I => \N__4809\
        );

    \I__728\ : Span12Mux_h
    port map (
            O => \N__4814\,
            I => \N__4809\
        );

    \I__727\ : Odrv12
    port map (
            O => \N__4809\,
            I => \CASLn_c\
        );

    \I__726\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4803\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4803\,
            I => \U712_REG_SM.N_431\
        );

    \I__724\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4796\
        );

    \I__723\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4793\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4796\,
            I => \U712_REG_SM.N_358\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4793\,
            I => \U712_REG_SM.N_358\
        );

    \I__720\ : InMux
    port map (
            O => \N__4788\,
            I => \N__4783\
        );

    \I__719\ : InMux
    port map (
            O => \N__4787\,
            I => \N__4780\
        );

    \I__718\ : InMux
    port map (
            O => \N__4786\,
            I => \N__4777\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4783\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4780\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4777\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__4770\,
            I => \U712_CHIP_RAM.N_341_cascade_\
        );

    \I__713\ : InMux
    port map (
            O => \N__4767\,
            I => \N__4763\
        );

    \I__712\ : InMux
    port map (
            O => \N__4766\,
            I => \N__4760\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__4763\,
            I => \U712_CHIP_RAM.N_560\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4760\,
            I => \U712_CHIP_RAM.N_560\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__4755\,
            I => \U712_CHIP_RAM.N_450_cascade_\
        );

    \I__708\ : CascadeMux
    port map (
            O => \N__4752\,
            I => \U712_CHIP_RAM.N_326_cascade_\
        );

    \I__707\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4743\
        );

    \I__706\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4743\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__4743\,
            I => \U712_CHIP_RAM.N_326\
        );

    \I__704\ : IoInMux
    port map (
            O => \N__4740\,
            I => \N__4737\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4737\,
            I => \N__4734\
        );

    \I__702\ : Span4Mux_s3_v
    port map (
            O => \N__4734\,
            I => \N__4731\
        );

    \I__701\ : Span4Mux_h
    port map (
            O => \N__4731\,
            I => \N__4724\
        );

    \I__700\ : InMux
    port map (
            O => \N__4730\,
            I => \N__4719\
        );

    \I__699\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4719\
        );

    \I__698\ : InMux
    port map (
            O => \N__4728\,
            I => \N__4714\
        );

    \I__697\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4714\
        );

    \I__696\ : Sp12to4
    port map (
            O => \N__4724\,
            I => \N__4711\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4719\,
            I => \N__4708\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4714\,
            I => \N__4705\
        );

    \I__693\ : Span12Mux_v
    port map (
            O => \N__4711\,
            I => \N__4701\
        );

    \I__692\ : Span4Mux_v
    port map (
            O => \N__4708\,
            I => \N__4696\
        );

    \I__691\ : Span4Mux_v
    port map (
            O => \N__4705\,
            I => \N__4696\
        );

    \I__690\ : InMux
    port map (
            O => \N__4704\,
            I => \N__4693\
        );

    \I__689\ : Odrv12
    port map (
            O => \N__4701\,
            I => \DBENn_c\
        );

    \I__688\ : Odrv4
    port map (
            O => \N__4696\,
            I => \DBENn_c\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__4693\,
            I => \DBENn_c\
        );

    \I__686\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4682\
        );

    \I__685\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4679\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__4682\,
            I => \U712_CHIP_RAM.N_450\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4679\,
            I => \U712_CHIP_RAM.N_450\
        );

    \I__682\ : InMux
    port map (
            O => \N__4674\,
            I => \N__4670\
        );

    \I__681\ : InMux
    port map (
            O => \N__4673\,
            I => \N__4667\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__4670\,
            I => \N__4664\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__4667\,
            I => \N__4661\
        );

    \I__678\ : Span4Mux_v
    port map (
            O => \N__4664\,
            I => \N__4658\
        );

    \I__677\ : Span4Mux_v
    port map (
            O => \N__4661\,
            I => \N__4655\
        );

    \I__676\ : Sp12to4
    port map (
            O => \N__4658\,
            I => \N__4650\
        );

    \I__675\ : Sp12to4
    port map (
            O => \N__4655\,
            I => \N__4650\
        );

    \I__674\ : Span12Mux_h
    port map (
            O => \N__4650\,
            I => \N__4647\
        );

    \I__673\ : Span12Mux_v
    port map (
            O => \N__4647\,
            I => \N__4644\
        );

    \I__672\ : Odrv12
    port map (
            O => \N__4644\,
            I => \AWEn_c\
        );

    \I__671\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4637\
        );

    \I__670\ : InMux
    port map (
            O => \N__4640\,
            I => \N__4634\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__4637\,
            I => \N__4627\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4634\,
            I => \N__4627\
        );

    \I__667\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4622\
        );

    \I__666\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4622\
        );

    \I__665\ : Span4Mux_v
    port map (
            O => \N__4627\,
            I => \N__4617\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4622\,
            I => \N__4617\
        );

    \I__663\ : Odrv4
    port map (
            O => \N__4617\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__662\ : CEMux
    port map (
            O => \N__4614\,
            I => \N__4611\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4611\,
            I => \N__4608\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__4608\,
            I => \U712_CHIP_RAM.N_450_0\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__4605\,
            I => \N__4601\
        );

    \I__658\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4596\
        );

    \I__657\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4596\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__4596\,
            I => \U712_CHIP_RAM.DMA_CYCLE_7\
        );

    \I__655\ : InMux
    port map (
            O => \N__4593\,
            I => \N__4590\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4590\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a3_0\
        );

    \I__653\ : CascadeMux
    port map (
            O => \N__4587\,
            I => \U712_CHIP_RAM.N_332_cascade_\
        );

    \I__652\ : InMux
    port map (
            O => \N__4584\,
            I => \N__4578\
        );

    \I__651\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4575\
        );

    \I__650\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4570\
        );

    \I__649\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4570\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4578\,
            I => \U712_CHIP_RAM.N_493\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__4575\,
            I => \U712_CHIP_RAM.N_493\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__4570\,
            I => \U712_CHIP_RAM.N_493\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__4563\,
            I => \N__4560\
        );

    \I__644\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4556\
        );

    \I__643\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4551\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__4556\,
            I => \N__4548\
        );

    \I__641\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4545\
        );

    \I__640\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4542\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4551\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__638\ : Odrv4
    port map (
            O => \N__4548\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4545\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__4542\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__635\ : InMux
    port map (
            O => \N__4533\,
            I => \N__4528\
        );

    \I__634\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4525\
        );

    \I__633\ : InMux
    port map (
            O => \N__4531\,
            I => \N__4522\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__4528\,
            I => \N__4517\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4525\,
            I => \N__4517\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4522\,
            I => \U712_CHIP_RAM.N_351\
        );

    \I__629\ : Odrv4
    port map (
            O => \N__4517\,
            I => \U712_CHIP_RAM.N_351\
        );

    \I__628\ : CascadeMux
    port map (
            O => \N__4512\,
            I => \U712_CHIP_RAM.N_351_cascade_\
        );

    \I__627\ : InMux
    port map (
            O => \N__4509\,
            I => \N__4504\
        );

    \I__626\ : InMux
    port map (
            O => \N__4508\,
            I => \N__4501\
        );

    \I__625\ : InMux
    port map (
            O => \N__4507\,
            I => \N__4498\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__4504\,
            I => \N__4487\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__4501\,
            I => \N__4487\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__4498\,
            I => \N__4487\
        );

    \I__621\ : InMux
    port map (
            O => \N__4497\,
            I => \N__4478\
        );

    \I__620\ : InMux
    port map (
            O => \N__4496\,
            I => \N__4478\
        );

    \I__619\ : InMux
    port map (
            O => \N__4495\,
            I => \N__4478\
        );

    \I__618\ : InMux
    port map (
            O => \N__4494\,
            I => \N__4478\
        );

    \I__617\ : Odrv4
    port map (
            O => \N__4487\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4478\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__615\ : InMux
    port map (
            O => \N__4473\,
            I => \N__4470\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__4470\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_o2_1\
        );

    \I__613\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4464\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4464\,
            I => \N__4461\
        );

    \I__611\ : Odrv4
    port map (
            O => \N__4461\,
            I => \U712_CHIP_RAM.N_402\
        );

    \I__610\ : InMux
    port map (
            O => \N__4458\,
            I => \N__4455\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__4455\,
            I => \U712_CHIP_RAM.N_341\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__4452\,
            I => \U712_CHIP_RAM.N_471_cascade_\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__4449\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0_cascade_\
        );

    \I__606\ : IoInMux
    port map (
            O => \N__4446\,
            I => \N__4443\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4443\,
            I => \N__4440\
        );

    \I__604\ : Span12Mux_s6_h
    port map (
            O => \N__4440\,
            I => \N__4437\
        );

    \I__603\ : Span12Mux_h
    port map (
            O => \N__4437\,
            I => \N__4433\
        );

    \I__602\ : InMux
    port map (
            O => \N__4436\,
            I => \N__4430\
        );

    \I__601\ : Odrv12
    port map (
            O => \N__4433\,
            I => \CLK_EN_c\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__4430\,
            I => \CLK_EN_c\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__4425\,
            I => \U712_CHIP_RAM.N_447_cascade_\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__4422\,
            I => \N__4416\
        );

    \I__597\ : InMux
    port map (
            O => \N__4421\,
            I => \N__4413\
        );

    \I__596\ : InMux
    port map (
            O => \N__4420\,
            I => \N__4410\
        );

    \I__595\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4407\
        );

    \I__594\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4404\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4413\,
            I => \N__4401\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4410\,
            I => \U712_CHIP_RAM.N_333\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4407\,
            I => \U712_CHIP_RAM.N_333\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__4404\,
            I => \U712_CHIP_RAM.N_333\
        );

    \I__589\ : Odrv4
    port map (
            O => \N__4401\,
            I => \U712_CHIP_RAM.N_333\
        );

    \I__588\ : InMux
    port map (
            O => \N__4392\,
            I => \N__4385\
        );

    \I__587\ : InMux
    port map (
            O => \N__4391\,
            I => \N__4385\
        );

    \I__586\ : InMux
    port map (
            O => \N__4390\,
            I => \N__4382\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__4385\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4382\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__4377\,
            I => \N__4374\
        );

    \I__582\ : InMux
    port map (
            O => \N__4374\,
            I => \N__4367\
        );

    \I__581\ : InMux
    port map (
            O => \N__4373\,
            I => \N__4367\
        );

    \I__580\ : InMux
    port map (
            O => \N__4372\,
            I => \N__4364\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__4367\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4364\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__4359\,
            I => \N__4355\
        );

    \I__576\ : CascadeMux
    port map (
            O => \N__4358\,
            I => \N__4351\
        );

    \I__575\ : InMux
    port map (
            O => \N__4355\,
            I => \N__4346\
        );

    \I__574\ : InMux
    port map (
            O => \N__4354\,
            I => \N__4346\
        );

    \I__573\ : InMux
    port map (
            O => \N__4351\,
            I => \N__4343\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4346\,
            I => \N__4338\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4343\,
            I => \N__4338\
        );

    \I__570\ : Odrv4
    port map (
            O => \N__4338\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__569\ : CascadeMux
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__568\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4328\
        );

    \I__567\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4325\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4328\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__4325\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__4320\,
            I => \U712_CHIP_RAM.N_330_cascade_\
        );

    \I__563\ : CascadeMux
    port map (
            O => \N__4317\,
            I => \N__4314\
        );

    \I__562\ : InMux
    port map (
            O => \N__4314\,
            I => \N__4311\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__4311\,
            I => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\
        );

    \I__560\ : InMux
    port map (
            O => \N__4308\,
            I => \N__4305\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4305\,
            I => \N__4301\
        );

    \I__558\ : InMux
    port map (
            O => \N__4304\,
            I => \N__4298\
        );

    \I__557\ : Span4Mux_h
    port map (
            O => \N__4301\,
            I => \N__4295\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4298\,
            I => \CPU_TACKm\
        );

    \I__555\ : Odrv4
    port map (
            O => \N__4295\,
            I => \CPU_TACKm\
        );

    \I__554\ : CascadeMux
    port map (
            O => \N__4290\,
            I => \U712_CHIP_RAM.N_554_cascade_\
        );

    \I__553\ : InMux
    port map (
            O => \N__4287\,
            I => \N__4284\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__4284\,
            I => \U712_CHIP_RAM.N_565\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__4281\,
            I => \U712_CHIP_RAM.N_565_cascade_\
        );

    \I__550\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4275\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4275\,
            I => \U712_CHIP_RAM.N_563\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__4272\,
            I => \U712_CHIP_RAM.N_445_cascade_\
        );

    \I__547\ : InMux
    port map (
            O => \N__4269\,
            I => \N__4266\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__4266\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_a3_2_1\
        );

    \I__545\ : CascadeMux
    port map (
            O => \N__4263\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_1_1_cascade_\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__4260\,
            I => \U712_CHIP_RAM.N_333_cascade_\
        );

    \I__543\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4253\
        );

    \I__542\ : InMux
    port map (
            O => \N__4256\,
            I => \N__4250\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__4253\,
            I => \U712_CHIP_RAM.N_564\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4250\,
            I => \U712_CHIP_RAM.N_564\
        );

    \I__539\ : IoInMux
    port map (
            O => \N__4245\,
            I => \N__4242\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4242\,
            I => \N__4239\
        );

    \I__537\ : Span4Mux_s0_v
    port map (
            O => \N__4239\,
            I => \N__4236\
        );

    \I__536\ : Span4Mux_h
    port map (
            O => \N__4236\,
            I => \N__4233\
        );

    \I__535\ : Span4Mux_v
    port map (
            O => \N__4233\,
            I => \N__4230\
        );

    \I__534\ : Span4Mux_v
    port map (
            O => \N__4230\,
            I => \N__4227\
        );

    \I__533\ : Sp12to4
    port map (
            O => \N__4227\,
            I => \N__4224\
        );

    \I__532\ : Span12Mux_h
    port map (
            O => \N__4224\,
            I => \N__4221\
        );

    \I__531\ : Odrv12
    port map (
            O => \N__4221\,
            I => \DRDENn_c\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__4218\,
            I => \U712_REG_SM.N_343_cascade_\
        );

    \I__529\ : CascadeMux
    port map (
            O => \N__4215\,
            I => \U712_REG_SM.N_358_cascade_\
        );

    \I__528\ : InMux
    port map (
            O => \N__4212\,
            I => \N__4209\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4209\,
            I => \N__4203\
        );

    \I__526\ : InMux
    port map (
            O => \N__4208\,
            I => \N__4196\
        );

    \I__525\ : InMux
    port map (
            O => \N__4207\,
            I => \N__4196\
        );

    \I__524\ : InMux
    port map (
            O => \N__4206\,
            I => \N__4196\
        );

    \I__523\ : Odrv12
    port map (
            O => \N__4203\,
            I => \REG_CYCLEm\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4196\,
            I => \REG_CYCLEm\
        );

    \I__521\ : CascadeMux
    port map (
            O => \N__4191\,
            I => \N__4188\
        );

    \I__520\ : InMux
    port map (
            O => \N__4188\,
            I => \N__4184\
        );

    \I__519\ : InMux
    port map (
            O => \N__4187\,
            I => \N__4181\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4184\,
            I => \REG_TACK\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4181\,
            I => \REG_TACK\
        );

    \I__516\ : CascadeMux
    port map (
            O => \N__4176\,
            I => \U712_CHIP_RAM.N_563_cascade_\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__4173\,
            I => \U712_CHIP_RAM.N_215_cascade_\
        );

    \I__514\ : InMux
    port map (
            O => \N__4170\,
            I => \N__4167\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4167\,
            I => \N__4164\
        );

    \I__512\ : Span4Mux_h
    port map (
            O => \N__4164\,
            I => \N__4161\
        );

    \I__511\ : Sp12to4
    port map (
            O => \N__4161\,
            I => \N__4158\
        );

    \I__510\ : Span12Mux_v
    port map (
            O => \N__4158\,
            I => \N__4155\
        );

    \I__509\ : Odrv12
    port map (
            O => \N__4155\,
            I => \A_c_18\
        );

    \I__508\ : CascadeMux
    port map (
            O => \N__4152\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_7_cascade_\
        );

    \I__507\ : InMux
    port map (
            O => \N__4149\,
            I => \N__4146\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4146\,
            I => \N__4143\
        );

    \I__505\ : Sp12to4
    port map (
            O => \N__4143\,
            I => \N__4140\
        );

    \I__504\ : Span12Mux_v
    port map (
            O => \N__4140\,
            I => \N__4137\
        );

    \I__503\ : Span12Mux_h
    port map (
            O => \N__4137\,
            I => \N__4134\
        );

    \I__502\ : Odrv12
    port map (
            O => \N__4134\,
            I => \A_c_16\
        );

    \I__501\ : InMux
    port map (
            O => \N__4131\,
            I => \N__4125\
        );

    \I__500\ : InMux
    port map (
            O => \N__4130\,
            I => \N__4125\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4125\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_ac0_7_0\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__4122\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6_cascade_\
        );

    \I__497\ : InMux
    port map (
            O => \N__4119\,
            I => \N__4116\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__4116\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6\
        );

    \I__495\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4110\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4110\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0\
        );

    \I__493\ : IoInMux
    port map (
            O => \N__4107\,
            I => \N__4104\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__4104\,
            I => \N__4101\
        );

    \I__491\ : Span4Mux_s1_v
    port map (
            O => \N__4101\,
            I => \N__4098\
        );

    \I__490\ : Span4Mux_v
    port map (
            O => \N__4098\,
            I => \N__4095\
        );

    \I__489\ : Span4Mux_v
    port map (
            O => \N__4095\,
            I => \N__4092\
        );

    \I__488\ : Span4Mux_v
    port map (
            O => \N__4092\,
            I => \N__4087\
        );

    \I__487\ : InMux
    port map (
            O => \N__4091\,
            I => \N__4084\
        );

    \I__486\ : InMux
    port map (
            O => \N__4090\,
            I => \N__4081\
        );

    \I__485\ : Odrv4
    port map (
            O => \N__4087\,
            I => \DBDIR_c\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4084\,
            I => \DBDIR_c\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__4081\,
            I => \DBDIR_c\
        );

    \I__482\ : IoInMux
    port map (
            O => \N__4074\,
            I => \N__4071\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4071\,
            I => \N__4068\
        );

    \I__480\ : Span4Mux_s2_h
    port map (
            O => \N__4068\,
            I => \N__4065\
        );

    \I__479\ : Span4Mux_v
    port map (
            O => \N__4065\,
            I => \N__4062\
        );

    \I__478\ : Sp12to4
    port map (
            O => \N__4062\,
            I => \N__4059\
        );

    \I__477\ : Span12Mux_s11_h
    port map (
            O => \N__4059\,
            I => \N__4056\
        );

    \I__476\ : Span12Mux_v
    port map (
            O => \N__4056\,
            I => \N__4053\
        );

    \I__475\ : Odrv12
    port map (
            O => \N__4053\,
            I => \DRDDIR_i_0\
        );

    \I__474\ : InMux
    port map (
            O => \N__4050\,
            I => \N__4046\
        );

    \I__473\ : InMux
    port map (
            O => \N__4049\,
            I => \N__4043\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4046\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4043\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0\
        );

    \I__470\ : CascadeMux
    port map (
            O => \N__4038\,
            I => \U712_BYTE_ENABLE.N_459_cascade_\
        );

    \I__469\ : InMux
    port map (
            O => \N__4035\,
            I => \N__4032\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4032\,
            I => \U712_BYTE_ENABLE.N_352\
        );

    \I__467\ : IoInMux
    port map (
            O => \N__4029\,
            I => \N__4026\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4026\,
            I => \N__4023\
        );

    \I__465\ : Span12Mux_s4_v
    port map (
            O => \N__4023\,
            I => \N__4020\
        );

    \I__464\ : Odrv12
    port map (
            O => \N__4020\,
            I => \N_47_i\
        );

    \I__463\ : CascadeMux
    port map (
            O => \N__4017\,
            I => \N__4012\
        );

    \I__462\ : InMux
    port map (
            O => \N__4016\,
            I => \N__4009\
        );

    \I__461\ : InMux
    port map (
            O => \N__4015\,
            I => \N__4004\
        );

    \I__460\ : InMux
    port map (
            O => \N__4012\,
            I => \N__4004\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__4009\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4004\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__3999\,
            I => \N__3996\
        );

    \I__456\ : InMux
    port map (
            O => \N__3996\,
            I => \N__3992\
        );

    \I__455\ : InMux
    port map (
            O => \N__3995\,
            I => \N__3989\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__3992\,
            I => \N__3984\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3989\,
            I => \N__3984\
        );

    \I__452\ : Odrv4
    port map (
            O => \N__3984\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__451\ : CascadeMux
    port map (
            O => \N__3981\,
            I => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\
        );

    \I__450\ : InMux
    port map (
            O => \N__3978\,
            I => \N__3973\
        );

    \I__449\ : InMux
    port map (
            O => \N__3977\,
            I => \N__3970\
        );

    \I__448\ : InMux
    port map (
            O => \N__3976\,
            I => \N__3967\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3973\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__3970\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3967\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__3960\,
            I => \U712_CYCLE_TERM.N_362_i_0_en_cascade_\
        );

    \I__443\ : CEMux
    port map (
            O => \N__3957\,
            I => \N__3954\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__3954\,
            I => \N__3951\
        );

    \I__441\ : Odrv4
    port map (
            O => \N__3951\,
            I => \U712_CYCLE_TERM.N_362_i_0_en_0\
        );

    \I__440\ : IoInMux
    port map (
            O => \N__3948\,
            I => \N__3945\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3945\,
            I => \N__3942\
        );

    \I__438\ : Span12Mux_s10_v
    port map (
            O => \N__3942\,
            I => \N__3939\
        );

    \I__437\ : Odrv12
    port map (
            O => \N__3939\,
            I => \VBENn_c\
        );

    \I__436\ : InMux
    port map (
            O => \N__3936\,
            I => \N__3932\
        );

    \I__435\ : InMux
    port map (
            O => \N__3935\,
            I => \N__3929\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3932\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3929\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__432\ : InMux
    port map (
            O => \N__3924\,
            I => \N__3920\
        );

    \I__431\ : InMux
    port map (
            O => \N__3923\,
            I => \N__3917\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3920\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3917\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__428\ : CascadeMux
    port map (
            O => \N__3912\,
            I => \N__3908\
        );

    \I__427\ : InMux
    port map (
            O => \N__3911\,
            I => \N__3905\
        );

    \I__426\ : InMux
    port map (
            O => \N__3908\,
            I => \N__3902\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3905\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3902\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__423\ : InMux
    port map (
            O => \N__3897\,
            I => \N__3893\
        );

    \I__422\ : InMux
    port map (
            O => \N__3896\,
            I => \N__3890\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3893\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3890\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__419\ : InMux
    port map (
            O => \N__3885\,
            I => \N__3881\
        );

    \I__418\ : InMux
    port map (
            O => \N__3884\,
            I => \N__3878\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3881\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3878\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__415\ : InMux
    port map (
            O => \N__3873\,
            I => \N__3869\
        );

    \I__414\ : InMux
    port map (
            O => \N__3872\,
            I => \N__3866\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__3869\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__3866\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__3861\,
            I => \N__3858\
        );

    \I__410\ : InMux
    port map (
            O => \N__3858\,
            I => \N__3854\
        );

    \I__409\ : InMux
    port map (
            O => \N__3857\,
            I => \N__3850\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3854\,
            I => \N__3847\
        );

    \I__407\ : InMux
    port map (
            O => \N__3853\,
            I => \N__3844\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3850\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__405\ : Odrv12
    port map (
            O => \N__3847\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__3844\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__403\ : IoInMux
    port map (
            O => \N__3837\,
            I => \N__3834\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3834\,
            I => \N__3831\
        );

    \I__401\ : IoSpan4Mux
    port map (
            O => \N__3831\,
            I => \N__3828\
        );

    \I__400\ : Span4Mux_s3_h
    port map (
            O => \N__3828\,
            I => \N__3825\
        );

    \I__399\ : Span4Mux_h
    port map (
            O => \N__3825\,
            I => \N__3822\
        );

    \I__398\ : Sp12to4
    port map (
            O => \N__3822\,
            I => \N__3819\
        );

    \I__397\ : Span12Mux_v
    port map (
            O => \N__3819\,
            I => \N__3815\
        );

    \I__396\ : InMux
    port map (
            O => \N__3818\,
            I => \N__3812\
        );

    \I__395\ : Odrv12
    port map (
            O => \N__3815\,
            I => \TACK_OUTn\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3812\,
            I => \TACK_OUTn\
        );

    \I__393\ : InMux
    port map (
            O => \N__3807\,
            I => \N__3803\
        );

    \I__392\ : InMux
    port map (
            O => \N__3806\,
            I => \N__3800\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__3803\,
            I => \N__3797\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3800\,
            I => \N__3794\
        );

    \I__389\ : Odrv4
    port map (
            O => \N__3797\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__388\ : Odrv4
    port map (
            O => \N__3794\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__387\ : InMux
    port map (
            O => \N__3789\,
            I => \N__3786\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__3786\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\
        );

    \I__385\ : InMux
    port map (
            O => \N__3783\,
            I => \N__3780\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3780\,
            I => \N__3774\
        );

    \I__383\ : InMux
    port map (
            O => \N__3779\,
            I => \N__3767\
        );

    \I__382\ : InMux
    port map (
            O => \N__3778\,
            I => \N__3767\
        );

    \I__381\ : InMux
    port map (
            O => \N__3777\,
            I => \N__3767\
        );

    \I__380\ : Span4Mux_h
    port map (
            O => \N__3774\,
            I => \N__3762\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__3767\,
            I => \N__3762\
        );

    \I__378\ : Span4Mux_v
    port map (
            O => \N__3762\,
            I => \N__3759\
        );

    \I__377\ : Span4Mux_h
    port map (
            O => \N__3759\,
            I => \N__3756\
        );

    \I__376\ : Span4Mux_v
    port map (
            O => \N__3756\,
            I => \N__3753\
        );

    \I__375\ : Span4Mux_v
    port map (
            O => \N__3753\,
            I => \N__3750\
        );

    \I__374\ : Odrv4
    port map (
            O => \N__3750\,
            I => \CLK40_OUT_i\
        );

    \I__373\ : InMux
    port map (
            O => \N__3747\,
            I => \N__3735\
        );

    \I__372\ : InMux
    port map (
            O => \N__3746\,
            I => \N__3735\
        );

    \I__371\ : InMux
    port map (
            O => \N__3745\,
            I => \N__3735\
        );

    \I__370\ : InMux
    port map (
            O => \N__3744\,
            I => \N__3735\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__3735\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__368\ : InMux
    port map (
            O => \N__3732\,
            I => \N__3729\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__3729\,
            I => \U712_BYTE_ENABLE.N_455\
        );

    \I__366\ : InMux
    port map (
            O => \N__3726\,
            I => \N__3720\
        );

    \I__365\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3720\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3720\,
            I => \N__3717\
        );

    \I__363\ : Span4Mux_v
    port map (
            O => \N__3717\,
            I => \N__3714\
        );

    \I__362\ : Sp12to4
    port map (
            O => \N__3714\,
            I => \N__3711\
        );

    \I__361\ : Span12Mux_h
    port map (
            O => \N__3711\,
            I => \N__3708\
        );

    \I__360\ : Span12Mux_v
    port map (
            O => \N__3708\,
            I => \N__3705\
        );

    \I__359\ : Odrv12
    port map (
            O => \N__3705\,
            I => \SIZ_c_1\
        );

    \I__358\ : CascadeMux
    port map (
            O => \N__3702\,
            I => \U712_BYTE_ENABLE.N_352_cascade_\
        );

    \I__357\ : IoInMux
    port map (
            O => \N__3699\,
            I => \N__3696\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__3696\,
            I => \N__3693\
        );

    \I__355\ : IoSpan4Mux
    port map (
            O => \N__3693\,
            I => \N__3690\
        );

    \I__354\ : Span4Mux_s3_v
    port map (
            O => \N__3690\,
            I => \N__3687\
        );

    \I__353\ : Sp12to4
    port map (
            O => \N__3687\,
            I => \N__3684\
        );

    \I__352\ : Span12Mux_v
    port map (
            O => \N__3684\,
            I => \N__3681\
        );

    \I__351\ : Span12Mux_h
    port map (
            O => \N__3681\,
            I => \N__3678\
        );

    \I__350\ : Odrv12
    port map (
            O => \N__3678\,
            I => \N_49_i\
        );

    \I__349\ : IoInMux
    port map (
            O => \N__3675\,
            I => \N__3672\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3672\,
            I => \N__3669\
        );

    \I__347\ : Span12Mux_s5_h
    port map (
            O => \N__3669\,
            I => \N__3666\
        );

    \I__346\ : Odrv12
    port map (
            O => \N__3666\,
            I => \CLK40_OUT_i_i\
        );

    \I__345\ : InMux
    port map (
            O => \N__3663\,
            I => \N__3657\
        );

    \I__344\ : InMux
    port map (
            O => \N__3662\,
            I => \N__3657\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3657\,
            I => \N__3654\
        );

    \I__342\ : Sp12to4
    port map (
            O => \N__3654\,
            I => \N__3651\
        );

    \I__341\ : Span12Mux_v
    port map (
            O => \N__3651\,
            I => \N__3648\
        );

    \I__340\ : Odrv12
    port map (
            O => \N__3648\,
            I => \A_c_1\
        );

    \I__339\ : InMux
    port map (
            O => \N__3645\,
            I => \N__3642\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__3642\,
            I => \N__3639\
        );

    \I__337\ : Odrv4
    port map (
            O => \N__3639\,
            I => \U712_BYTE_ENABLE.N_457\
        );

    \I__336\ : InMux
    port map (
            O => \N__3636\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__335\ : InMux
    port map (
            O => \N__3633\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__334\ : InMux
    port map (
            O => \N__3630\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__333\ : InMux
    port map (
            O => \N__3627\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__332\ : InMux
    port map (
            O => \N__3624\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__331\ : ClkMux
    port map (
            O => \N__3621\,
            I => \N__3618\
        );

    \I__330\ : GlobalMux
    port map (
            O => \N__3618\,
            I => \N__3615\
        );

    \I__329\ : gio2CtrlBuf
    port map (
            O => \N__3615\,
            I => \C1_c_g\
        );

    \I__328\ : InMux
    port map (
            O => \N__3612\,
            I => \N__3609\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__3609\,
            I => \TACK_EN_i_ess\
        );

    \I__326\ : IoInMux
    port map (
            O => \N__3606\,
            I => \N__3603\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__3603\,
            I => \N__3600\
        );

    \I__324\ : Span12Mux_s5_h
    port map (
            O => \N__3600\,
            I => \N__3597\
        );

    \I__323\ : Span12Mux_v
    port map (
            O => \N__3597\,
            I => \N__3594\
        );

    \I__322\ : Odrv12
    port map (
            O => \N__3594\,
            I => \N_888_i\
        );

    \I__321\ : CascadeMux
    port map (
            O => \N__3591\,
            I => \U712_BYTE_ENABLE.N_451_cascade_\
        );

    \I__320\ : IoInMux
    port map (
            O => \N__3588\,
            I => \N__3585\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__3585\,
            I => \N__3582\
        );

    \I__318\ : Span4Mux_s2_h
    port map (
            O => \N__3582\,
            I => \N__3579\
        );

    \I__317\ : Span4Mux_h
    port map (
            O => \N__3579\,
            I => \N__3576\
        );

    \I__316\ : Sp12to4
    port map (
            O => \N__3576\,
            I => \N__3573\
        );

    \I__315\ : Span12Mux_v
    port map (
            O => \N__3573\,
            I => \N__3570\
        );

    \I__314\ : Span12Mux_h
    port map (
            O => \N__3570\,
            I => \N__3567\
        );

    \I__313\ : Odrv12
    port map (
            O => \N__3567\,
            I => \N_48_i\
        );

    \I__312\ : IoInMux
    port map (
            O => \N__3564\,
            I => \N__3561\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__3561\,
            I => \N__3558\
        );

    \I__310\ : Span4Mux_s2_v
    port map (
            O => \N__3558\,
            I => \N__3555\
        );

    \I__309\ : Span4Mux_v
    port map (
            O => \N__3555\,
            I => \N__3552\
        );

    \I__308\ : Odrv4
    port map (
            O => \N__3552\,
            I => \CLK80_OUT_i_i\
        );

    \I__307\ : InMux
    port map (
            O => \N__3549\,
            I => \bfn_7_7_0_\
        );

    \I__306\ : InMux
    port map (
            O => \N__3546\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__305\ : InMux
    port map (
            O => \N__3543\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__304\ : IoInMux
    port map (
            O => \N__3540\,
            I => \N__3537\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__3537\,
            I => \N__3534\
        );

    \I__302\ : Span4Mux_s0_v
    port map (
            O => \N__3534\,
            I => \N__3531\
        );

    \I__301\ : Span4Mux_v
    port map (
            O => \N__3531\,
            I => \N__3528\
        );

    \I__300\ : Sp12to4
    port map (
            O => \N__3528\,
            I => \N__3525\
        );

    \I__299\ : Span12Mux_h
    port map (
            O => \N__3525\,
            I => \N__3522\
        );

    \I__298\ : Span12Mux_v
    port map (
            O => \N__3522\,
            I => \N__3519\
        );

    \I__297\ : Odrv12
    port map (
            O => \N__3519\,
            I => \CLK40_IN_c\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7437\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5888\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_3_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9162\,
            lcout => \CLK80_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3897\,
            in2 => \_gnd_net_\,
            in3 => \N__3549\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__3621\,
            ce => 'H',
            sr => \N__4953\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3924\,
            in2 => \_gnd_net_\,
            in3 => \N__3546\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__3621\,
            ce => 'H',
            sr => \N__4953\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3936\,
            in2 => \_gnd_net_\,
            in3 => \N__3543\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__3621\,
            ce => 'H',
            sr => \N__4953\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5459\,
            in2 => \_gnd_net_\,
            in3 => \N__3636\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__3621\,
            ce => 'H',
            sr => \N__4953\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3911\,
            in2 => \_gnd_net_\,
            in3 => \N__3633\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__3621\,
            ce => 'H',
            sr => \N__4953\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3873\,
            in2 => \_gnd_net_\,
            in3 => \N__3630\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__3621\,
            ce => 'H',
            sr => \N__4953\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3885\,
            in2 => \_gnd_net_\,
            in3 => \N__3627\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__3621\,
            ce => 'H',
            sr => \N__4953\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5429\,
            in2 => \_gnd_net_\,
            in3 => \N__3624\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3621\,
            ce => 'H',
            sr => \N__4953\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__3978\,
            in1 => \N__7520\,
            in2 => \_gnd_net_\,
            in3 => \N__4016\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9157\,
            ce => \N__3957\,
            sr => \N__8965\
        );

    \TACKn_obuft_RNO_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3612\,
            lcout => \N_888_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__7374\,
            in1 => \N__3726\,
            in2 => \_gnd_net_\,
            in3 => \N__8155\,
            lcout => \U712_BYTE_ENABLE.N_451\,
            ltout => \U712_BYTE_ENABLE.N_451_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_48_i_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__3645\,
            in1 => \N__6892\,
            in2 => \N__3591\,
            in3 => \N__4049\,
            lcout => \N_48_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_o2_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__6893\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3725\,
            lcout => \U712_BYTE_ENABLE.N_352\,
            ltout => \U712_BYTE_ENABLE.N_352_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_49_i_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__3732\,
            in1 => \N__7058\,
            in2 => \N__3702\,
            in3 => \N__7039\,
            lcout => \N_49_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK40C_obuf_RNO_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3783\,
            lcout => \CLK40_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3662\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8156\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_1_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__3663\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8157\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3807\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9145\,
            ce => 'H',
            sr => \N__8972\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3857\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9145\,
            ce => 'H',
            sr => \N__8972\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3853\,
            in2 => \_gnd_net_\,
            in3 => \N__3806\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__6111\,
            in1 => \_gnd_net_\,
            in2 => \N__4893\,
            in3 => \N__4730\,
            lcout => \U712_BYTE_ENABLE.N_453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_0_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4729\,
            in1 => \N__4888\,
            in2 => \_gnd_net_\,
            in3 => \N__6110\,
            lcout => \U712_BYTE_ENABLE.N_457\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__3935\,
            in1 => \N__3923\,
            in2 => \N__3912\,
            in3 => \N__3896\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3884\,
            in2 => \_gnd_net_\,
            in3 => \N__3872\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110011110100"
        )
    port map (
            in0 => \N__3746\,
            in1 => \N__3818\,
            in2 => \N__3861\,
            in3 => \N__3777\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9153\,
            ce => 'H',
            sr => \N__8951\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__3779\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3745\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9153\,
            ce => 'H',
            sr => \N__8951\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__3789\,
            in1 => \N__4015\,
            in2 => \N__3999\,
            in3 => \N__3744\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9153\,
            ce => 'H',
            sr => \N__8951\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110001000"
        )
    port map (
            in0 => \N__3747\,
            in1 => \N__3778\,
            in2 => \N__4017\,
            in3 => \N__3977\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9153\,
            ce => 'H',
            sr => \N__8951\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__4728\,
            in1 => \_gnd_net_\,
            in2 => \N__4848\,
            in3 => \N__6109\,
            lcout => \U712_BYTE_ENABLE.N_455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6108\,
            in1 => \N__4844\,
            in2 => \_gnd_net_\,
            in3 => \N__4727\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_459_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_47_i_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__7046\,
            in1 => \N__4050\,
            in2 => \N__4038\,
            in3 => \N__4035\,
            lcout => \N_47_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4187\,
            in2 => \_gnd_net_\,
            in3 => \N__4308\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__7503\,
            in1 => \N__3995\,
            in2 => \N__3981\,
            in3 => \N__3976\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_362_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9019\,
            in1 => \_gnd_net_\,
            in2 => \N__3960\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.N_362_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__5400\,
            in1 => \N__7523\,
            in2 => \N__4563\,
            in3 => \N__4507\,
            lcout => \U712_CHIP_RAM.N_492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a3_0_a3_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4212\,
            in2 => \_gnd_net_\,
            in3 => \N__8118\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4532\,
            in1 => \N__5609\,
            in2 => \N__7527\,
            in3 => \N__5700\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_a3_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__5798\,
            in1 => \N__9026\,
            in2 => \N__4359\,
            in3 => \N__5827\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9136\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7743\,
            in1 => \N__8115\,
            in2 => \N__8817\,
            in3 => \N__8241\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__8116\,
            in1 => \N__4170\,
            in2 => \N__4152\,
            in3 => \N__4149\,
            lcout => \U712_CHIP_RAM.N_374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_4_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5797\,
            in2 => \_gnd_net_\,
            in3 => \N__4354\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_ac0_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__4131\,
            in1 => \N__9022\,
            in2 => \N__4377\,
            in3 => \N__5829\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5828\,
            in1 => \N__4130\,
            in2 => \_gnd_net_\,
            in3 => \N__4373\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9023\,
            in2 => \N__4122\,
            in3 => \N__4391\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__4119\,
            in1 => \N__9024\,
            in2 => \N__4335\,
            in3 => \N__4392\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000001"
        )
    port map (
            in0 => \N__4531\,
            in1 => \N__5711\,
            in2 => \N__5613\,
            in3 => \N__4421\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__4113\,
            in1 => \N__4559\,
            in2 => \_gnd_net_\,
            in3 => \N__5186\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9149\,
            ce => 'H',
            sr => \N__8943\
        );

    \U712_CHIP_RAM.DBDIR_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__4673\,
            in1 => \N__4090\,
            in2 => \_gnd_net_\,
            in3 => \N__4686\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9149\,
            ce => 'H',
            sr => \N__8943\
        );

    \U712_BUFFERS.DRDDIR_i_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__4207\,
            in1 => \N__7413\,
            in2 => \N__6097\,
            in3 => \N__4091\,
            lcout => \DRDDIR_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4208\,
            in2 => \_gnd_net_\,
            in3 => \N__6090\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__4934\,
            in1 => \N__7114\,
            in2 => \_gnd_net_\,
            in3 => \N__7149\,
            lcout => \U712_REG_SM.N_343\,
            ltout => \U712_REG_SM.N_343_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5916\,
            in2 => \N__4218\,
            in3 => \N__5952\,
            lcout => \U712_REG_SM.N_358\,
            ltout => \U712_REG_SM.N_358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001010"
        )
    port map (
            in0 => \N__4787\,
            in1 => \N__6966\,
            in2 => \N__4215\,
            in3 => \N__4206\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9154\,
            ce => 'H',
            sr => \N__8936\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__6476\,
            in1 => \N__4786\,
            in2 => \N__6458\,
            in3 => \N__4800\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9158\,
            ce => 'H',
            sr => \N__8931\
        );

    \U712_REG_SM.REG_TACK_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101010000"
        )
    port map (
            in0 => \N__6965\,
            in1 => \N__6454\,
            in2 => \N__4191\,
            in3 => \N__6475\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9158\,
            ce => 'H',
            sr => \N__8931\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIM76F1_1_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5273\,
            in2 => \_gnd_net_\,
            in3 => \N__5608\,
            lcout => \U712_CHIP_RAM.N_563\,
            ltout => \U712_CHIP_RAM.N_563_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__7518\,
            in1 => \N__4640\,
            in2 => \N__4176\,
            in3 => \N__4287\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5243\,
            in2 => \N__4173\,
            in3 => \N__8650\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000011"
        )
    port map (
            in0 => \N__5607\,
            in1 => \N__4509\,
            in2 => \N__4422\,
            in3 => \N__5699\,
            lcout => \U712_CHIP_RAM.N_565\,
            ltout => \U712_CHIP_RAM.N_565_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOF0DC_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__5181\,
            in1 => \N__7519\,
            in2 => \N__4281\,
            in3 => \N__4257\,
            lcout => \U712_CHIP_RAM.N_445\,
            ltout => \U712_CHIP_RAM.N_445_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101100000001"
        )
    port map (
            in0 => \N__5244\,
            in1 => \N__4278\,
            in2 => \N__4272\,
            in3 => \N__7846\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__4533\,
            in1 => \N__4256\,
            in2 => \_gnd_net_\,
            in3 => \N__5178\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__7522\,
            in1 => \N__4269\,
            in2 => \N__4263\,
            in3 => \N__4419\,
            lcout => \U712_CHIP_RAM.N_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5778\,
            in1 => \N__5501\,
            in2 => \_gnd_net_\,
            in3 => \N__5119\,
            lcout => \U712_CHIP_RAM.N_333\,
            ltout => \U712_CHIP_RAM.N_333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__5669\,
            in1 => \_gnd_net_\,
            in2 => \N__4260\,
            in3 => \N__5573\,
            lcout => \U712_CHIP_RAM.N_346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__4581\,
            in1 => \N__5502\,
            in2 => \N__5796\,
            in3 => \N__4508\,
            lcout => \U712_CHIP_RAM.N_564\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5503\,
            in1 => \N__5218\,
            in2 => \N__5802\,
            in3 => \N__4582\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_471_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110101"
        )
    port map (
            in0 => \N__5219\,
            in1 => \_gnd_net_\,
            in2 => \N__4452\,
            in3 => \N__5179\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101011111010"
        )
    port map (
            in0 => \N__4436\,
            in1 => \N__4641\,
            in2 => \N__4449\,
            in3 => \N__5707\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9127\,
            ce => 'H',
            sr => \N__8966\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8117\,
            in1 => \N__4632\,
            in2 => \N__5520\,
            in3 => \N__4583\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_447_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__4633\,
            in1 => \N__5672\,
            in2 => \N__4425\,
            in3 => \N__4420\,
            lcout => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4390\,
            in1 => \N__4372\,
            in2 => \N__4358\,
            in3 => \N__4331\,
            lcout => \U712_CHIP_RAM.N_330\,
            ltout => \U712_CHIP_RAM.N_330_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5574\,
            in2 => \N__4320\,
            in3 => \N__5670\,
            lcout => \U712_CHIP_RAM.N_493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__5130\,
            in1 => \N__4593\,
            in2 => \N__4317\,
            in3 => \N__4304\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9132\,
            ce => 'H',
            sr => \N__8952\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIU9AV6_0_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__4766\,
            in1 => \N__5255\,
            in2 => \N__5133\,
            in3 => \N__5671\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_554_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRDCDD_0_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__9025\,
            in1 => \N__4467\,
            in2 => \N__4290\,
            in3 => \N__5180\,
            lcout => \U712_CHIP_RAM.N_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__5784\,
            in1 => \N__5710\,
            in2 => \N__5603\,
            in3 => \N__5217\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__4494\,
            in1 => \N__5393\,
            in2 => \_gnd_net_\,
            in3 => \N__4554\,
            lcout => \U712_CHIP_RAM.N_332\,
            ltout => \U712_CHIP_RAM.N_332_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__5783\,
            in1 => \N__5576\,
            in2 => \N__4587\,
            in3 => \N__5510\,
            lcout => \U712_CHIP_RAM.N_560\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__4497\,
            in1 => \N__4584\,
            in2 => \N__5519\,
            in3 => \N__5785\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9137\,
            ce => 'H',
            sr => \N__8944\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__5392\,
            in1 => \N__4555\,
            in2 => \_gnd_net_\,
            in3 => \N__4496\,
            lcout => \U712_CHIP_RAM.N_351\,
            ltout => \U712_CHIP_RAM.N_351_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOMFN2_2_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000000000"
        )
    port map (
            in0 => \N__5509\,
            in1 => \N__5586\,
            in2 => \N__4512\,
            in3 => \N__4473\,
            lcout => \U712_CHIP_RAM.N_331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP0891_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001100110"
        )
    port map (
            in0 => \N__5782\,
            in1 => \N__5575\,
            in2 => \_gnd_net_\,
            in3 => \N__4495\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_o2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5207\,
            in2 => \_gnd_net_\,
            in3 => \N__4458\,
            lcout => \U712_CHIP_RAM.N_402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5300\,
            in1 => \N__5937\,
            in2 => \N__6050\,
            in3 => \N__5902\,
            lcout => \U712_CHIP_RAM.N_341\,
            ltout => \U712_CHIP_RAM.N_341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI7Q5U5_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5208\,
            in2 => \N__4770\,
            in3 => \N__5185\,
            lcout => \U712_CHIP_RAM.N_450\,
            ltout => \U712_CHIP_RAM.N_450_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_0_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__4767\,
            in1 => \N__5708\,
            in2 => \N__4755\,
            in3 => \N__5132\,
            lcout => \U712_CHIP_RAM.N_326\,
            ltout => \U712_CHIP_RAM.N_326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__5709\,
            in1 => \N__8076\,
            in2 => \N__4752\,
            in3 => \N__6037\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9147\,
            ce => 'H',
            sr => \N__8937\
        );

    \U712_CHIP_RAM.DMA_CYCLE_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__4749\,
            in1 => \N__6084\,
            in2 => \_gnd_net_\,
            in3 => \N__4604\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9147\,
            ce => 'H',
            sr => \N__8937\
        );

    \U712_CHIP_RAM.DBENn_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101111111001100"
        )
    port map (
            in0 => \N__7752\,
            in1 => \N__4704\,
            in2 => \N__4605\,
            in3 => \N__4748\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9147\,
            ce => 'H',
            sr => \N__8937\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9018\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4685\,
            lcout => \U712_CHIP_RAM.N_450_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001100"
        )
    port map (
            in0 => \N__4674\,
            in1 => \N__5307\,
            in2 => \N__7424\,
            in3 => \N__6053\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9150\,
            ce => \N__4614\,
            sr => \N__8932\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__6052\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5715\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7146\,
            in1 => \N__4935\,
            in2 => \_gnd_net_\,
            in3 => \N__7115\,
            lcout => \U712_REG_SM.N_361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__6435\,
            in1 => \N__6766\,
            in2 => \N__6402\,
            in3 => \N__6722\,
            lcout => \U712_REG_SM.N_338\,
            ltout => \U712_REG_SM.N_338_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__7147\,
            in1 => \N__5989\,
            in2 => \N__4923\,
            in3 => \N__7116\,
            lcout => \U712_REG_SM.N_431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6767\,
            in2 => \_gnd_net_\,
            in3 => \N__6721\,
            lcout => \U712_REG_SM.N_354\,
            ltout => \U712_REG_SM.N_354_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000001"
        )
    port map (
            in0 => \N__6808\,
            in1 => \N__6983\,
            in2 => \N__4920\,
            in3 => \N__6270\,
            lcout => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001101"
        )
    port map (
            in0 => \N__5375\,
            in1 => \N__6260\,
            in2 => \N__4917\,
            in3 => \N__6225\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9155\,
            ce => 'H',
            sr => \N__8928\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4892\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4838\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9155\,
            ce => 'H',
            sr => \N__8928\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6149\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9155\,
            ce => 'H',
            sr => \N__8928\
        );

    \U712_REG_SM.DS_EN_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__7559\,
            in1 => \N__4806\,
            in2 => \N__5079\,
            in3 => \N__6132\,
            lcout => \U712_REG_SM.DS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9155\,
            ce => 'H',
            sr => \N__8928\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000000000"
        )
    port map (
            in0 => \N__4788\,
            in1 => \N__6009\,
            in2 => \N__5997\,
            in3 => \N__4799\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9155\,
            ce => 'H',
            sr => \N__8928\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__7420\,
            in1 => \N__6391\,
            in2 => \_gnd_net_\,
            in3 => \N__6733\,
            lcout => \U712_REG_SM.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__5001\,
            in1 => \N__8577\,
            in2 => \_gnd_net_\,
            in3 => \N__8654\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9116\,
            ce => \N__8475\,
            sr => \N__8978\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__8539\,
            in1 => \N__8788\,
            in2 => \_gnd_net_\,
            in3 => \N__8614\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__5043\,
            in1 => \N__6279\,
            in2 => \N__5025\,
            in3 => \N__8153\,
            lcout => \U712_CHIP_RAM.N_369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__8538\,
            in1 => \N__5242\,
            in2 => \_gnd_net_\,
            in3 => \N__4995\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8161\,
            in1 => \N__4989\,
            in2 => \N__5739\,
            in3 => \N__4971\,
            lcout => \U712_CHIP_RAM.N_370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8536\,
            in1 => \N__8613\,
            in2 => \N__8769\,
            in3 => \N__7838\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => \U712_CHIP_RAM.REFRESH_RST_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__8537\,
            in1 => \N__8733\,
            in2 => \N__4938\,
            in3 => \N__7839\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVNIQ6_3_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5123\,
            in1 => \N__5791\,
            in2 => \N__5838\,
            in3 => \N__5139\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNICDSCD_0_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__5091\,
            in1 => \N__5277\,
            in2 => \N__5262\,
            in3 => \N__5259\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5229\,
            in2 => \N__5223\,
            in3 => \N__8768\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000100"
        )
    port map (
            in0 => \N__5220\,
            in1 => \N__5085\,
            in2 => \N__5187\,
            in3 => \N__5679\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_0_0_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__9021\,
            in1 => \_gnd_net_\,
            in2 => \N__5142\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__5590\,
            in1 => \N__5677\,
            in2 => \_gnd_net_\,
            in3 => \N__5514\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__5678\,
            in1 => \_gnd_net_\,
            in2 => \N__5131\,
            in3 => \N__7521\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__5912\,
            in1 => \N__5948\,
            in2 => \N__6051\,
            in3 => \N__5302\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_0_i_a3_0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI7TES1_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5578\,
            in1 => \N__5674\,
            in2 => \N__5518\,
            in3 => \N__6038\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIRB433_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__5911\,
            in1 => \N__5947\,
            in2 => \N__5841\,
            in3 => \N__5301\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5577\,
            in1 => \N__5673\,
            in2 => \_gnd_net_\,
            in3 => \N__5504\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5795\,
            in2 => \N__5805\,
            in3 => \N__5727\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110101"
        )
    port map (
            in0 => \N__6573\,
            in1 => \N__6660\,
            in2 => \N__8789\,
            in3 => \N__8104\,
            lcout => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5675\,
            in1 => \N__5582\,
            in2 => \_gnd_net_\,
            in3 => \N__5725\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__5726\,
            in1 => \N__5676\,
            in2 => \N__5599\,
            in3 => \N__5505\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111111011"
        )
    port map (
            in0 => \N__5460\,
            in1 => \N__5445\,
            in2 => \N__5436\,
            in3 => \N__5415\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9133\,
            ce => 'H',
            sr => \N__8938\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__8074\,
            in1 => \N__5406\,
            in2 => \_gnd_net_\,
            in3 => \N__6086\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9133\,
            ce => 'H',
            sr => \N__8938\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__5379\,
            in1 => \N__8075\,
            in2 => \N__5343\,
            in3 => \N__5306\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9133\,
            ce => 'H',
            sr => \N__8938\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__6168\,
            in1 => \N__6153\,
            in2 => \N__6054\,
            in3 => \N__6085\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9133\,
            ce => 'H',
            sr => \N__8938\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__5993\,
            in1 => \N__6861\,
            in2 => \_gnd_net_\,
            in3 => \N__6008\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9138\,
            ce => 'H',
            sr => \N__8933\
        );

    \U712_CHIP_RAM.DBR_SYNC_0_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5973\,
            lcout => \U712_REG_SM_DBR_SYNC_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9138\,
            ce => 'H',
            sr => \N__8933\
        );

    \U712_REG_SM.C1_SYNC_1_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6732\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9138\,
            ce => 'H',
            sr => \N__8933\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5946\,
            lcout => \U712_REG_SM_DBR_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9138\,
            ce => 'H',
            sr => \N__8933\
        );

    \U712_REG_SM.C1_SYNC_0_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5889\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9138\,
            ce => 'H',
            sr => \N__8933\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__6860\,
            in1 => \N__5853\,
            in2 => \N__6240\,
            in3 => \N__6259\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9148\,
            ce => 'H',
            sr => \N__8929\
        );

    \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__7142\,
            in1 => \N__5852\,
            in2 => \_gnd_net_\,
            in3 => \N__7100\,
            lcout => \U712_REG_SM.N_394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_1_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6398\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9148\,
            ce => 'H',
            sr => \N__8929\
        );

    \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7099\,
            in2 => \_gnd_net_\,
            in3 => \N__7141\,
            lcout => \U712_REG_SM.N_347\,
            ltout => \U712_REG_SM.N_347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6925\,
            in1 => \N__6768\,
            in2 => \N__6273\,
            in3 => \N__6720\,
            lcout => \U712_REG_SM.N_559\,
            ltout => \U712_REG_SM.N_559_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__6235\,
            in1 => \N__6258\,
            in2 => \N__6264\,
            in3 => \N__6809\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9148\,
            ce => 'H',
            sr => \N__8929\
        );

    \U712_REG_SM.REG_CYCLE_GO_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__6224\,
            in1 => \N__6261\,
            in2 => \N__6870\,
            in3 => \N__6236\,
            lcout => \U712_REG_SM.REG_CYCLE_GOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9148\,
            ce => 'H',
            sr => \N__8929\
        );

    \U712_REG_SM.REGENn_1_ess_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6779\,
            in1 => \N__6926\,
            in2 => \N__6743\,
            in3 => \N__6691\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9151\,
            ce => \N__6120\,
            sr => \N__8923\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__9016\,
            in1 => \N__6164\,
            in2 => \_gnd_net_\,
            in3 => \N__6148\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_1_ess_RNO_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9017\,
            in2 => \_gnd_net_\,
            in3 => \N__6131\,
            lcout => \U712_REG_SM.N_186_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6387\,
            in2 => \_gnd_net_\,
            in3 => \N__6428\,
            lcout => \U712_REG_SM.N_348\,
            ltout => \U712_REG_SM.N_348_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7001\,
            in2 => \N__6114\,
            in3 => \N__6692\,
            lcout => \U712_REG_SM.N_364\,
            ltout => \U712_REG_SM.N_364_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__6483\,
            in1 => \N__6952\,
            in2 => \N__6462\,
            in3 => \N__6459\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9156\,
            ce => 'H',
            sr => \N__8922\
        );

    \U712_REG_SM.C1_SYNC_2_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6780\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9156\,
            ce => 'H',
            sr => \N__8922\
        );

    \U712_REG_SM.C3_SYNC_0_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6417\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9156\,
            ce => 'H',
            sr => \N__8922\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8676\,
            in1 => \N__6366\,
            in2 => \_gnd_net_\,
            in3 => \N__8559\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9115\,
            ce => \N__8464\,
            sr => \N__8964\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000001"
        )
    port map (
            in0 => \N__8558\,
            in1 => \N__8677\,
            in2 => \N__8813\,
            in3 => \N__6285\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9115\,
            ce => \N__8464\,
            sr => \N__8964\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__8159\,
            in1 => \N__6648\,
            in2 => \N__6495\,
            in3 => \N__8758\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__6327\,
            in1 => \N__6306\,
            in2 => \N__6288\,
            in3 => \N__8160\,
            lcout => \U712_CHIP_RAM.N_368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__6540\,
            in1 => \N__8158\,
            in2 => \N__8790\,
            in3 => \N__6654\,
            lcout => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__6666\,
            in1 => \N__9020\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6567\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9119\,
            ce => \N__8193\,
            sr => \N__8942\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6527\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9119\,
            ce => \N__8193\,
            sr => \N__8942\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7983\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9119\,
            ce => \N__8193\,
            sr => \N__8942\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__9221\,
            in1 => \N__7281\,
            in2 => \N__6642\,
            in3 => \N__8154\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9122\,
            ce => \N__8467\,
            sr => \N__8935\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__6603\,
            in1 => \N__8576\,
            in2 => \_gnd_net_\,
            in3 => \N__8671\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9122\,
            ce => \N__8467\,
            sr => \N__8935\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8423\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9126\,
            ce => \N__7923\,
            sr => \N__8930\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6566\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9126\,
            ce => \N__7923\,
            sr => \N__8930\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6531\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9126\,
            ce => \N__7923\,
            sr => \N__8930\
        );

    \U712_REG_SM.C3_SYNC_2_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7148\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9131\,
            ce => 'H',
            sr => \N__8927\
        );

    \U712_BYTE_ENABLE.N_50_i_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100011"
        )
    port map (
            in0 => \N__6909\,
            in1 => \N__7083\,
            in2 => \N__7071\,
            in3 => \N__7047\,
            lcout => \N_50_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7002\,
            in1 => \N__6984\,
            in2 => \_gnd_net_\,
            in3 => \N__6810\,
            lcout => \U712_REG_SM.N_395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101010000"
        )
    port map (
            in0 => \N__6672\,
            in1 => \N__6972\,
            in2 => \N__6930\,
            in3 => \N__6951\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9141\,
            ce => 'H',
            sr => \N__8921\
        );

    \U712_REG_SM.LDS_OUT_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101111"
        )
    port map (
            in0 => \N__6907\,
            in1 => \N__6836\,
            in2 => \N__7340\,
            in3 => \N__6862\,
            lcout => \U712_REG_SM.LDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9141\,
            ce => 'H',
            sr => \N__8921\
        );

    \U712_REG_SM.UDS_OUT_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011111"
        )
    port map (
            in0 => \N__6908\,
            in1 => \N__7583\,
            in2 => \N__7341\,
            in3 => \N__6863\,
            lcout => \U712_REG_SM.UDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9141\,
            ce => 'H',
            sr => \N__8921\
        );

    \U712_REG_SM.LDS_OUT_RNIL31J_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7571\,
            lcout => \U712_REG_SM_un1_LDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6807\,
            in1 => \N__6778\,
            in2 => \N__6744\,
            in3 => \N__6693\,
            lcout => \U712_REG_SM.N_433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_RNIUP9B_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__7587\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7572\,
            lcout => \U712_REG_SM_un1_UDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7473\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDS_OUT_2_0_a3_0_a3_0_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__7425\,
            in1 => \N__7373\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.LDS_OUT_2_0_a3_0_a3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_13_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8578\,
            in1 => \N__8679\,
            in2 => \N__8820\,
            in3 => \N__7853\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9117\,
            ce => \N__8466\,
            sr => \N__8973\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8678\,
            in1 => \N__7653\,
            in2 => \_gnd_net_\,
            in3 => \N__8579\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9117\,
            ce => \N__8466\,
            sr => \N__8973\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_13_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__7280\,
            in1 => \N__7263\,
            in2 => \N__8358\,
            in3 => \N__8162\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9117\,
            ce => \N__8466\,
            sr => \N__8973\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__7224\,
            in1 => \N__7155\,
            in2 => \N__7203\,
            in3 => \N__8144\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_367_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8580\,
            in2 => \N__7176\,
            in3 => \N__8672\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9125\,
            ce => \N__8465\,
            sr => \N__8953\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7950\,
            in1 => \N__8142\,
            in2 => \N__8818\,
            in3 => \N__8202\,
            lcout => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8231\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9139\,
            ce => \N__7924\,
            sr => \N__8934\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8381\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9139\,
            ce => \N__7924\,
            sr => \N__8934\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001100100011"
        )
    port map (
            in0 => \N__7731\,
            in1 => \N__7611\,
            in2 => \N__8163\,
            in3 => \N__7716\,
            lcout => \U712_CHIP_RAM.N_372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__7695\,
            in1 => \N__8152\,
            in2 => \N__7677\,
            in3 => \N__7599\,
            lcout => \U712_CHIP_RAM.N_371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__7647\,
            in1 => \N__8151\,
            in2 => \N__7629\,
            in3 => \N__7989\,
            lcout => \U712_CHIP_RAM.N_373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__8130\,
            in1 => \N__7605\,
            in2 => \N__8800\,
            in3 => \N__8310\,
            lcout => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8304\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9129\,
            ce => \N__7935\,
            sr => \N__8967\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010011"
        )
    port map (
            in0 => \N__8391\,
            in1 => \N__7593\,
            in2 => \N__8802\,
            in3 => \N__8143\,
            lcout => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8339\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9129\,
            ce => \N__7935\,
            sr => \N__8967\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__8131\,
            in1 => \N__7944\,
            in2 => \N__8801\,
            in3 => \N__8280\,
            lcout => \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7976\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9134\,
            ce => \N__7931\,
            sr => \N__8954\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8274\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9134\,
            ce => \N__7931\,
            sr => \N__8954\
        );

    \U712_CHIP_RAM.CASn_LC_15_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8812\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9118\,
            ce => 'H',
            sr => \N__8982\
        );

    \U712_CHIP_RAM.WEn_LC_15_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8673\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9118\,
            ce => 'H',
            sr => \N__8982\
        );

    \U712_CHIP_RAM.CRCSn_LC_15_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7857\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9121\,
            ce => 'H',
            sr => \N__8981\
        );

    \U712_CHIP_RAM.RASn_LC_15_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8583\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9121\,
            ce => 'H',
            sr => \N__8981\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__7779\,
            in1 => \_gnd_net_\,
            in2 => \N__8675\,
            in3 => \N__8581\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9130\,
            ce => \N__8474\,
            sr => \N__8979\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100011"
        )
    port map (
            in0 => \N__8826\,
            in1 => \N__8819\,
            in2 => \N__8674\,
            in3 => \N__8582\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9130\,
            ce => \N__8474\,
            sr => \N__8979\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8424\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9135\,
            ce => \N__8186\,
            sr => \N__8974\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8385\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9135\,
            ce => \N__8186\,
            sr => \N__8974\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8343\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9135\,
            ce => \N__8186\,
            sr => \N__8974\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8303\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9135\,
            ce => \N__8186\,
            sr => \N__8974\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8270\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9140\,
            ce => \N__8185\,
            sr => \N__8968\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8232\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9140\,
            ce => \N__8185\,
            sr => \N__8968\
        );

    \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__9027\,
            in1 => \N__8169\,
            in2 => \_gnd_net_\,
            in3 => \N__9173\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9174\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9152\,
            ce => 'H',
            sr => \N__8980\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9222\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9189\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9152\,
            ce => 'H',
            sr => \N__8980\
        );
end \INTERFACE\;

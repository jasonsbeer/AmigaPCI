-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 8 2025 20:42:07

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    TSn : in std_logic;
    RASn : out std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__10182\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \N_981_i\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_2\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.un5_DMA_CYCLE_START_0\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_1_cascade_\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_1_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_i_i_a3_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_e_1_cascade_\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.N_176_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_166_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_313\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_9_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.N_232_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0_a3_1\ : std_logic;
signal \U712_CHIP_RAM.N_232\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_167_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_9_0_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNIIGLS1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_176\ : std_logic;
signal \U712_CHIP_RAM.N_230_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_a3_1_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_285_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\ : std_logic;
signal \U712_CHIP_RAM.N_314\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.N_167\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_53\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_196_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_315\ : std_logic;
signal \U712_CHIP_RAM.N_197_i_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_233\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8RZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_219_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_166\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_7_i_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_258\ : std_logic;
signal \U712_CHIP_RAM.N_49_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_206\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_BYTE_ENABLE.N_268\ : std_logic;
signal \N_185_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_270_cascade_\ : std_logic;
signal \N_186_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_272\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0\ : std_logic;
signal \N_187_i\ : std_logic;
signal \A_c_1\ : std_logic;
signal \U712_BYTE_ENABLE.N_265\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_266_cascade_\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \N_184_i\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \DRDDIR_i_m2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \A_c_14\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_324_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \RnW_c\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_248\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2Z0Z_1\ : std_logic;
signal \U712_REG_SM.N_171_cascade_\ : std_logic;
signal \U712_REG_SM.DS_EN_0_sqmuxa_0_a2_0_a3_1_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \U712_REG_SM.N_199_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.N_208_i_0_en_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_208_i_0_en_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a3_0_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_165\ : std_logic;
signal \U712_CHIP_RAM.N_249\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_REG_SM.N_199\ : std_logic;
signal \U712_REG_SM.N_171\ : std_logic;
signal \U712_REG_SM.N_174_cascade_\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_210\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_5\ : std_logic;
signal \U712_REG_SM.N_174\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \CASn_c\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_2\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_RNITQLC2Z0Z_1\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_GOZ0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.DS_EN_0_sqmuxa\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_205\ : std_logic;
signal \U712_REG_SM.N_202\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \N_118\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \DS_ENm\ : std_logic;
signal \N_113\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CLK40_OUT_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    CLK_EN <= \CLK_EN_wire\;
    \RESETn_wire\ <= RESETn;
    LDSn <= \LDSn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CLK40_OUT <= \CLK40_OUT_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__3620\,
            RESETB => \N__4373\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10182\,
            DIN => \N__10181\,
            DOUT => \N__10180\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10182\,
            PADOUT => \N__10181\,
            PADIN => \N__10180\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5645\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10173\,
            DIN => \N__10172\,
            DOUT => \N__10171\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10173\,
            PADOUT => \N__10172\,
            PADIN => \N__10171\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10164\,
            DIN => \N__10163\,
            DOUT => \N__10162\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10164\,
            PADOUT => \N__10163\,
            PADIN => \N__10162\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6950\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10155\,
            DIN => \N__10154\,
            DOUT => \N__10153\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10155\,
            PADOUT => \N__10154\,
            PADIN => \N__10153\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5297\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10146\,
            DIN => \N__10145\,
            DOUT => \N__10144\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10146\,
            PADOUT => \N__10145\,
            PADIN => \N__10144\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10137\,
            DIN => \N__10136\,
            DOUT => \N__10135\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10137\,
            PADOUT => \N__10136\,
            PADIN => \N__10135\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10128\,
            DIN => \N__10127\,
            DOUT => \N__10126\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10128\,
            PADOUT => \N__10127\,
            PADIN => \N__10126\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10119\,
            DIN => \N__10118\,
            DOUT => \N__10117\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10119\,
            PADOUT => \N__10118\,
            PADIN => \N__10117\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10110\,
            DIN => \N__10109\,
            DOUT => \N__10108\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10110\,
            PADOUT => \N__10109\,
            PADIN => \N__10108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10101\,
            DIN => \N__10100\,
            DOUT => \N__10099\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10101\,
            PADOUT => \N__10100\,
            PADIN => \N__10099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5741\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10092\,
            DIN => \N__10091\,
            DOUT => \N__10090\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10092\,
            PADOUT => \N__10091\,
            PADIN => \N__10090\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10083\,
            DIN => \N__10082\,
            DOUT => \N__10081\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10083\,
            PADOUT => \N__10082\,
            PADIN => \N__10081\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10074\,
            DIN => \N__10073\,
            DOUT => \N__10072\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10074\,
            PADOUT => \N__10073\,
            PADIN => \N__10072\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10065\,
            DIN => \N__10064\,
            DOUT => \N__10063\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10065\,
            PADOUT => \N__10064\,
            PADIN => \N__10063\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3893\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10056\,
            DIN => \N__10055\,
            DOUT => \N__10054\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10056\,
            PADOUT => \N__10055\,
            PADIN => \N__10054\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10047\,
            DIN => \N__10046\,
            DOUT => \N__10045\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10047\,
            PADOUT => \N__10046\,
            PADIN => \N__10045\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10038\,
            DIN => \N__10037\,
            DOUT => \N__10036\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10038\,
            PADOUT => \N__10037\,
            PADIN => \N__10036\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5270\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10029\,
            DIN => \N__10028\,
            DOUT => \N__10027\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10029\,
            PADOUT => \N__10028\,
            PADIN => \N__10027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10020\,
            DIN => \N__10019\,
            DOUT => \N__10018\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10020\,
            PADOUT => \N__10019\,
            PADIN => \N__10018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8162\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10011\,
            DIN => \N__10010\,
            DOUT => \N__10009\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10011\,
            PADOUT => \N__10010\,
            PADIN => \N__10009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10002\,
            DIN => \N__10001\,
            DOUT => \N__10000\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10002\,
            PADOUT => \N__10001\,
            PADIN => \N__10000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9993\,
            DIN => \N__9992\,
            DOUT => \N__9991\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9993\,
            PADOUT => \N__9992\,
            PADIN => \N__9991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9984\,
            DIN => \N__9983\,
            DOUT => \N__9982\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9984\,
            PADOUT => \N__9983\,
            PADIN => \N__9982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9975\,
            DIN => \N__9974\,
            DOUT => \N__9973\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9975\,
            PADOUT => \N__9974\,
            PADIN => \N__9973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9966\,
            DIN => \N__9965\,
            DOUT => \N__9964\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9966\,
            PADOUT => \N__9965\,
            PADIN => \N__9964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4238\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9957\,
            DIN => \N__9956\,
            DOUT => \N__9955\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9957\,
            PADOUT => \N__9956\,
            PADIN => \N__9955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9948\,
            DIN => \N__9947\,
            DOUT => \N__9946\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9948\,
            PADOUT => \N__9947\,
            PADIN => \N__9946\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9939\,
            DIN => \N__9938\,
            DOUT => \N__9937\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9939\,
            PADOUT => \N__9938\,
            PADIN => \N__9937\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9930\,
            DIN => \N__9929\,
            DOUT => \N__9928\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9930\,
            PADOUT => \N__9929\,
            PADIN => \N__9928\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9921\,
            DIN => \N__9920\,
            DOUT => \N__9919\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9921\,
            PADOUT => \N__9920\,
            PADIN => \N__9919\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9912\,
            DIN => \N__9911\,
            DOUT => \N__9910\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9912\,
            PADOUT => \N__9911\,
            PADIN => \N__9910\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5714\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9903\,
            DIN => \N__9902\,
            DOUT => \N__9901\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9903\,
            PADOUT => \N__9902\,
            PADIN => \N__9901\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9894\,
            DIN => \N__9893\,
            DOUT => \N__9892\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9894\,
            PADOUT => \N__9893\,
            PADIN => \N__9892\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9885\,
            DIN => \N__9884\,
            DOUT => \N__9883\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9885\,
            PADOUT => \N__9884\,
            PADIN => \N__9883\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9876\,
            DIN => \N__9875\,
            DOUT => \N__9874\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9876\,
            PADOUT => \N__9875\,
            PADIN => \N__9874\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9867\,
            DIN => \N__9866\,
            DOUT => \N__9865\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9867\,
            PADOUT => \N__9866\,
            PADIN => \N__9865\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8342\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9858\,
            DIN => \N__9857\,
            DOUT => \N__9856\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9858\,
            PADOUT => \N__9857\,
            PADIN => \N__9856\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9849\,
            DIN => \N__9848\,
            DOUT => \N__9847\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9849\,
            PADOUT => \N__9848\,
            PADIN => \N__9847\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8030\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9840\,
            DIN => \N__9839\,
            DOUT => \N__9838\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9840\,
            PADOUT => \N__9839\,
            PADIN => \N__9838\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9831\,
            DIN => \N__9830\,
            DOUT => \N__9829\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9831\,
            PADOUT => \N__9830\,
            PADIN => \N__9829\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9822\,
            DIN => \N__9821\,
            DOUT => \N__9820\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9822\,
            PADOUT => \N__9821\,
            PADIN => \N__9820\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3728\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9813\,
            DIN => \N__9812\,
            DOUT => \N__9811\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9813\,
            PADOUT => \N__9812\,
            PADIN => \N__9811\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7709\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9804\,
            DIN => \N__9803\,
            DOUT => \N__9802\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9804\,
            PADOUT => \N__9803\,
            PADIN => \N__9802\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6815\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9795\,
            DIN => \N__9794\,
            DOUT => \N__9793\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9795\,
            PADOUT => \N__9794\,
            PADIN => \N__9793\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9786\,
            DIN => \N__9785\,
            DOUT => \N__9784\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9786\,
            PADOUT => \N__9785\,
            PADIN => \N__9784\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9777\,
            DIN => \N__9776\,
            DOUT => \N__9775\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9777\,
            PADOUT => \N__9776\,
            PADIN => \N__9775\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9768\,
            DIN => \N__9767\,
            DOUT => \N__9766\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9768\,
            PADOUT => \N__9767\,
            PADIN => \N__9766\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6935\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9759\,
            DIN => \N__9758\,
            DOUT => \N__9757\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9759\,
            PADOUT => \N__9758\,
            PADIN => \N__9757\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9750\,
            DIN => \N__9749\,
            DOUT => \N__9748\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9750\,
            PADOUT => \N__9749\,
            PADIN => \N__9748\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5681\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9741\,
            DIN => \N__9740\,
            DOUT => \N__9739\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9741\,
            PADOUT => \N__9740\,
            PADIN => \N__9739\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4022\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9732\,
            DIN => \N__9731\,
            DOUT => \N__9730\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9732\,
            PADOUT => \N__9731\,
            PADIN => \N__9730\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5480\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9723\,
            DIN => \N__9722\,
            DOUT => \N__9721\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9723\,
            PADOUT => \N__9722\,
            PADIN => \N__9721\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7988\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9714\,
            DIN => \N__9713\,
            DOUT => \N__9712\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9714\,
            PADOUT => \N__9713\,
            PADIN => \N__9712\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7708\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9705\,
            DIN => \N__9704\,
            DOUT => \N__9703\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9705\,
            PADOUT => \N__9704\,
            PADIN => \N__9703\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9696\,
            DIN => \N__9695\,
            DOUT => \N__9694\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9696\,
            PADOUT => \N__9695\,
            PADIN => \N__9694\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9687\,
            DIN => \N__9686\,
            DOUT => \N__9685\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9687\,
            PADOUT => \N__9686\,
            PADIN => \N__9685\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5570\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9678\,
            DIN => \N__9677\,
            DOUT => \N__9676\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9678\,
            PADOUT => \N__9677\,
            PADIN => \N__9676\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8093\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9669\,
            DIN => \N__9668\,
            DOUT => \N__9667\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9669\,
            PADOUT => \N__9668\,
            PADIN => \N__9667\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3923\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9660\,
            DIN => \N__9659\,
            DOUT => \N__9658\,
            PACKAGEPIN => \CLK40_OUT_wire\
        );

    \CLK40_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9660\,
            PADOUT => \N__9659\,
            PADIN => \N__9658\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3647\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9651\,
            DIN => \N__9650\,
            DOUT => \N__9649\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9651\,
            PADOUT => \N__9650\,
            PADIN => \N__9649\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5597\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9642\,
            DIN => \N__9641\,
            DOUT => \N__9640\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9642\,
            PADOUT => \N__9641\,
            PADIN => \N__9640\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9633\,
            DIN => \N__9632\,
            DOUT => \N__9631\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9633\,
            PADOUT => \N__9632\,
            PADIN => \N__9631\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9624\,
            DIN => \N__9623\,
            DOUT => \N__9622\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9624\,
            PADOUT => \N__9623\,
            PADIN => \N__9622\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9615\,
            DIN => \N__9614\,
            DOUT => \N__9613\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9615\,
            PADOUT => \N__9614\,
            PADIN => \N__9613\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9606\,
            DIN => \N__9605\,
            DOUT => \N__9604\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9606\,
            PADOUT => \N__9605\,
            PADIN => \N__9604\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5831\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9597\,
            DIN => \N__9596\,
            DOUT => \N__9595\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9597\,
            PADOUT => \N__9596\,
            PADIN => \N__9595\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9588\,
            DIN => \N__9587\,
            DOUT => \N__9586\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9588\,
            PADOUT => \N__9587\,
            PADIN => \N__9586\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5366\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9579\,
            DIN => \N__9578\,
            DOUT => \N__9577\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9579\,
            PADOUT => \N__9578\,
            PADIN => \N__9577\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3638\,
            DIN0 => OPEN,
            DOUT0 => \N__3689\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9570\,
            DIN => \N__9569\,
            DOUT => \N__9568\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9570\,
            PADOUT => \N__9569\,
            PADIN => \N__9568\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6902\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9561\,
            DIN => \N__9560\,
            DOUT => \N__9559\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9561\,
            PADOUT => \N__9560\,
            PADIN => \N__9559\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9552\,
            DIN => \N__9551\,
            DOUT => \N__9550\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9552\,
            PADOUT => \N__9551\,
            PADIN => \N__9550\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9543\,
            DIN => \N__9542\,
            DOUT => \N__9541\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9543\,
            PADOUT => \N__9542\,
            PADIN => \N__9541\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7763\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9534\,
            DIN => \N__9533\,
            DOUT => \N__9532\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9534\,
            PADOUT => \N__9533\,
            PADIN => \N__9532\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9525\,
            DIN => \N__9524\,
            DOUT => \N__9523\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9525\,
            PADOUT => \N__9524\,
            PADIN => \N__9523\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9516\,
            DIN => \N__9515\,
            DOUT => \N__9514\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9516\,
            PADOUT => \N__9515\,
            PADIN => \N__9514\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9507\,
            DIN => \N__9506\,
            DOUT => \N__9505\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9507\,
            PADOUT => \N__9506\,
            PADIN => \N__9505\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9498\,
            DIN => \N__9497\,
            DOUT => \N__9496\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9498\,
            PADOUT => \N__9497\,
            PADIN => \N__9496\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5798\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9489\,
            DIN => \N__9488\,
            DOUT => \N__9487\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9489\,
            PADOUT => \N__9488\,
            PADIN => \N__9487\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8216\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2267\ : InMux
    port map (
            O => \N__9470\,
            I => \N__9466\
        );

    \I__2266\ : InMux
    port map (
            O => \N__9469\,
            I => \N__9463\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__9466\,
            I => \N__9458\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__9463\,
            I => \N__9458\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__2262\ : Span4Mux_v
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__2261\ : Sp12to4
    port map (
            O => \N__9452\,
            I => \N__9449\
        );

    \I__2260\ : Span12Mux_h
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__2259\ : Odrv12
    port map (
            O => \N__9446\,
            I => \DRA_c_3\
        );

    \I__2258\ : InMux
    port map (
            O => \N__9443\,
            I => \N__9440\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__9440\,
            I => \N__9437\
        );

    \I__2256\ : Span4Mux_h
    port map (
            O => \N__9437\,
            I => \N__9434\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__9434\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2254\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__9428\,
            I => \N__9424\
        );

    \I__2252\ : InMux
    port map (
            O => \N__9427\,
            I => \N__9421\
        );

    \I__2251\ : Span12Mux_v
    port map (
            O => \N__9424\,
            I => \N__9416\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__9421\,
            I => \N__9416\
        );

    \I__2249\ : Span12Mux_h
    port map (
            O => \N__9416\,
            I => \N__9413\
        );

    \I__2248\ : Odrv12
    port map (
            O => \N__9413\,
            I => \DRA_c_8\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__9410\,
            I => \N__9407\
        );

    \I__2246\ : InMux
    port map (
            O => \N__9407\,
            I => \N__9404\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__9404\,
            I => \N__9401\
        );

    \I__2244\ : Span4Mux_h
    port map (
            O => \N__9401\,
            I => \N__9398\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__9398\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9395\,
            I => \N__9392\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__9392\,
            I => \N__9382\
        );

    \I__2240\ : ClkMux
    port map (
            O => \N__9391\,
            I => \N__9365\
        );

    \I__2239\ : ClkMux
    port map (
            O => \N__9390\,
            I => \N__9365\
        );

    \I__2238\ : ClkMux
    port map (
            O => \N__9389\,
            I => \N__9365\
        );

    \I__2237\ : ClkMux
    port map (
            O => \N__9388\,
            I => \N__9365\
        );

    \I__2236\ : ClkMux
    port map (
            O => \N__9387\,
            I => \N__9365\
        );

    \I__2235\ : ClkMux
    port map (
            O => \N__9386\,
            I => \N__9365\
        );

    \I__2234\ : ClkMux
    port map (
            O => \N__9385\,
            I => \N__9365\
        );

    \I__2233\ : Glb2LocalMux
    port map (
            O => \N__9382\,
            I => \N__9365\
        );

    \I__2232\ : GlobalMux
    port map (
            O => \N__9365\,
            I => \N__9362\
        );

    \I__2231\ : gio2CtrlBuf
    port map (
            O => \N__9362\,
            I => \C3_c_g\
        );

    \I__2230\ : CEMux
    port map (
            O => \N__9359\,
            I => \N__9356\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__9356\,
            I => \N__9348\
        );

    \I__2228\ : CEMux
    port map (
            O => \N__9355\,
            I => \N__9345\
        );

    \I__2227\ : CEMux
    port map (
            O => \N__9354\,
            I => \N__9342\
        );

    \I__2226\ : CEMux
    port map (
            O => \N__9353\,
            I => \N__9338\
        );

    \I__2225\ : CEMux
    port map (
            O => \N__9352\,
            I => \N__9335\
        );

    \I__2224\ : CEMux
    port map (
            O => \N__9351\,
            I => \N__9332\
        );

    \I__2223\ : Span4Mux_v
    port map (
            O => \N__9348\,
            I => \N__9329\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__9345\,
            I => \N__9324\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__9342\,
            I => \N__9324\
        );

    \I__2220\ : CEMux
    port map (
            O => \N__9341\,
            I => \N__9321\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__9338\,
            I => \N__9318\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__9335\,
            I => \N__9315\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__9332\,
            I => \N__9312\
        );

    \I__2216\ : Span4Mux_h
    port map (
            O => \N__9329\,
            I => \N__9305\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__9324\,
            I => \N__9305\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__9321\,
            I => \N__9305\
        );

    \I__2213\ : Span4Mux_v
    port map (
            O => \N__9318\,
            I => \N__9302\
        );

    \I__2212\ : Span4Mux_h
    port map (
            O => \N__9315\,
            I => \N__9299\
        );

    \I__2211\ : Span4Mux_v
    port map (
            O => \N__9312\,
            I => \N__9294\
        );

    \I__2210\ : Span4Mux_h
    port map (
            O => \N__9305\,
            I => \N__9294\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__9302\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\
        );

    \I__2208\ : Odrv4
    port map (
            O => \N__9299\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\
        );

    \I__2207\ : Odrv4
    port map (
            O => \N__9294\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\
        );

    \I__2206\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9280\
        );

    \I__2205\ : InMux
    port map (
            O => \N__9286\,
            I => \N__9277\
        );

    \I__2204\ : InMux
    port map (
            O => \N__9285\,
            I => \N__9274\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9271\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9268\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__9280\,
            I => \N__9250\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__9277\,
            I => \N__9240\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__9274\,
            I => \N__9224\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__9271\,
            I => \N__9218\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__9268\,
            I => \N__9213\
        );

    \I__2196\ : SRMux
    port map (
            O => \N__9267\,
            I => \N__9122\
        );

    \I__2195\ : SRMux
    port map (
            O => \N__9266\,
            I => \N__9122\
        );

    \I__2194\ : SRMux
    port map (
            O => \N__9265\,
            I => \N__9122\
        );

    \I__2193\ : SRMux
    port map (
            O => \N__9264\,
            I => \N__9122\
        );

    \I__2192\ : SRMux
    port map (
            O => \N__9263\,
            I => \N__9122\
        );

    \I__2191\ : SRMux
    port map (
            O => \N__9262\,
            I => \N__9122\
        );

    \I__2190\ : SRMux
    port map (
            O => \N__9261\,
            I => \N__9122\
        );

    \I__2189\ : SRMux
    port map (
            O => \N__9260\,
            I => \N__9122\
        );

    \I__2188\ : SRMux
    port map (
            O => \N__9259\,
            I => \N__9122\
        );

    \I__2187\ : SRMux
    port map (
            O => \N__9258\,
            I => \N__9122\
        );

    \I__2186\ : SRMux
    port map (
            O => \N__9257\,
            I => \N__9122\
        );

    \I__2185\ : SRMux
    port map (
            O => \N__9256\,
            I => \N__9122\
        );

    \I__2184\ : SRMux
    port map (
            O => \N__9255\,
            I => \N__9122\
        );

    \I__2183\ : SRMux
    port map (
            O => \N__9254\,
            I => \N__9122\
        );

    \I__2182\ : SRMux
    port map (
            O => \N__9253\,
            I => \N__9122\
        );

    \I__2181\ : Glb2LocalMux
    port map (
            O => \N__9250\,
            I => \N__9122\
        );

    \I__2180\ : SRMux
    port map (
            O => \N__9249\,
            I => \N__9122\
        );

    \I__2179\ : SRMux
    port map (
            O => \N__9248\,
            I => \N__9122\
        );

    \I__2178\ : SRMux
    port map (
            O => \N__9247\,
            I => \N__9122\
        );

    \I__2177\ : SRMux
    port map (
            O => \N__9246\,
            I => \N__9122\
        );

    \I__2176\ : SRMux
    port map (
            O => \N__9245\,
            I => \N__9122\
        );

    \I__2175\ : SRMux
    port map (
            O => \N__9244\,
            I => \N__9122\
        );

    \I__2174\ : SRMux
    port map (
            O => \N__9243\,
            I => \N__9122\
        );

    \I__2173\ : Glb2LocalMux
    port map (
            O => \N__9240\,
            I => \N__9122\
        );

    \I__2172\ : SRMux
    port map (
            O => \N__9239\,
            I => \N__9122\
        );

    \I__2171\ : SRMux
    port map (
            O => \N__9238\,
            I => \N__9122\
        );

    \I__2170\ : SRMux
    port map (
            O => \N__9237\,
            I => \N__9122\
        );

    \I__2169\ : SRMux
    port map (
            O => \N__9236\,
            I => \N__9122\
        );

    \I__2168\ : SRMux
    port map (
            O => \N__9235\,
            I => \N__9122\
        );

    \I__2167\ : SRMux
    port map (
            O => \N__9234\,
            I => \N__9122\
        );

    \I__2166\ : SRMux
    port map (
            O => \N__9233\,
            I => \N__9122\
        );

    \I__2165\ : SRMux
    port map (
            O => \N__9232\,
            I => \N__9122\
        );

    \I__2164\ : SRMux
    port map (
            O => \N__9231\,
            I => \N__9122\
        );

    \I__2163\ : SRMux
    port map (
            O => \N__9230\,
            I => \N__9122\
        );

    \I__2162\ : SRMux
    port map (
            O => \N__9229\,
            I => \N__9122\
        );

    \I__2161\ : SRMux
    port map (
            O => \N__9228\,
            I => \N__9122\
        );

    \I__2160\ : SRMux
    port map (
            O => \N__9227\,
            I => \N__9122\
        );

    \I__2159\ : Glb2LocalMux
    port map (
            O => \N__9224\,
            I => \N__9122\
        );

    \I__2158\ : SRMux
    port map (
            O => \N__9223\,
            I => \N__9122\
        );

    \I__2157\ : SRMux
    port map (
            O => \N__9222\,
            I => \N__9122\
        );

    \I__2156\ : SRMux
    port map (
            O => \N__9221\,
            I => \N__9122\
        );

    \I__2155\ : Glb2LocalMux
    port map (
            O => \N__9218\,
            I => \N__9122\
        );

    \I__2154\ : SRMux
    port map (
            O => \N__9217\,
            I => \N__9122\
        );

    \I__2153\ : SRMux
    port map (
            O => \N__9216\,
            I => \N__9122\
        );

    \I__2152\ : Glb2LocalMux
    port map (
            O => \N__9213\,
            I => \N__9122\
        );

    \I__2151\ : GlobalMux
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__2150\ : gio2CtrlBuf
    port map (
            O => \N__9119\,
            I => \RESETn_c_i_g\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9116\,
            I => \N__9113\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9113\,
            I => \N__9109\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9112\,
            I => \N__9106\
        );

    \I__2146\ : Sp12to4
    port map (
            O => \N__9109\,
            I => \N__9101\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__9106\,
            I => \N__9101\
        );

    \I__2144\ : Span12Mux_v
    port map (
            O => \N__9101\,
            I => \N__9098\
        );

    \I__2143\ : Span12Mux_h
    port map (
            O => \N__9098\,
            I => \N__9095\
        );

    \I__2142\ : Odrv12
    port map (
            O => \N__9095\,
            I => \DRA_c_6\
        );

    \I__2141\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9089\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__9089\,
            I => \N__9086\
        );

    \I__2139\ : Span4Mux_v
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__9083\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9077\,
            I => \N__9073\
        );

    \I__2135\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9070\
        );

    \I__2134\ : Span4Mux_h
    port map (
            O => \N__9073\,
            I => \N__9065\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__9070\,
            I => \N__9065\
        );

    \I__2132\ : Span4Mux_v
    port map (
            O => \N__9065\,
            I => \N__9062\
        );

    \I__2131\ : Sp12to4
    port map (
            O => \N__9062\,
            I => \N__9059\
        );

    \I__2130\ : Span12Mux_h
    port map (
            O => \N__9059\,
            I => \N__9056\
        );

    \I__2129\ : Span12Mux_v
    port map (
            O => \N__9056\,
            I => \N__9053\
        );

    \I__2128\ : Odrv12
    port map (
            O => \N__9053\,
            I => \DRA_c_4\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9050\,
            I => \N__9047\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__9047\,
            I => \N__9044\
        );

    \I__2125\ : Span4Mux_h
    port map (
            O => \N__9044\,
            I => \N__9041\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__9041\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__2121\ : Span4Mux_h
    port map (
            O => \N__9032\,
            I => \N__9029\
        );

    \I__2120\ : Odrv4
    port map (
            O => \N__9029\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9026\,
            I => \N__9023\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9023\,
            I => \N__9020\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__9020\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__9017\,
            I => \N__9014\
        );

    \I__2115\ : InMux
    port map (
            O => \N__9014\,
            I => \N__9011\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__9011\,
            I => \N__9008\
        );

    \I__2113\ : Span4Mux_h
    port map (
            O => \N__9008\,
            I => \N__9005\
        );

    \I__2112\ : Odrv4
    port map (
            O => \N__9005\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2111\ : InMux
    port map (
            O => \N__9002\,
            I => \N__8999\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__8999\,
            I => \N__8995\
        );

    \I__2109\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8992\
        );

    \I__2108\ : Sp12to4
    port map (
            O => \N__8995\,
            I => \N__8987\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__8992\,
            I => \N__8987\
        );

    \I__2106\ : Span12Mux_v
    port map (
            O => \N__8987\,
            I => \N__8984\
        );

    \I__2105\ : Span12Mux_h
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__2104\ : Odrv12
    port map (
            O => \N__8981\,
            I => \DRA_c_2\
        );

    \I__2103\ : InMux
    port map (
            O => \N__8978\,
            I => \N__8972\
        );

    \I__2102\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8972\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__8972\,
            I => \N__8969\
        );

    \I__2100\ : Span4Mux_h
    port map (
            O => \N__8969\,
            I => \N__8966\
        );

    \I__2099\ : Odrv4
    port map (
            O => \N__8966\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2098\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8959\
        );

    \I__2097\ : InMux
    port map (
            O => \N__8962\,
            I => \N__8956\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__8959\,
            I => \N__8951\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__8956\,
            I => \N__8951\
        );

    \I__2094\ : Span12Mux_v
    port map (
            O => \N__8951\,
            I => \N__8948\
        );

    \I__2093\ : Span12Mux_h
    port map (
            O => \N__8948\,
            I => \N__8945\
        );

    \I__2092\ : Span12Mux_v
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__2091\ : Odrv12
    port map (
            O => \N__8942\,
            I => \DRA_c_9\
        );

    \I__2090\ : InMux
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__8936\,
            I => \N__8933\
        );

    \I__2088\ : Span12Mux_v
    port map (
            O => \N__8933\,
            I => \N__8930\
        );

    \I__2087\ : Odrv12
    port map (
            O => \N__8930\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2086\ : CEMux
    port map (
            O => \N__8927\,
            I => \N__8924\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__8924\,
            I => \N__8917\
        );

    \I__2084\ : CEMux
    port map (
            O => \N__8923\,
            I => \N__8914\
        );

    \I__2083\ : CEMux
    port map (
            O => \N__8922\,
            I => \N__8911\
        );

    \I__2082\ : CEMux
    port map (
            O => \N__8921\,
            I => \N__8908\
        );

    \I__2081\ : CEMux
    port map (
            O => \N__8920\,
            I => \N__8905\
        );

    \I__2080\ : Span4Mux_h
    port map (
            O => \N__8917\,
            I => \N__8899\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__8914\,
            I => \N__8899\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__8911\,
            I => \N__8896\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__8908\,
            I => \N__8893\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__8905\,
            I => \N__8890\
        );

    \I__2075\ : CEMux
    port map (
            O => \N__8904\,
            I => \N__8887\
        );

    \I__2074\ : Span4Mux_v
    port map (
            O => \N__8899\,
            I => \N__8884\
        );

    \I__2073\ : Span4Mux_v
    port map (
            O => \N__8896\,
            I => \N__8875\
        );

    \I__2072\ : Span4Mux_h
    port map (
            O => \N__8893\,
            I => \N__8875\
        );

    \I__2071\ : Span4Mux_v
    port map (
            O => \N__8890\,
            I => \N__8875\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__8887\,
            I => \N__8875\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__8884\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__8875\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\
        );

    \I__2067\ : InMux
    port map (
            O => \N__8870\,
            I => \N__8867\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__8867\,
            I => \N__8864\
        );

    \I__2065\ : Span4Mux_v
    port map (
            O => \N__8864\,
            I => \N__8861\
        );

    \I__2064\ : Sp12to4
    port map (
            O => \N__8861\,
            I => \N__8858\
        );

    \I__2063\ : Span12Mux_h
    port map (
            O => \N__8858\,
            I => \N__8855\
        );

    \I__2062\ : Odrv12
    port map (
            O => \N__8855\,
            I => \RAS0n_c\
        );

    \I__2061\ : InMux
    port map (
            O => \N__8852\,
            I => \N__8849\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__8849\,
            I => \N__8846\
        );

    \I__2059\ : Span4Mux_v
    port map (
            O => \N__8846\,
            I => \N__8843\
        );

    \I__2058\ : Odrv4
    port map (
            O => \N__8843\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2057\ : InMux
    port map (
            O => \N__8840\,
            I => \N__8837\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__8837\,
            I => \N__8810\
        );

    \I__2055\ : ClkMux
    port map (
            O => \N__8836\,
            I => \N__8732\
        );

    \I__2054\ : ClkMux
    port map (
            O => \N__8835\,
            I => \N__8732\
        );

    \I__2053\ : ClkMux
    port map (
            O => \N__8834\,
            I => \N__8732\
        );

    \I__2052\ : ClkMux
    port map (
            O => \N__8833\,
            I => \N__8732\
        );

    \I__2051\ : ClkMux
    port map (
            O => \N__8832\,
            I => \N__8732\
        );

    \I__2050\ : ClkMux
    port map (
            O => \N__8831\,
            I => \N__8732\
        );

    \I__2049\ : ClkMux
    port map (
            O => \N__8830\,
            I => \N__8732\
        );

    \I__2048\ : ClkMux
    port map (
            O => \N__8829\,
            I => \N__8732\
        );

    \I__2047\ : ClkMux
    port map (
            O => \N__8828\,
            I => \N__8732\
        );

    \I__2046\ : ClkMux
    port map (
            O => \N__8827\,
            I => \N__8732\
        );

    \I__2045\ : ClkMux
    port map (
            O => \N__8826\,
            I => \N__8732\
        );

    \I__2044\ : ClkMux
    port map (
            O => \N__8825\,
            I => \N__8732\
        );

    \I__2043\ : ClkMux
    port map (
            O => \N__8824\,
            I => \N__8732\
        );

    \I__2042\ : ClkMux
    port map (
            O => \N__8823\,
            I => \N__8732\
        );

    \I__2041\ : ClkMux
    port map (
            O => \N__8822\,
            I => \N__8732\
        );

    \I__2040\ : ClkMux
    port map (
            O => \N__8821\,
            I => \N__8732\
        );

    \I__2039\ : ClkMux
    port map (
            O => \N__8820\,
            I => \N__8732\
        );

    \I__2038\ : ClkMux
    port map (
            O => \N__8819\,
            I => \N__8732\
        );

    \I__2037\ : ClkMux
    port map (
            O => \N__8818\,
            I => \N__8732\
        );

    \I__2036\ : ClkMux
    port map (
            O => \N__8817\,
            I => \N__8732\
        );

    \I__2035\ : ClkMux
    port map (
            O => \N__8816\,
            I => \N__8732\
        );

    \I__2034\ : ClkMux
    port map (
            O => \N__8815\,
            I => \N__8732\
        );

    \I__2033\ : ClkMux
    port map (
            O => \N__8814\,
            I => \N__8732\
        );

    \I__2032\ : ClkMux
    port map (
            O => \N__8813\,
            I => \N__8732\
        );

    \I__2031\ : Glb2LocalMux
    port map (
            O => \N__8810\,
            I => \N__8732\
        );

    \I__2030\ : ClkMux
    port map (
            O => \N__8809\,
            I => \N__8732\
        );

    \I__2029\ : ClkMux
    port map (
            O => \N__8808\,
            I => \N__8732\
        );

    \I__2028\ : ClkMux
    port map (
            O => \N__8807\,
            I => \N__8732\
        );

    \I__2027\ : ClkMux
    port map (
            O => \N__8806\,
            I => \N__8732\
        );

    \I__2026\ : ClkMux
    port map (
            O => \N__8805\,
            I => \N__8732\
        );

    \I__2025\ : ClkMux
    port map (
            O => \N__8804\,
            I => \N__8732\
        );

    \I__2024\ : ClkMux
    port map (
            O => \N__8803\,
            I => \N__8732\
        );

    \I__2023\ : ClkMux
    port map (
            O => \N__8802\,
            I => \N__8732\
        );

    \I__2022\ : ClkMux
    port map (
            O => \N__8801\,
            I => \N__8732\
        );

    \I__2021\ : GlobalMux
    port map (
            O => \N__8732\,
            I => \CLK80_PLL\
        );

    \I__2020\ : CEMux
    port map (
            O => \N__8729\,
            I => \N__8726\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__8726\,
            I => \N__8721\
        );

    \I__2018\ : CEMux
    port map (
            O => \N__8725\,
            I => \N__8718\
        );

    \I__2017\ : CEMux
    port map (
            O => \N__8724\,
            I => \N__8715\
        );

    \I__2016\ : Span4Mux_h
    port map (
            O => \N__8721\,
            I => \N__8712\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__8718\,
            I => \N__8708\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__8715\,
            I => \N__8705\
        );

    \I__2013\ : Span4Mux_h
    port map (
            O => \N__8712\,
            I => \N__8700\
        );

    \I__2012\ : CEMux
    port map (
            O => \N__8711\,
            I => \N__8697\
        );

    \I__2011\ : Span12Mux_h
    port map (
            O => \N__8708\,
            I => \N__8692\
        );

    \I__2010\ : Sp12to4
    port map (
            O => \N__8705\,
            I => \N__8692\
        );

    \I__2009\ : CEMux
    port map (
            O => \N__8704\,
            I => \N__8689\
        );

    \I__2008\ : CEMux
    port map (
            O => \N__8703\,
            I => \N__8686\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__8700\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__8697\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2005\ : Odrv12
    port map (
            O => \N__8692\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__8689\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__8686\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2002\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__8672\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2000\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8663\
        );

    \I__1999\ : InMux
    port map (
            O => \N__8668\,
            I => \N__8663\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__1997\ : Odrv4
    port map (
            O => \N__8660\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1996\ : InMux
    port map (
            O => \N__8657\,
            I => \N__8654\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__8654\,
            I => \N__8650\
        );

    \I__1994\ : InMux
    port map (
            O => \N__8653\,
            I => \N__8647\
        );

    \I__1993\ : Span4Mux_h
    port map (
            O => \N__8650\,
            I => \N__8642\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__8647\,
            I => \N__8642\
        );

    \I__1991\ : Sp12to4
    port map (
            O => \N__8642\,
            I => \N__8639\
        );

    \I__1990\ : Span12Mux_v
    port map (
            O => \N__8639\,
            I => \N__8636\
        );

    \I__1989\ : Span12Mux_h
    port map (
            O => \N__8636\,
            I => \N__8633\
        );

    \I__1988\ : Odrv12
    port map (
            O => \N__8633\,
            I => \DRA_c_5\
        );

    \I__1987\ : InMux
    port map (
            O => \N__8630\,
            I => \N__8627\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__1985\ : Span4Mux_h
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__1984\ : Odrv4
    port map (
            O => \N__8621\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1983\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8614\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8617\,
            I => \N__8611\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__8614\,
            I => \N__8606\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__8611\,
            I => \N__8606\
        );

    \I__1979\ : Span4Mux_v
    port map (
            O => \N__8606\,
            I => \N__8603\
        );

    \I__1978\ : Sp12to4
    port map (
            O => \N__8603\,
            I => \N__8600\
        );

    \I__1977\ : Span12Mux_h
    port map (
            O => \N__8600\,
            I => \N__8597\
        );

    \I__1976\ : Odrv12
    port map (
            O => \N__8597\,
            I => \DRA_c_7\
        );

    \I__1975\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8591\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__8591\,
            I => \N__8588\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__8588\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1972\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8582\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__8582\,
            I => \N__8579\
        );

    \I__1970\ : Span4Mux_h
    port map (
            O => \N__8579\,
            I => \N__8576\
        );

    \I__1969\ : Odrv4
    port map (
            O => \N__8576\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1968\ : InMux
    port map (
            O => \N__8573\,
            I => \N__8570\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__8570\,
            I => \N__8567\
        );

    \I__1966\ : Span4Mux_h
    port map (
            O => \N__8567\,
            I => \N__8564\
        );

    \I__1965\ : Span4Mux_v
    port map (
            O => \N__8564\,
            I => \N__8561\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__8561\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8554\
        );

    \I__1962\ : InMux
    port map (
            O => \N__8557\,
            I => \N__8551\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__8554\,
            I => \N__8546\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__8551\,
            I => \N__8546\
        );

    \I__1959\ : Sp12to4
    port map (
            O => \N__8546\,
            I => \N__8543\
        );

    \I__1958\ : Span12Mux_v
    port map (
            O => \N__8543\,
            I => \N__8540\
        );

    \I__1957\ : Span12Mux_h
    port map (
            O => \N__8540\,
            I => \N__8537\
        );

    \I__1956\ : Odrv12
    port map (
            O => \N__8537\,
            I => \DRA_c_1\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__8531\,
            I => \N__8528\
        );

    \I__1953\ : Span4Mux_v
    port map (
            O => \N__8528\,
            I => \N__8525\
        );

    \I__1952\ : Span4Mux_h
    port map (
            O => \N__8525\,
            I => \N__8522\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__8522\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8514\
        );

    \I__1949\ : InMux
    port map (
            O => \N__8518\,
            I => \N__8511\
        );

    \I__1948\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8508\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__8514\,
            I => \N__8503\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__8511\,
            I => \N__8503\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__8508\,
            I => \N__8500\
        );

    \I__1944\ : Span4Mux_v
    port map (
            O => \N__8503\,
            I => \N__8497\
        );

    \I__1943\ : Span4Mux_v
    port map (
            O => \N__8500\,
            I => \N__8494\
        );

    \I__1942\ : Sp12to4
    port map (
            O => \N__8497\,
            I => \N__8489\
        );

    \I__1941\ : Sp12to4
    port map (
            O => \N__8494\,
            I => \N__8489\
        );

    \I__1940\ : Span12Mux_h
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__1939\ : Span12Mux_v
    port map (
            O => \N__8486\,
            I => \N__8483\
        );

    \I__1938\ : Odrv12
    port map (
            O => \N__8483\,
            I => \DBRn_c\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8477\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8477\,
            I => \N__8467\
        );

    \I__1935\ : ClkMux
    port map (
            O => \N__8476\,
            I => \N__8450\
        );

    \I__1934\ : ClkMux
    port map (
            O => \N__8475\,
            I => \N__8450\
        );

    \I__1933\ : ClkMux
    port map (
            O => \N__8474\,
            I => \N__8450\
        );

    \I__1932\ : ClkMux
    port map (
            O => \N__8473\,
            I => \N__8450\
        );

    \I__1931\ : ClkMux
    port map (
            O => \N__8472\,
            I => \N__8450\
        );

    \I__1930\ : ClkMux
    port map (
            O => \N__8471\,
            I => \N__8450\
        );

    \I__1929\ : ClkMux
    port map (
            O => \N__8470\,
            I => \N__8450\
        );

    \I__1928\ : Glb2LocalMux
    port map (
            O => \N__8467\,
            I => \N__8450\
        );

    \I__1927\ : GlobalMux
    port map (
            O => \N__8450\,
            I => \N__8447\
        );

    \I__1926\ : gio2CtrlBuf
    port map (
            O => \N__8447\,
            I => \C1_c_g\
        );

    \I__1925\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8440\
        );

    \I__1924\ : InMux
    port map (
            O => \N__8443\,
            I => \N__8430\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__8440\,
            I => \N__8426\
        );

    \I__1922\ : InMux
    port map (
            O => \N__8439\,
            I => \N__8417\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8417\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8417\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8436\,
            I => \N__8417\
        );

    \I__1918\ : InMux
    port map (
            O => \N__8435\,
            I => \N__8414\
        );

    \I__1917\ : InMux
    port map (
            O => \N__8434\,
            I => \N__8411\
        );

    \I__1916\ : InMux
    port map (
            O => \N__8433\,
            I => \N__8408\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__8430\,
            I => \N__8405\
        );

    \I__1914\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8402\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__8426\,
            I => \N__8395\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__8417\,
            I => \N__8395\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__8414\,
            I => \N__8395\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__8411\,
            I => \N__8391\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__8408\,
            I => \N__8388\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__8405\,
            I => \N__8385\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8402\,
            I => \N__8380\
        );

    \I__1906\ : Span4Mux_v
    port map (
            O => \N__8395\,
            I => \N__8380\
        );

    \I__1905\ : InMux
    port map (
            O => \N__8394\,
            I => \N__8377\
        );

    \I__1904\ : Span12Mux_v
    port map (
            O => \N__8391\,
            I => \N__8374\
        );

    \I__1903\ : Span12Mux_v
    port map (
            O => \N__8388\,
            I => \N__8365\
        );

    \I__1902\ : Sp12to4
    port map (
            O => \N__8385\,
            I => \N__8365\
        );

    \I__1901\ : Sp12to4
    port map (
            O => \N__8380\,
            I => \N__8365\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__8377\,
            I => \N__8365\
        );

    \I__1899\ : Span12Mux_h
    port map (
            O => \N__8374\,
            I => \N__8362\
        );

    \I__1898\ : Span12Mux_h
    port map (
            O => \N__8365\,
            I => \N__8359\
        );

    \I__1897\ : Odrv12
    port map (
            O => \N__8362\,
            I => \RESETn_c\
        );

    \I__1896\ : Odrv12
    port map (
            O => \N__8359\,
            I => \RESETn_c\
        );

    \I__1895\ : IoInMux
    port map (
            O => \N__8354\,
            I => \N__8351\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__8351\,
            I => \N__8348\
        );

    \I__1893\ : Span12Mux_s4_v
    port map (
            O => \N__8348\,
            I => \N__8345\
        );

    \I__1892\ : Odrv12
    port map (
            O => \N__8345\,
            I => \RESETn_c_i\
        );

    \I__1891\ : IoInMux
    port map (
            O => \N__8342\,
            I => \N__8339\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__8339\,
            I => \N__8336\
        );

    \I__1889\ : Span12Mux_s10_v
    port map (
            O => \N__8336\,
            I => \N__8333\
        );

    \I__1888\ : Span12Mux_h
    port map (
            O => \N__8333\,
            I => \N__8330\
        );

    \I__1887\ : Odrv12
    port map (
            O => \N__8330\,
            I => \N_118\
        );

    \I__1886\ : InMux
    port map (
            O => \N__8327\,
            I => \N__8319\
        );

    \I__1885\ : InMux
    port map (
            O => \N__8326\,
            I => \N__8319\
        );

    \I__1884\ : InMux
    port map (
            O => \N__8325\,
            I => \N__8314\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8324\,
            I => \N__8314\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__8319\,
            I => \N__8309\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__8314\,
            I => \N__8306\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8313\,
            I => \N__8301\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8312\,
            I => \N__8301\
        );

    \I__1878\ : Span4Mux_v
    port map (
            O => \N__8309\,
            I => \N__8298\
        );

    \I__1877\ : Span4Mux_v
    port map (
            O => \N__8306\,
            I => \N__8295\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8301\,
            I => \N__8292\
        );

    \I__1875\ : Span4Mux_h
    port map (
            O => \N__8298\,
            I => \N__8289\
        );

    \I__1874\ : Span4Mux_h
    port map (
            O => \N__8295\,
            I => \N__8284\
        );

    \I__1873\ : Span4Mux_v
    port map (
            O => \N__8292\,
            I => \N__8284\
        );

    \I__1872\ : Sp12to4
    port map (
            O => \N__8289\,
            I => \N__8279\
        );

    \I__1871\ : Sp12to4
    port map (
            O => \N__8284\,
            I => \N__8279\
        );

    \I__1870\ : Odrv12
    port map (
            O => \N__8279\,
            I => \A_c_0\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8276\,
            I => \N__8272\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__8275\,
            I => \N__8269\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8272\,
            I => \N__8265\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8269\,
            I => \N__8260\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8268\,
            I => \N__8260\
        );

    \I__1864\ : Span4Mux_h
    port map (
            O => \N__8265\,
            I => \N__8257\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__8260\,
            I => \N__8254\
        );

    \I__1862\ : Sp12to4
    port map (
            O => \N__8257\,
            I => \N__8251\
        );

    \I__1861\ : Span12Mux_v
    port map (
            O => \N__8254\,
            I => \N__8248\
        );

    \I__1860\ : Span12Mux_v
    port map (
            O => \N__8251\,
            I => \N__8245\
        );

    \I__1859\ : Span12Mux_h
    port map (
            O => \N__8248\,
            I => \N__8242\
        );

    \I__1858\ : Odrv12
    port map (
            O => \N__8245\,
            I => \SIZ_c_0\
        );

    \I__1857\ : Odrv12
    port map (
            O => \N__8242\,
            I => \SIZ_c_0\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8237\,
            I => \N__8231\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8231\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8231\,
            I => \N__8228\
        );

    \I__1853\ : Span12Mux_s9_v
    port map (
            O => \N__8228\,
            I => \N__8224\
        );

    \I__1852\ : InMux
    port map (
            O => \N__8227\,
            I => \N__8221\
        );

    \I__1851\ : Odrv12
    port map (
            O => \N__8224\,
            I => \DS_ENm\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8221\,
            I => \DS_ENm\
        );

    \I__1849\ : IoInMux
    port map (
            O => \N__8216\,
            I => \N__8213\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8213\,
            I => \N__8210\
        );

    \I__1847\ : Span4Mux_s3_v
    port map (
            O => \N__8210\,
            I => \N__8207\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__8207\,
            I => \N__8204\
        );

    \I__1845\ : Sp12to4
    port map (
            O => \N__8204\,
            I => \N__8201\
        );

    \I__1844\ : Odrv12
    port map (
            O => \N__8201\,
            I => \N_113\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8198\,
            I => \N__8195\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__8195\,
            I => \N__8191\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8194\,
            I => \N__8188\
        );

    \I__1840\ : Span4Mux_v
    port map (
            O => \N__8191\,
            I => \N__8182\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8188\,
            I => \N__8182\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__8187\,
            I => \N__8178\
        );

    \I__1837\ : Span4Mux_v
    port map (
            O => \N__8182\,
            I => \N__8175\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8181\,
            I => \N__8172\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8178\,
            I => \N__8169\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__8175\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__8172\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8169\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1831\ : IoInMux
    port map (
            O => \N__8162\,
            I => \N__8159\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8159\,
            I => \N__8156\
        );

    \I__1829\ : Span4Mux_s2_v
    port map (
            O => \N__8156\,
            I => \N__8153\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__8153\,
            I => \N__8150\
        );

    \I__1827\ : Span4Mux_h
    port map (
            O => \N__8150\,
            I => \N__8147\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__8147\,
            I => \CRCSn_c\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__8144\,
            I => \N__8141\
        );

    \I__1824\ : InMux
    port map (
            O => \N__8141\,
            I => \N__8137\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8140\,
            I => \N__8134\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__8137\,
            I => \N__8128\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8134\,
            I => \N__8123\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8133\,
            I => \N__8118\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8132\,
            I => \N__8118\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8115\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__8128\,
            I => \N__8112\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8127\,
            I => \N__8107\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8126\,
            I => \N__8107\
        );

    \I__1814\ : Span4Mux_h
    port map (
            O => \N__8123\,
            I => \N__8102\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8118\,
            I => \N__8102\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8115\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__8112\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8107\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__8102\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1808\ : IoInMux
    port map (
            O => \N__8093\,
            I => \N__8090\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8090\,
            I => \N__8087\
        );

    \I__1806\ : IoSpan4Mux
    port map (
            O => \N__8087\,
            I => \N__8084\
        );

    \I__1805\ : Span4Mux_s2_h
    port map (
            O => \N__8084\,
            I => \N__8081\
        );

    \I__1804\ : Sp12to4
    port map (
            O => \N__8081\,
            I => \N__8078\
        );

    \I__1803\ : Span12Mux_h
    port map (
            O => \N__8078\,
            I => \N__8075\
        );

    \I__1802\ : Odrv12
    port map (
            O => \N__8075\,
            I => \WEn_c\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8072\,
            I => \N__8068\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8071\,
            I => \N__8065\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8068\,
            I => \N__8060\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8065\,
            I => \N__8057\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8052\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8063\,
            I => \N__8052\
        );

    \I__1795\ : Span4Mux_v
    port map (
            O => \N__8060\,
            I => \N__8047\
        );

    \I__1794\ : Span4Mux_v
    port map (
            O => \N__8057\,
            I => \N__8042\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8052\,
            I => \N__8042\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8051\,
            I => \N__8037\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8050\,
            I => \N__8037\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__8047\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1789\ : Odrv4
    port map (
            O => \N__8042\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8037\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1787\ : IoInMux
    port map (
            O => \N__8030\,
            I => \N__8027\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8027\,
            I => \N__8024\
        );

    \I__1785\ : Span4Mux_s2_v
    port map (
            O => \N__8024\,
            I => \N__8021\
        );

    \I__1784\ : Span4Mux_v
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__1782\ : Span4Mux_h
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__8012\,
            I => \RASn_c\
        );

    \I__1780\ : InMux
    port map (
            O => \N__8009\,
            I => \N__8006\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8006\,
            I => \N__8003\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__8003\,
            I => \N__8000\
        );

    \I__1777\ : Span4Mux_v
    port map (
            O => \N__8000\,
            I => \N__7997\
        );

    \I__1776\ : Sp12to4
    port map (
            O => \N__7997\,
            I => \N__7994\
        );

    \I__1775\ : Span12Mux_h
    port map (
            O => \N__7994\,
            I => \N__7991\
        );

    \I__1774\ : Odrv12
    port map (
            O => \N__7991\,
            I => \A_c_19\
        );

    \I__1773\ : IoInMux
    port map (
            O => \N__7988\,
            I => \N__7985\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__7985\,
            I => \N__7982\
        );

    \I__1771\ : IoSpan4Mux
    port map (
            O => \N__7982\,
            I => \N__7979\
        );

    \I__1770\ : Span4Mux_s1_h
    port map (
            O => \N__7979\,
            I => \N__7976\
        );

    \I__1769\ : Sp12to4
    port map (
            O => \N__7976\,
            I => \N__7973\
        );

    \I__1768\ : Span12Mux_h
    port map (
            O => \N__7973\,
            I => \N__7970\
        );

    \I__1767\ : Odrv12
    port map (
            O => \N__7970\,
            I => \CMA_c_9\
        );

    \I__1766\ : InMux
    port map (
            O => \N__7967\,
            I => \N__7960\
        );

    \I__1765\ : InMux
    port map (
            O => \N__7966\,
            I => \N__7960\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__7965\,
            I => \N__7957\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__7960\,
            I => \N__7953\
        );

    \I__1762\ : InMux
    port map (
            O => \N__7957\,
            I => \N__7948\
        );

    \I__1761\ : InMux
    port map (
            O => \N__7956\,
            I => \N__7948\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__7953\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__7948\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1758\ : InMux
    port map (
            O => \N__7943\,
            I => \N__7940\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__7940\,
            I => \N__7937\
        );

    \I__1756\ : Span4Mux_v
    port map (
            O => \N__7937\,
            I => \N__7934\
        );

    \I__1755\ : Span4Mux_v
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__1754\ : Sp12to4
    port map (
            O => \N__7931\,
            I => \N__7928\
        );

    \I__1753\ : Span12Mux_h
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__1752\ : Odrv12
    port map (
            O => \N__7925\,
            I => \A_c_17\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__7922\,
            I => \N__7915\
        );

    \I__1750\ : InMux
    port map (
            O => \N__7921\,
            I => \N__7907\
        );

    \I__1749\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7904\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__7919\,
            I => \N__7899\
        );

    \I__1747\ : InMux
    port map (
            O => \N__7918\,
            I => \N__7891\
        );

    \I__1746\ : InMux
    port map (
            O => \N__7915\,
            I => \N__7891\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__7914\,
            I => \N__7881\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__7913\,
            I => \N__7878\
        );

    \I__1743\ : InMux
    port map (
            O => \N__7912\,
            I => \N__7875\
        );

    \I__1742\ : InMux
    port map (
            O => \N__7911\,
            I => \N__7870\
        );

    \I__1741\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7870\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__7907\,
            I => \N__7865\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__7904\,
            I => \N__7865\
        );

    \I__1738\ : InMux
    port map (
            O => \N__7903\,
            I => \N__7858\
        );

    \I__1737\ : InMux
    port map (
            O => \N__7902\,
            I => \N__7858\
        );

    \I__1736\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7858\
        );

    \I__1735\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7853\
        );

    \I__1734\ : InMux
    port map (
            O => \N__7897\,
            I => \N__7853\
        );

    \I__1733\ : InMux
    port map (
            O => \N__7896\,
            I => \N__7850\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__7891\,
            I => \N__7847\
        );

    \I__1731\ : InMux
    port map (
            O => \N__7890\,
            I => \N__7840\
        );

    \I__1730\ : InMux
    port map (
            O => \N__7889\,
            I => \N__7840\
        );

    \I__1729\ : InMux
    port map (
            O => \N__7888\,
            I => \N__7840\
        );

    \I__1728\ : InMux
    port map (
            O => \N__7887\,
            I => \N__7837\
        );

    \I__1727\ : InMux
    port map (
            O => \N__7886\,
            I => \N__7832\
        );

    \I__1726\ : InMux
    port map (
            O => \N__7885\,
            I => \N__7832\
        );

    \I__1725\ : InMux
    port map (
            O => \N__7884\,
            I => \N__7825\
        );

    \I__1724\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7825\
        );

    \I__1723\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7825\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__7875\,
            I => \N__7819\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__7870\,
            I => \N__7819\
        );

    \I__1720\ : Span4Mux_v
    port map (
            O => \N__7865\,
            I => \N__7812\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__7858\,
            I => \N__7812\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__7853\,
            I => \N__7812\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__7850\,
            I => \N__7808\
        );

    \I__1716\ : Span4Mux_v
    port map (
            O => \N__7847\,
            I => \N__7801\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__7840\,
            I => \N__7801\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__7837\,
            I => \N__7801\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__7832\,
            I => \N__7798\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__7825\,
            I => \N__7795\
        );

    \I__1711\ : InMux
    port map (
            O => \N__7824\,
            I => \N__7792\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__7819\,
            I => \N__7789\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__7812\,
            I => \N__7786\
        );

    \I__1708\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7783\
        );

    \I__1707\ : Span4Mux_v
    port map (
            O => \N__7808\,
            I => \N__7778\
        );

    \I__1706\ : Span4Mux_h
    port map (
            O => \N__7801\,
            I => \N__7778\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__7798\,
            I => \CPU_CYCLEm\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__7795\,
            I => \CPU_CYCLEm\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__7792\,
            I => \CPU_CYCLEm\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__7789\,
            I => \CPU_CYCLEm\
        );

    \I__1701\ : Odrv4
    port map (
            O => \N__7786\,
            I => \CPU_CYCLEm\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__7783\,
            I => \CPU_CYCLEm\
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__7778\,
            I => \CPU_CYCLEm\
        );

    \I__1698\ : IoInMux
    port map (
            O => \N__7763\,
            I => \N__7760\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__7760\,
            I => \N__7757\
        );

    \I__1696\ : IoSpan4Mux
    port map (
            O => \N__7757\,
            I => \N__7754\
        );

    \I__1695\ : Span4Mux_s2_h
    port map (
            O => \N__7754\,
            I => \N__7751\
        );

    \I__1694\ : Sp12to4
    port map (
            O => \N__7751\,
            I => \N__7748\
        );

    \I__1693\ : Span12Mux_h
    port map (
            O => \N__7748\,
            I => \N__7745\
        );

    \I__1692\ : Odrv12
    port map (
            O => \N__7745\,
            I => \CMA_c_8\
        );

    \I__1691\ : InMux
    port map (
            O => \N__7742\,
            I => \N__7738\
        );

    \I__1690\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7735\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__7738\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__7735\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__7730\,
            I => \N__7726\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__7729\,
            I => \N__7722\
        );

    \I__1685\ : InMux
    port map (
            O => \N__7726\,
            I => \N__7717\
        );

    \I__1684\ : InMux
    port map (
            O => \N__7725\,
            I => \N__7717\
        );

    \I__1683\ : InMux
    port map (
            O => \N__7722\,
            I => \N__7714\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__7717\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__7714\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1680\ : IoInMux
    port map (
            O => \N__7709\,
            I => \N__7705\
        );

    \I__1679\ : IoInMux
    port map (
            O => \N__7708\,
            I => \N__7702\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__7705\,
            I => \N__7699\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__7702\,
            I => \N__7696\
        );

    \I__1676\ : Span4Mux_s3_v
    port map (
            O => \N__7699\,
            I => \N__7693\
        );

    \I__1675\ : Span4Mux_s2_v
    port map (
            O => \N__7696\,
            I => \N__7690\
        );

    \I__1674\ : Sp12to4
    port map (
            O => \N__7693\,
            I => \N__7687\
        );

    \I__1673\ : Span4Mux_h
    port map (
            O => \N__7690\,
            I => \N__7684\
        );

    \I__1672\ : Span12Mux_s11_h
    port map (
            O => \N__7687\,
            I => \N__7681\
        );

    \I__1671\ : Sp12to4
    port map (
            O => \N__7684\,
            I => \N__7678\
        );

    \I__1670\ : Span12Mux_v
    port map (
            O => \N__7681\,
            I => \N__7672\
        );

    \I__1669\ : Span12Mux_v
    port map (
            O => \N__7678\,
            I => \N__7672\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7677\,
            I => \N__7669\
        );

    \I__1667\ : Odrv12
    port map (
            O => \N__7672\,
            I => \ASn_c\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__7669\,
            I => \ASn_c\
        );

    \I__1665\ : InMux
    port map (
            O => \N__7664\,
            I => \N__7652\
        );

    \I__1664\ : InMux
    port map (
            O => \N__7663\,
            I => \N__7652\
        );

    \I__1663\ : InMux
    port map (
            O => \N__7662\,
            I => \N__7652\
        );

    \I__1662\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7652\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__7652\,
            I => \U712_REG_SM.STATE_COUNT_RNITQLC2Z0Z_1\
        );

    \I__1660\ : InMux
    port map (
            O => \N__7649\,
            I => \N__7646\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__7643\,
            I => \N__7640\
        );

    \I__1657\ : Sp12to4
    port map (
            O => \N__7640\,
            I => \N__7637\
        );

    \I__1656\ : Span12Mux_h
    port map (
            O => \N__7637\,
            I => \N__7634\
        );

    \I__1655\ : Span12Mux_v
    port map (
            O => \N__7634\,
            I => \N__7631\
        );

    \I__1654\ : Odrv12
    port map (
            O => \N__7631\,
            I => \REGSPACEn_c\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__7628\,
            I => \N__7624\
        );

    \I__1652\ : InMux
    port map (
            O => \N__7627\,
            I => \N__7619\
        );

    \I__1651\ : InMux
    port map (
            O => \N__7624\,
            I => \N__7619\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__7619\,
            I => \U712_REG_SM.REG_CYCLE_GOZ0\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__7616\,
            I => \N__7612\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7615\,
            I => \N__7609\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7606\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__7609\,
            I => \N__7603\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__7606\,
            I => \N__7600\
        );

    \I__1644\ : Span4Mux_v
    port map (
            O => \N__7603\,
            I => \N__7597\
        );

    \I__1643\ : Span4Mux_v
    port map (
            O => \N__7600\,
            I => \N__7594\
        );

    \I__1642\ : Sp12to4
    port map (
            O => \N__7597\,
            I => \N__7589\
        );

    \I__1641\ : Sp12to4
    port map (
            O => \N__7594\,
            I => \N__7589\
        );

    \I__1640\ : Span12Mux_h
    port map (
            O => \N__7589\,
            I => \N__7586\
        );

    \I__1639\ : Span12Mux_v
    port map (
            O => \N__7586\,
            I => \N__7583\
        );

    \I__1638\ : Odrv12
    port map (
            O => \N__7583\,
            I => \TSn_c\
        );

    \I__1637\ : InMux
    port map (
            O => \N__7580\,
            I => \N__7568\
        );

    \I__1636\ : InMux
    port map (
            O => \N__7579\,
            I => \N__7568\
        );

    \I__1635\ : InMux
    port map (
            O => \N__7578\,
            I => \N__7568\
        );

    \I__1634\ : InMux
    port map (
            O => \N__7577\,
            I => \N__7568\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7568\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__7565\,
            I => \N__7561\
        );

    \I__1631\ : InMux
    port map (
            O => \N__7564\,
            I => \N__7556\
        );

    \I__1630\ : InMux
    port map (
            O => \N__7561\,
            I => \N__7553\
        );

    \I__1629\ : InMux
    port map (
            O => \N__7560\,
            I => \N__7548\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7559\,
            I => \N__7548\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__7556\,
            I => \N__7545\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__7553\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__7548\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa\
        );

    \I__1624\ : Odrv12
    port map (
            O => \N__7545\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa\
        );

    \I__1623\ : InMux
    port map (
            O => \N__7538\,
            I => \N__7529\
        );

    \I__1622\ : InMux
    port map (
            O => \N__7537\,
            I => \N__7529\
        );

    \I__1621\ : InMux
    port map (
            O => \N__7536\,
            I => \N__7529\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__7529\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__7526\,
            I => \N__7521\
        );

    \I__1618\ : InMux
    port map (
            O => \N__7525\,
            I => \N__7514\
        );

    \I__1617\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7514\
        );

    \I__1616\ : InMux
    port map (
            O => \N__7521\,
            I => \N__7514\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__7514\,
            I => \U712_REG_SM.N_205\
        );

    \I__1614\ : InMux
    port map (
            O => \N__7511\,
            I => \N__7507\
        );

    \I__1613\ : InMux
    port map (
            O => \N__7510\,
            I => \N__7503\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__7507\,
            I => \N__7500\
        );

    \I__1611\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7497\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__7503\,
            I => \U712_REG_SM.N_202\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__7500\,
            I => \U712_REG_SM.N_202\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__7497\,
            I => \U712_REG_SM.N_202\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__7490\,
            I => \N__7485\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7489\,
            I => \N__7482\
        );

    \I__1605\ : InMux
    port map (
            O => \N__7488\,
            I => \N__7479\
        );

    \I__1604\ : InMux
    port map (
            O => \N__7485\,
            I => \N__7476\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__7482\,
            I => \N__7473\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__7479\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__7476\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1600\ : Odrv12
    port map (
            O => \N__7473\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7466\,
            I => \N__7461\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__7465\,
            I => \N__7458\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__7464\,
            I => \N__7455\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__7461\,
            I => \N__7442\
        );

    \I__1595\ : InMux
    port map (
            O => \N__7458\,
            I => \N__7439\
        );

    \I__1594\ : InMux
    port map (
            O => \N__7455\,
            I => \N__7436\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__7454\,
            I => \N__7433\
        );

    \I__1592\ : InMux
    port map (
            O => \N__7453\,
            I => \N__7428\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7452\,
            I => \N__7425\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7451\,
            I => \N__7416\
        );

    \I__1589\ : InMux
    port map (
            O => \N__7450\,
            I => \N__7416\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7449\,
            I => \N__7416\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7448\,
            I => \N__7416\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7447\,
            I => \N__7413\
        );

    \I__1585\ : CascadeMux
    port map (
            O => \N__7446\,
            I => \N__7410\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__7445\,
            I => \N__7407\
        );

    \I__1583\ : Span4Mux_v
    port map (
            O => \N__7442\,
            I => \N__7400\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7439\,
            I => \N__7400\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__7436\,
            I => \N__7400\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7433\,
            I => \N__7397\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7432\,
            I => \N__7392\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__7431\,
            I => \N__7388\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7428\,
            I => \N__7383\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__7425\,
            I => \N__7380\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7416\,
            I => \N__7377\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__7413\,
            I => \N__7374\
        );

    \I__1573\ : InMux
    port map (
            O => \N__7410\,
            I => \N__7369\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7407\,
            I => \N__7369\
        );

    \I__1571\ : Span4Mux_h
    port map (
            O => \N__7400\,
            I => \N__7363\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__7397\,
            I => \N__7360\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7396\,
            I => \N__7355\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7395\,
            I => \N__7355\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__7392\,
            I => \N__7352\
        );

    \I__1566\ : InMux
    port map (
            O => \N__7391\,
            I => \N__7349\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7388\,
            I => \N__7342\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7387\,
            I => \N__7342\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7342\
        );

    \I__1562\ : Span4Mux_v
    port map (
            O => \N__7383\,
            I => \N__7331\
        );

    \I__1561\ : Span4Mux_v
    port map (
            O => \N__7380\,
            I => \N__7331\
        );

    \I__1560\ : Span4Mux_v
    port map (
            O => \N__7377\,
            I => \N__7331\
        );

    \I__1559\ : Span4Mux_h
    port map (
            O => \N__7374\,
            I => \N__7331\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7369\,
            I => \N__7331\
        );

    \I__1557\ : InMux
    port map (
            O => \N__7368\,
            I => \N__7324\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7367\,
            I => \N__7324\
        );

    \I__1555\ : InMux
    port map (
            O => \N__7366\,
            I => \N__7324\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__7363\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__7360\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7355\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__7352\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7349\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7342\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__7331\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7324\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7307\,
            I => \N__7303\
        );

    \I__1545\ : InMux
    port map (
            O => \N__7306\,
            I => \N__7300\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7303\,
            I => \N__7291\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__7300\,
            I => \N__7291\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7299\,
            I => \N__7286\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7298\,
            I => \N__7286\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7297\,
            I => \N__7281\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7296\,
            I => \N__7281\
        );

    \I__1538\ : Odrv4
    port map (
            O => \N__7291\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__7286\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__7281\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7274\,
            I => \N__7271\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7271\,
            I => \N__7268\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__7268\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7265\,
            I => \N__7262\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__7262\,
            I => \N__7259\
        );

    \I__1530\ : Span4Mux_h
    port map (
            O => \N__7259\,
            I => \N__7256\
        );

    \I__1529\ : Odrv4
    port map (
            O => \N__7256\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__1528\ : IoInMux
    port map (
            O => \N__7253\,
            I => \N__7249\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7252\,
            I => \N__7246\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__7249\,
            I => \N__7243\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7246\,
            I => \N__7240\
        );

    \I__1524\ : IoSpan4Mux
    port map (
            O => \N__7243\,
            I => \N__7237\
        );

    \I__1523\ : Span12Mux_v
    port map (
            O => \N__7240\,
            I => \N__7234\
        );

    \I__1522\ : IoSpan4Mux
    port map (
            O => \N__7237\,
            I => \N__7231\
        );

    \I__1521\ : Span12Mux_h
    port map (
            O => \N__7234\,
            I => \N__7228\
        );

    \I__1520\ : IoSpan4Mux
    port map (
            O => \N__7231\,
            I => \N__7225\
        );

    \I__1519\ : Odrv12
    port map (
            O => \N__7228\,
            I => \C3_c\
        );

    \I__1518\ : Odrv4
    port map (
            O => \N__7225\,
            I => \C3_c\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7220\,
            I => \N__7211\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7219\,
            I => \N__7211\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7218\,
            I => \N__7211\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__7211\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__1513\ : IoInMux
    port map (
            O => \N__7208\,
            I => \N__7204\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7207\,
            I => \N__7201\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7204\,
            I => \N__7198\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7201\,
            I => \N__7195\
        );

    \I__1509\ : Span4Mux_s3_h
    port map (
            O => \N__7198\,
            I => \N__7192\
        );

    \I__1508\ : Span12Mux_v
    port map (
            O => \N__7195\,
            I => \N__7189\
        );

    \I__1507\ : Sp12to4
    port map (
            O => \N__7192\,
            I => \N__7186\
        );

    \I__1506\ : Span12Mux_h
    port map (
            O => \N__7189\,
            I => \N__7183\
        );

    \I__1505\ : Span12Mux_v
    port map (
            O => \N__7186\,
            I => \N__7180\
        );

    \I__1504\ : Odrv12
    port map (
            O => \N__7183\,
            I => \C1_c\
        );

    \I__1503\ : Odrv12
    port map (
            O => \N__7180\,
            I => \C1_c\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__7175\,
            I => \N__7170\
        );

    \I__1501\ : CascadeMux
    port map (
            O => \N__7174\,
            I => \N__7167\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7163\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7170\,
            I => \N__7160\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7155\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7166\,
            I => \N__7155\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__7163\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7160\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7155\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7148\,
            I => \N__7142\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7147\,
            I => \N__7142\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7142\,
            I => \N__7135\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7141\,
            I => \N__7132\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7129\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7124\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7138\,
            I => \N__7124\
        );

    \I__1486\ : Sp12to4
    port map (
            O => \N__7135\,
            I => \N__7121\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7132\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7129\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7124\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1482\ : Odrv12
    port map (
            O => \N__7121\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7112\,
            I => \N__7101\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7111\,
            I => \N__7101\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7110\,
            I => \N__7101\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7109\,
            I => \N__7096\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7108\,
            I => \N__7096\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7101\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__7096\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7091\,
            I => \N__7085\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7090\,
            I => \N__7078\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7089\,
            I => \N__7078\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7088\,
            I => \N__7078\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7085\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7078\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__7073\,
            I => \N__7067\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7072\,
            I => \N__7064\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7071\,
            I => \N__7057\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7057\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7067\,
            I => \N__7057\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7064\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7057\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7052\,
            I => \N__7048\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7051\,
            I => \N__7045\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7048\,
            I => \N__7042\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7045\,
            I => \N__7039\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__7042\,
            I => \U712_REG_SM.N_210\
        );

    \I__1456\ : Odrv4
    port map (
            O => \N__7039\,
            I => \U712_REG_SM.N_210\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7034\,
            I => \N__7025\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7033\,
            I => \N__7025\
        );

    \I__1453\ : InMux
    port map (
            O => \N__7032\,
            I => \N__7025\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__7025\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1451\ : CascadeMux
    port map (
            O => \N__7022\,
            I => \N__7018\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7021\,
            I => \N__7015\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7018\,
            I => \N__7012\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7015\,
            I => \N__7005\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7012\,
            I => \N__7005\
        );

    \I__1446\ : InMux
    port map (
            O => \N__7011\,
            I => \N__7000\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7010\,
            I => \N__7000\
        );

    \I__1444\ : Span4Mux_v
    port map (
            O => \N__7005\,
            I => \N__6997\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7000\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__6997\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__6992\,
            I => \N__6989\
        );

    \I__1440\ : InMux
    port map (
            O => \N__6989\,
            I => \N__6980\
        );

    \I__1439\ : InMux
    port map (
            O => \N__6988\,
            I => \N__6980\
        );

    \I__1438\ : InMux
    port map (
            O => \N__6987\,
            I => \N__6980\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__6980\,
            I => \U712_REG_SM.N_174\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__6977\,
            I => \N__6974\
        );

    \I__1435\ : InMux
    port map (
            O => \N__6974\,
            I => \N__6970\
        );

    \I__1434\ : InMux
    port map (
            O => \N__6973\,
            I => \N__6967\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__6970\,
            I => \REG_TACK\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__6967\,
            I => \REG_TACK\
        );

    \I__1431\ : InMux
    port map (
            O => \N__6962\,
            I => \N__6958\
        );

    \I__1430\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6955\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__6958\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__6955\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__1427\ : IoInMux
    port map (
            O => \N__6950\,
            I => \N__6947\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__6947\,
            I => \N__6944\
        );

    \I__1425\ : Span12Mux_s1_v
    port map (
            O => \N__6944\,
            I => \N__6941\
        );

    \I__1424\ : Span12Mux_h
    port map (
            O => \N__6941\,
            I => \N__6938\
        );

    \I__1423\ : Odrv12
    port map (
            O => \N__6938\,
            I => \CASn_c\
        );

    \I__1422\ : IoInMux
    port map (
            O => \N__6935\,
            I => \N__6932\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__6932\,
            I => \N__6929\
        );

    \I__1420\ : Span4Mux_s3_v
    port map (
            O => \N__6929\,
            I => \N__6926\
        );

    \I__1419\ : Span4Mux_v
    port map (
            O => \N__6926\,
            I => \N__6923\
        );

    \I__1418\ : Span4Mux_h
    port map (
            O => \N__6923\,
            I => \N__6920\
        );

    \I__1417\ : Span4Mux_h
    port map (
            O => \N__6920\,
            I => \N__6917\
        );

    \I__1416\ : Odrv4
    port map (
            O => \N__6917\,
            I => \CMA_c_10\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6914\,
            I => \N__6911\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__6911\,
            I => \N__6908\
        );

    \I__1413\ : Odrv12
    port map (
            O => \N__6908\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__6905\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\
        );

    \I__1411\ : IoInMux
    port map (
            O => \N__6902\,
            I => \N__6899\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__6899\,
            I => \N__6896\
        );

    \I__1409\ : IoSpan4Mux
    port map (
            O => \N__6896\,
            I => \N__6893\
        );

    \I__1408\ : Span4Mux_s3_v
    port map (
            O => \N__6893\,
            I => \N__6890\
        );

    \I__1407\ : Span4Mux_v
    port map (
            O => \N__6890\,
            I => \N__6887\
        );

    \I__1406\ : Odrv4
    port map (
            O => \N__6887\,
            I => \CMA_c_2\
        );

    \I__1405\ : CascadeMux
    port map (
            O => \N__6884\,
            I => \N__6878\
        );

    \I__1404\ : CascadeMux
    port map (
            O => \N__6883\,
            I => \N__6873\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__6882\,
            I => \N__6868\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6863\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6878\,
            I => \N__6863\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__6877\,
            I => \N__6860\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6876\,
            I => \N__6856\
        );

    \I__1398\ : InMux
    port map (
            O => \N__6873\,
            I => \N__6851\
        );

    \I__1397\ : InMux
    port map (
            O => \N__6872\,
            I => \N__6851\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6871\,
            I => \N__6848\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6868\,
            I => \N__6845\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6863\,
            I => \N__6842\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6860\,
            I => \N__6837\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6859\,
            I => \N__6837\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6856\,
            I => \N__6834\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6851\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__6848\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__6845\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__6842\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__6837\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1385\ : Odrv4
    port map (
            O => \N__6834\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6821\,
            I => \N__6818\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__6818\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1382\ : IoInMux
    port map (
            O => \N__6815\,
            I => \N__6812\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__6812\,
            I => \N__6809\
        );

    \I__1380\ : IoSpan4Mux
    port map (
            O => \N__6809\,
            I => \N__6806\
        );

    \I__1379\ : IoSpan4Mux
    port map (
            O => \N__6806\,
            I => \N__6803\
        );

    \I__1378\ : Span4Mux_s2_h
    port map (
            O => \N__6803\,
            I => \N__6800\
        );

    \I__1377\ : Sp12to4
    port map (
            O => \N__6800\,
            I => \N__6797\
        );

    \I__1376\ : Span12Mux_h
    port map (
            O => \N__6797\,
            I => \N__6794\
        );

    \I__1375\ : Odrv12
    port map (
            O => \N__6794\,
            I => \CMA_c_3\
        );

    \I__1374\ : CascadeMux
    port map (
            O => \N__6791\,
            I => \U712_REG_SM.N_199_cascade_\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__6788\,
            I => \N__6784\
        );

    \I__1372\ : InMux
    port map (
            O => \N__6787\,
            I => \N__6781\
        );

    \I__1371\ : InMux
    port map (
            O => \N__6784\,
            I => \N__6778\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__6781\,
            I => \N__6775\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__6778\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1368\ : Odrv12
    port map (
            O => \N__6775\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__6770\,
            I => \N__6767\
        );

    \I__1366\ : InMux
    port map (
            O => \N__6767\,
            I => \N__6762\
        );

    \I__1365\ : InMux
    port map (
            O => \N__6766\,
            I => \N__6759\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6756\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__6762\,
            I => \N__6753\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__6759\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6756\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1360\ : Odrv12
    port map (
            O => \N__6753\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__6746\,
            I => \U712_CYCLE_TERM.N_208_i_0_en_cascade_\
        );

    \I__1358\ : CEMux
    port map (
            O => \N__6743\,
            I => \N__6740\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__6740\,
            I => \N__6737\
        );

    \I__1356\ : Odrv12
    port map (
            O => \N__6737\,
            I => \U712_CYCLE_TERM.N_208_i_0_en_0\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6734\,
            I => \N__6731\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6731\,
            I => \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a3_0_2\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__6728\,
            I => \N__6724\
        );

    \I__1352\ : InMux
    port map (
            O => \N__6727\,
            I => \N__6721\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6715\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6721\,
            I => \N__6711\
        );

    \I__1349\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6708\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6702\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6718\,
            I => \N__6702\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__6715\,
            I => \N__6698\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6714\,
            I => \N__6688\
        );

    \I__1344\ : Span4Mux_v
    port map (
            O => \N__6711\,
            I => \N__6685\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__6708\,
            I => \N__6682\
        );

    \I__1342\ : InMux
    port map (
            O => \N__6707\,
            I => \N__6679\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__6702\,
            I => \N__6676\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6701\,
            I => \N__6673\
        );

    \I__1339\ : Span4Mux_v
    port map (
            O => \N__6698\,
            I => \N__6670\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6697\,
            I => \N__6667\
        );

    \I__1337\ : InMux
    port map (
            O => \N__6696\,
            I => \N__6662\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6695\,
            I => \N__6662\
        );

    \I__1335\ : InMux
    port map (
            O => \N__6694\,
            I => \N__6657\
        );

    \I__1334\ : InMux
    port map (
            O => \N__6693\,
            I => \N__6657\
        );

    \I__1333\ : InMux
    port map (
            O => \N__6692\,
            I => \N__6652\
        );

    \I__1332\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6652\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__6688\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__6685\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__6682\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__6679\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__6676\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__6673\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1325\ : Odrv4
    port map (
            O => \N__6670\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6667\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__6662\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6657\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6652\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6624\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__6628\,
            I => \N__6620\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__6627\,
            I => \N__6617\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6624\,
            I => \N__6607\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6623\,
            I => \N__6604\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6620\,
            I => \N__6599\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6617\,
            I => \N__6599\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6616\,
            I => \N__6596\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6615\,
            I => \N__6593\
        );

    \I__1311\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6588\
        );

    \I__1310\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6588\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6612\,
            I => \N__6585\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6611\,
            I => \N__6580\
        );

    \I__1307\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6580\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__6607\,
            I => \U712_CHIP_RAM.N_165\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6604\,
            I => \U712_CHIP_RAM.N_165\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__6599\,
            I => \U712_CHIP_RAM.N_165\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6596\,
            I => \U712_CHIP_RAM.N_165\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__6593\,
            I => \U712_CHIP_RAM.N_165\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__6588\,
            I => \U712_CHIP_RAM.N_165\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6585\,
            I => \U712_CHIP_RAM.N_165\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6580\,
            I => \U712_CHIP_RAM.N_165\
        );

    \I__1298\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6560\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6560\,
            I => \U712_CHIP_RAM.N_249\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6557\,
            I => \N__6553\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6550\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6553\,
            I => \N__6547\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6550\,
            I => \CPU_TACKm\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__6547\,
            I => \CPU_TACKm\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__6542\,
            I => \N__6537\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6541\,
            I => \N__6534\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6540\,
            I => \N__6529\
        );

    \I__1288\ : InMux
    port map (
            O => \N__6537\,
            I => \N__6529\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__6534\,
            I => \N__6523\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__6529\,
            I => \N__6523\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6528\,
            I => \N__6520\
        );

    \I__1284\ : Odrv12
    port map (
            O => \N__6523\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6520\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__6515\,
            I => \N__6512\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6512\,
            I => \N__6509\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__6509\,
            I => \N__6506\
        );

    \I__1279\ : Odrv4
    port map (
            O => \N__6506\,
            I => \U712_REG_SM.N_199\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6500\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6500\,
            I => \U712_REG_SM.N_171\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__6497\,
            I => \U712_REG_SM.N_174_cascade_\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6494\,
            I => \N__6490\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6493\,
            I => \N__6487\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__6490\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6487\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1271\ : InMux
    port map (
            O => \N__6482\,
            I => \N__6478\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6481\,
            I => \N__6475\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__6478\,
            I => \N__6472\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6475\,
            I => \N__6469\
        );

    \I__1267\ : Sp12to4
    port map (
            O => \N__6472\,
            I => \N__6466\
        );

    \I__1266\ : Span4Mux_v
    port map (
            O => \N__6469\,
            I => \N__6463\
        );

    \I__1265\ : Span12Mux_h
    port map (
            O => \N__6466\,
            I => \N__6460\
        );

    \I__1264\ : Sp12to4
    port map (
            O => \N__6463\,
            I => \N__6457\
        );

    \I__1263\ : Span12Mux_v
    port map (
            O => \N__6460\,
            I => \N__6452\
        );

    \I__1262\ : Span12Mux_h
    port map (
            O => \N__6457\,
            I => \N__6452\
        );

    \I__1261\ : Odrv12
    port map (
            O => \N__6452\,
            I => \RnW_c\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6449\,
            I => \N__6446\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6446\,
            I => \N__6441\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6445\,
            I => \N__6438\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6444\,
            I => \N__6435\
        );

    \I__1256\ : Span4Mux_h
    port map (
            O => \N__6441\,
            I => \N__6430\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__6438\,
            I => \N__6430\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6435\,
            I => \N__6427\
        );

    \I__1253\ : Span4Mux_h
    port map (
            O => \N__6430\,
            I => \N__6424\
        );

    \I__1252\ : Span4Mux_v
    port map (
            O => \N__6427\,
            I => \N__6421\
        );

    \I__1251\ : Sp12to4
    port map (
            O => \N__6424\,
            I => \N__6418\
        );

    \I__1250\ : IoSpan4Mux
    port map (
            O => \N__6421\,
            I => \N__6415\
        );

    \I__1249\ : Span12Mux_v
    port map (
            O => \N__6418\,
            I => \N__6412\
        );

    \I__1248\ : IoSpan4Mux
    port map (
            O => \N__6415\,
            I => \N__6409\
        );

    \I__1247\ : Odrv12
    port map (
            O => \N__6412\,
            I => \AWEn_c\
        );

    \I__1246\ : Odrv4
    port map (
            O => \N__6409\,
            I => \AWEn_c\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6404\,
            I => \N__6398\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6403\,
            I => \N__6391\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6402\,
            I => \N__6391\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6401\,
            I => \N__6388\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6398\,
            I => \N__6385\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6382\
        );

    \I__1239\ : CascadeMux
    port map (
            O => \N__6396\,
            I => \N__6377\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6391\,
            I => \N__6372\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6388\,
            I => \N__6369\
        );

    \I__1236\ : Span4Mux_h
    port map (
            O => \N__6385\,
            I => \N__6366\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6382\,
            I => \N__6363\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6381\,
            I => \N__6358\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6380\,
            I => \N__6358\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6377\,
            I => \N__6353\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6376\,
            I => \N__6353\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6375\,
            I => \N__6350\
        );

    \I__1229\ : Span4Mux_h
    port map (
            O => \N__6372\,
            I => \N__6347\
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__6369\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1227\ : Odrv4
    port map (
            O => \N__6366\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1226\ : Odrv4
    port map (
            O => \N__6363\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6358\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6353\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6350\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__6347\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6332\,
            I => \N__6329\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6329\,
            I => \N__6326\
        );

    \I__1219\ : Odrv4
    port map (
            O => \N__6326\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_RNOZ0Z_0\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__6323\,
            I => \N__6317\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__6322\,
            I => \N__6313\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6321\,
            I => \N__6309\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6320\,
            I => \N__6306\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6317\,
            I => \N__6302\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6299\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6290\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6290\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6309\,
            I => \N__6285\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6306\,
            I => \N__6285\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6282\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6302\,
            I => \N__6277\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__6299\,
            I => \N__6277\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__6298\,
            I => \N__6274\
        );

    \I__1204\ : CascadeMux
    port map (
            O => \N__6297\,
            I => \N__6270\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6296\,
            I => \N__6262\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6295\,
            I => \N__6259\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6290\,
            I => \N__6256\
        );

    \I__1200\ : Span4Mux_h
    port map (
            O => \N__6285\,
            I => \N__6251\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6282\,
            I => \N__6251\
        );

    \I__1198\ : Span4Mux_v
    port map (
            O => \N__6277\,
            I => \N__6248\
        );

    \I__1197\ : InMux
    port map (
            O => \N__6274\,
            I => \N__6245\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6273\,
            I => \N__6242\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6239\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6234\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6234\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6227\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6266\,
            I => \N__6227\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6265\,
            I => \N__6227\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__6262\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6259\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__6256\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1186\ : Odrv4
    port map (
            O => \N__6251\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1185\ : Odrv4
    port map (
            O => \N__6248\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6245\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6242\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6239\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6234\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6227\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6206\,
            I => \N__6203\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6203\,
            I => \N__6199\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6196\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__6199\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6196\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__6191\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1_cascade_\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6188\,
            I => \N__6182\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__6187\,
            I => \N__6178\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6186\,
            I => \N__6172\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6168\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6182\,
            I => \N__6165\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6162\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6178\,
            I => \N__6158\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6177\,
            I => \N__6152\
        );

    \I__1165\ : InMux
    port map (
            O => \N__6176\,
            I => \N__6152\
        );

    \I__1164\ : InMux
    port map (
            O => \N__6175\,
            I => \N__6148\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6172\,
            I => \N__6145\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6142\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__6168\,
            I => \N__6137\
        );

    \I__1160\ : Span4Mux_v
    port map (
            O => \N__6165\,
            I => \N__6137\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6162\,
            I => \N__6134\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6131\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6158\,
            I => \N__6128\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6125\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6152\,
            I => \N__6122\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6151\,
            I => \N__6119\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6148\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__6145\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__6142\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1150\ : Odrv4
    port map (
            O => \N__6137\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__6134\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6131\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1147\ : Odrv12
    port map (
            O => \N__6128\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6125\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__6122\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6119\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6098\,
            I => \N__6095\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__6095\,
            I => \N__6092\
        );

    \I__1141\ : Odrv4
    port map (
            O => \N__6092\,
            I => \U712_CHIP_RAM.N_248\
        );

    \I__1140\ : CascadeMux
    port map (
            O => \N__6089\,
            I => \N__6085\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__6088\,
            I => \N__6081\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6074\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6084\,
            I => \N__6071\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6068\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6080\,
            I => \N__6065\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6079\,
            I => \N__6062\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6057\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6050\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6074\,
            I => \N__6045\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__6071\,
            I => \N__6045\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6068\,
            I => \N__6038\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6065\,
            I => \N__6033\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__6062\,
            I => \N__6033\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6061\,
            I => \N__6030\
        );

    \I__1125\ : InMux
    port map (
            O => \N__6060\,
            I => \N__6027\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6057\,
            I => \N__6024\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6056\,
            I => \N__6021\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6055\,
            I => \N__6016\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6054\,
            I => \N__6016\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6053\,
            I => \N__6013\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6050\,
            I => \N__6008\
        );

    \I__1118\ : Span4Mux_v
    port map (
            O => \N__6045\,
            I => \N__6008\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6044\,
            I => \N__6003\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6043\,
            I => \N__6003\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6042\,
            I => \N__5998\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6041\,
            I => \N__5998\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__6038\,
            I => \N__5993\
        );

    \I__1112\ : Span4Mux_v
    port map (
            O => \N__6033\,
            I => \N__5993\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__6030\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6027\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__6024\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6021\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6016\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6013\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1105\ : Odrv4
    port map (
            O => \N__6008\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6003\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5998\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__5993\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5968\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5965\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5968\,
            I => \N__5958\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5965\,
            I => \N__5958\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5964\,
            I => \N__5955\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5963\,
            I => \N__5952\
        );

    \I__1095\ : Span4Mux_h
    port map (
            O => \N__5958\,
            I => \N__5949\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__5955\,
            I => \N__5946\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5952\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2Z0Z_1\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__5949\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2Z0Z_1\
        );

    \I__1091\ : Odrv4
    port map (
            O => \N__5946\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2Z0Z_1\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__5939\,
            I => \U712_REG_SM.N_171_cascade_\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__5936\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa_0_a2_0_a3_1_cascade_\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__5933\,
            I => \N__5929\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5932\,
            I => \N__5926\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5929\,
            I => \N__5923\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5926\,
            I => \N__5920\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__5923\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__1083\ : Odrv4
    port map (
            O => \N__5920\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__5915\,
            I => \N__5912\
        );

    \I__1081\ : InMux
    port map (
            O => \N__5912\,
            I => \N__5906\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5906\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__5906\,
            I => \N__5903\
        );

    \I__1078\ : Span4Mux_v
    port map (
            O => \N__5903\,
            I => \N__5900\
        );

    \I__1077\ : Span4Mux_v
    port map (
            O => \N__5900\,
            I => \N__5897\
        );

    \I__1076\ : Sp12to4
    port map (
            O => \N__5897\,
            I => \N__5894\
        );

    \I__1075\ : Span12Mux_h
    port map (
            O => \N__5894\,
            I => \N__5891\
        );

    \I__1074\ : Odrv12
    port map (
            O => \N__5891\,
            I => \A_c_14\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5885\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5885\,
            I => \N__5882\
        );

    \I__1071\ : Span4Mux_v
    port map (
            O => \N__5882\,
            I => \N__5879\
        );

    \I__1070\ : Sp12to4
    port map (
            O => \N__5879\,
            I => \N__5876\
        );

    \I__1069\ : Span12Mux_h
    port map (
            O => \N__5876\,
            I => \N__5873\
        );

    \I__1068\ : Span12Mux_v
    port map (
            O => \N__5873\,
            I => \N__5870\
        );

    \I__1067\ : Odrv12
    port map (
            O => \N__5870\,
            I => \A_c_3\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5864\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5864\,
            I => \N__5861\
        );

    \I__1064\ : Span4Mux_v
    port map (
            O => \N__5861\,
            I => \N__5858\
        );

    \I__1063\ : Sp12to4
    port map (
            O => \N__5858\,
            I => \N__5855\
        );

    \I__1062\ : Span12Mux_h
    port map (
            O => \N__5855\,
            I => \N__5852\
        );

    \I__1061\ : Odrv12
    port map (
            O => \N__5852\,
            I => \A_c_10\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__5849\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\
        );

    \I__1059\ : InMux
    port map (
            O => \N__5846\,
            I => \N__5843\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__5843\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__5840\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5834\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__5834\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1054\ : IoInMux
    port map (
            O => \N__5831\,
            I => \N__5828\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__5828\,
            I => \N__5825\
        );

    \I__1052\ : Span4Mux_s3_v
    port map (
            O => \N__5825\,
            I => \N__5822\
        );

    \I__1051\ : Span4Mux_v
    port map (
            O => \N__5822\,
            I => \N__5819\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__5819\,
            I => \N__5816\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__5816\,
            I => \CMA_c_1\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5813\,
            I => \N__5810\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5810\,
            I => \N__5807\
        );

    \I__1046\ : Odrv4
    port map (
            O => \N__5807\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1045\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5801\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__5801\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1043\ : IoInMux
    port map (
            O => \N__5798\,
            I => \N__5795\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5795\,
            I => \N__5792\
        );

    \I__1041\ : Span4Mux_s1_h
    port map (
            O => \N__5792\,
            I => \N__5789\
        );

    \I__1040\ : Span4Mux_h
    port map (
            O => \N__5789\,
            I => \N__5786\
        );

    \I__1039\ : Sp12to4
    port map (
            O => \N__5786\,
            I => \N__5783\
        );

    \I__1038\ : Span12Mux_s8_v
    port map (
            O => \N__5783\,
            I => \N__5780\
        );

    \I__1037\ : Span12Mux_h
    port map (
            O => \N__5780\,
            I => \N__5777\
        );

    \I__1036\ : Odrv12
    port map (
            O => \N__5777\,
            I => \CMA_c_5\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5774\,
            I => \N__5771\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5771\,
            I => \N__5768\
        );

    \I__1033\ : Span4Mux_v
    port map (
            O => \N__5768\,
            I => \N__5765\
        );

    \I__1032\ : Span4Mux_h
    port map (
            O => \N__5765\,
            I => \N__5762\
        );

    \I__1031\ : Sp12to4
    port map (
            O => \N__5762\,
            I => \N__5759\
        );

    \I__1030\ : Odrv12
    port map (
            O => \N__5759\,
            I => \A_c_7\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__5756\,
            I => \U712_CHIP_RAM.N_324_cascade_\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5753\,
            I => \N__5750\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5750\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5747\,
            I => \N__5744\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5744\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1024\ : IoInMux
    port map (
            O => \N__5741\,
            I => \N__5738\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__5738\,
            I => \N__5735\
        );

    \I__1022\ : IoSpan4Mux
    port map (
            O => \N__5735\,
            I => \N__5732\
        );

    \I__1021\ : Span4Mux_s3_h
    port map (
            O => \N__5732\,
            I => \N__5729\
        );

    \I__1020\ : Sp12to4
    port map (
            O => \N__5729\,
            I => \N__5726\
        );

    \I__1019\ : Span12Mux_h
    port map (
            O => \N__5726\,
            I => \N__5723\
        );

    \I__1018\ : Odrv12
    port map (
            O => \N__5723\,
            I => \CMA_c_7\
        );

    \I__1017\ : InMux
    port map (
            O => \N__5720\,
            I => \N__5717\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5717\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1015\ : IoInMux
    port map (
            O => \N__5714\,
            I => \N__5711\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5711\,
            I => \N__5708\
        );

    \I__1013\ : Span4Mux_s2_h
    port map (
            O => \N__5708\,
            I => \N__5705\
        );

    \I__1012\ : Span4Mux_v
    port map (
            O => \N__5705\,
            I => \N__5702\
        );

    \I__1011\ : Span4Mux_v
    port map (
            O => \N__5702\,
            I => \N__5699\
        );

    \I__1010\ : Sp12to4
    port map (
            O => \N__5699\,
            I => \N__5696\
        );

    \I__1009\ : Span12Mux_s9_h
    port map (
            O => \N__5696\,
            I => \N__5693\
        );

    \I__1008\ : Odrv12
    port map (
            O => \N__5693\,
            I => \CMA_c_6\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5690\,
            I => \N__5687\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__5687\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__5684\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_\
        );

    \I__1004\ : IoInMux
    port map (
            O => \N__5681\,
            I => \N__5678\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5678\,
            I => \N__5675\
        );

    \I__1002\ : IoSpan4Mux
    port map (
            O => \N__5675\,
            I => \N__5672\
        );

    \I__1001\ : Span4Mux_s1_h
    port map (
            O => \N__5672\,
            I => \N__5669\
        );

    \I__1000\ : Sp12to4
    port map (
            O => \N__5669\,
            I => \N__5666\
        );

    \I__999\ : Span12Mux_s11_v
    port map (
            O => \N__5666\,
            I => \N__5663\
        );

    \I__998\ : Span12Mux_h
    port map (
            O => \N__5663\,
            I => \N__5660\
        );

    \I__997\ : Odrv12
    port map (
            O => \N__5660\,
            I => \CMA_c_4\
        );

    \I__996\ : CascadeMux
    port map (
            O => \N__5657\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\
        );

    \I__995\ : InMux
    port map (
            O => \N__5654\,
            I => \N__5651\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5651\,
            I => \N__5648\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__5648\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__992\ : IoInMux
    port map (
            O => \N__5645\,
            I => \N__5642\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5642\,
            I => \N__5639\
        );

    \I__990\ : IoSpan4Mux
    port map (
            O => \N__5639\,
            I => \N__5636\
        );

    \I__989\ : Span4Mux_s2_v
    port map (
            O => \N__5636\,
            I => \N__5631\
        );

    \I__988\ : InMux
    port map (
            O => \N__5635\,
            I => \N__5626\
        );

    \I__987\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5626\
        );

    \I__986\ : Sp12to4
    port map (
            O => \N__5631\,
            I => \N__5623\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__5626\,
            I => \N__5620\
        );

    \I__984\ : Span12Mux_v
    port map (
            O => \N__5623\,
            I => \N__5616\
        );

    \I__983\ : Span4Mux_v
    port map (
            O => \N__5620\,
            I => \N__5613\
        );

    \I__982\ : InMux
    port map (
            O => \N__5619\,
            I => \N__5610\
        );

    \I__981\ : Odrv12
    port map (
            O => \N__5616\,
            I => \DBENn_c\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__5613\,
            I => \DBENn_c\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__5610\,
            I => \DBENn_c\
        );

    \I__978\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5600\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5600\,
            I => \U712_BYTE_ENABLE.N_268\
        );

    \I__976\ : IoInMux
    port map (
            O => \N__5597\,
            I => \N__5594\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__5594\,
            I => \N__5591\
        );

    \I__974\ : IoSpan4Mux
    port map (
            O => \N__5591\,
            I => \N__5588\
        );

    \I__973\ : IoSpan4Mux
    port map (
            O => \N__5588\,
            I => \N__5585\
        );

    \I__972\ : Sp12to4
    port map (
            O => \N__5585\,
            I => \N__5582\
        );

    \I__971\ : Span12Mux_s7_v
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__970\ : Span12Mux_h
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__969\ : Odrv12
    port map (
            O => \N__5576\,
            I => \N_185_i\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__5573\,
            I => \U712_BYTE_ENABLE.N_270_cascade_\
        );

    \I__967\ : IoInMux
    port map (
            O => \N__5570\,
            I => \N__5567\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5567\,
            I => \N__5564\
        );

    \I__965\ : IoSpan4Mux
    port map (
            O => \N__5564\,
            I => \N__5561\
        );

    \I__964\ : Sp12to4
    port map (
            O => \N__5561\,
            I => \N__5558\
        );

    \I__963\ : Span12Mux_s7_v
    port map (
            O => \N__5558\,
            I => \N__5555\
        );

    \I__962\ : Span12Mux_h
    port map (
            O => \N__5555\,
            I => \N__5552\
        );

    \I__961\ : Span12Mux_v
    port map (
            O => \N__5552\,
            I => \N__5549\
        );

    \I__960\ : Odrv12
    port map (
            O => \N__5549\,
            I => \N_186_i\
        );

    \I__959\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5543\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__5543\,
            I => \U712_BYTE_ENABLE.N_272\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__5540\,
            I => \N__5536\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__5539\,
            I => \N__5533\
        );

    \I__955\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5530\
        );

    \I__954\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5527\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5530\,
            I => \N__5523\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__5527\,
            I => \N__5520\
        );

    \I__951\ : InMux
    port map (
            O => \N__5526\,
            I => \N__5517\
        );

    \I__950\ : Span4Mux_v
    port map (
            O => \N__5523\,
            I => \N__5512\
        );

    \I__949\ : Span4Mux_v
    port map (
            O => \N__5520\,
            I => \N__5512\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5517\,
            I => \N__5509\
        );

    \I__947\ : Sp12to4
    port map (
            O => \N__5512\,
            I => \N__5506\
        );

    \I__946\ : Span12Mux_h
    port map (
            O => \N__5509\,
            I => \N__5503\
        );

    \I__945\ : Span12Mux_h
    port map (
            O => \N__5506\,
            I => \N__5500\
        );

    \I__944\ : Span12Mux_v
    port map (
            O => \N__5503\,
            I => \N__5497\
        );

    \I__943\ : Span12Mux_v
    port map (
            O => \N__5500\,
            I => \N__5494\
        );

    \I__942\ : Odrv12
    port map (
            O => \N__5497\,
            I => \CASLn_c\
        );

    \I__941\ : Odrv12
    port map (
            O => \N__5494\,
            I => \CASLn_c\
        );

    \I__940\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5483\
        );

    \I__939\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5483\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5483\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0\
        );

    \I__937\ : IoInMux
    port map (
            O => \N__5480\,
            I => \N__5477\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5477\,
            I => \N__5474\
        );

    \I__935\ : IoSpan4Mux
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__934\ : Sp12to4
    port map (
            O => \N__5471\,
            I => \N__5468\
        );

    \I__933\ : Span12Mux_s7_v
    port map (
            O => \N__5468\,
            I => \N__5465\
        );

    \I__932\ : Span12Mux_v
    port map (
            O => \N__5465\,
            I => \N__5462\
        );

    \I__931\ : Odrv12
    port map (
            O => \N__5462\,
            I => \N_187_i\
        );

    \I__930\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5453\
        );

    \I__929\ : InMux
    port map (
            O => \N__5458\,
            I => \N__5453\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5453\,
            I => \N__5448\
        );

    \I__927\ : InMux
    port map (
            O => \N__5452\,
            I => \N__5443\
        );

    \I__926\ : InMux
    port map (
            O => \N__5451\,
            I => \N__5443\
        );

    \I__925\ : Span4Mux_v
    port map (
            O => \N__5448\,
            I => \N__5440\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5443\,
            I => \N__5437\
        );

    \I__923\ : Span4Mux_v
    port map (
            O => \N__5440\,
            I => \N__5434\
        );

    \I__922\ : Span4Mux_v
    port map (
            O => \N__5437\,
            I => \N__5431\
        );

    \I__921\ : Span4Mux_h
    port map (
            O => \N__5434\,
            I => \N__5428\
        );

    \I__920\ : Span4Mux_v
    port map (
            O => \N__5431\,
            I => \N__5425\
        );

    \I__919\ : Sp12to4
    port map (
            O => \N__5428\,
            I => \N__5420\
        );

    \I__918\ : Sp12to4
    port map (
            O => \N__5425\,
            I => \N__5420\
        );

    \I__917\ : Odrv12
    port map (
            O => \N__5420\,
            I => \A_c_1\
        );

    \I__916\ : InMux
    port map (
            O => \N__5417\,
            I => \N__5405\
        );

    \I__915\ : InMux
    port map (
            O => \N__5416\,
            I => \N__5405\
        );

    \I__914\ : InMux
    port map (
            O => \N__5415\,
            I => \N__5405\
        );

    \I__913\ : InMux
    port map (
            O => \N__5414\,
            I => \N__5405\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__5405\,
            I => \U712_BYTE_ENABLE.N_265\
        );

    \I__911\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5396\
        );

    \I__910\ : InMux
    port map (
            O => \N__5401\,
            I => \N__5396\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5396\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0\
        );

    \I__908\ : CascadeMux
    port map (
            O => \N__5393\,
            I => \U712_BYTE_ENABLE.N_266_cascade_\
        );

    \I__907\ : InMux
    port map (
            O => \N__5390\,
            I => \N__5385\
        );

    \I__906\ : InMux
    port map (
            O => \N__5389\,
            I => \N__5380\
        );

    \I__905\ : InMux
    port map (
            O => \N__5388\,
            I => \N__5380\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5385\,
            I => \N__5375\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5380\,
            I => \N__5375\
        );

    \I__902\ : Span12Mux_v
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__901\ : Span12Mux_h
    port map (
            O => \N__5372\,
            I => \N__5369\
        );

    \I__900\ : Odrv12
    port map (
            O => \N__5369\,
            I => \CASUn_c\
        );

    \I__899\ : IoInMux
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__5363\,
            I => \N__5360\
        );

    \I__897\ : Span4Mux_s2_h
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__896\ : Span4Mux_h
    port map (
            O => \N__5357\,
            I => \N__5354\
        );

    \I__895\ : Sp12to4
    port map (
            O => \N__5354\,
            I => \N__5351\
        );

    \I__894\ : Span12Mux_v
    port map (
            O => \N__5351\,
            I => \N__5348\
        );

    \I__893\ : Span12Mux_h
    port map (
            O => \N__5348\,
            I => \N__5345\
        );

    \I__892\ : Odrv12
    port map (
            O => \N__5345\,
            I => \N_184_i\
        );

    \I__891\ : InMux
    port map (
            O => \N__5342\,
            I => \N__5339\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5339\,
            I => \N__5336\
        );

    \I__889\ : Span4Mux_v
    port map (
            O => \N__5336\,
            I => \N__5331\
        );

    \I__888\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5326\
        );

    \I__887\ : InMux
    port map (
            O => \N__5334\,
            I => \N__5326\
        );

    \I__886\ : Span4Mux_v
    port map (
            O => \N__5331\,
            I => \N__5320\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5326\,
            I => \N__5320\
        );

    \I__884\ : InMux
    port map (
            O => \N__5325\,
            I => \N__5317\
        );

    \I__883\ : Span4Mux_v
    port map (
            O => \N__5320\,
            I => \N__5312\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__5317\,
            I => \N__5309\
        );

    \I__881\ : InMux
    port map (
            O => \N__5316\,
            I => \N__5304\
        );

    \I__880\ : InMux
    port map (
            O => \N__5315\,
            I => \N__5304\
        );

    \I__879\ : Odrv4
    port map (
            O => \N__5312\,
            I => \DMA_CYCLEm\
        );

    \I__878\ : Odrv12
    port map (
            O => \N__5309\,
            I => \DMA_CYCLEm\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5304\,
            I => \DMA_CYCLEm\
        );

    \I__876\ : IoInMux
    port map (
            O => \N__5297\,
            I => \N__5294\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5294\,
            I => \N__5291\
        );

    \I__874\ : Span4Mux_s1_h
    port map (
            O => \N__5291\,
            I => \N__5288\
        );

    \I__873\ : Sp12to4
    port map (
            O => \N__5288\,
            I => \N__5285\
        );

    \I__872\ : Span12Mux_s6_v
    port map (
            O => \N__5285\,
            I => \N__5282\
        );

    \I__871\ : Span12Mux_h
    port map (
            O => \N__5282\,
            I => \N__5279\
        );

    \I__870\ : Odrv12
    port map (
            O => \N__5279\,
            I => \DRDDIR_i_m2\
        );

    \I__869\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5273\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5273\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__867\ : IoInMux
    port map (
            O => \N__5270\,
            I => \N__5267\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5267\,
            I => \N__5264\
        );

    \I__865\ : Span4Mux_s2_v
    port map (
            O => \N__5264\,
            I => \N__5261\
        );

    \I__864\ : Span4Mux_v
    port map (
            O => \N__5261\,
            I => \N__5258\
        );

    \I__863\ : Span4Mux_v
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__862\ : Span4Mux_h
    port map (
            O => \N__5255\,
            I => \N__5252\
        );

    \I__861\ : Odrv4
    port map (
            O => \N__5252\,
            I => \CMA_c_0\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__5249\,
            I => \U712_CHIP_RAM.N_219_cascade_\
        );

    \I__859\ : InMux
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5243\,
            I => \N__5236\
        );

    \I__857\ : InMux
    port map (
            O => \N__5242\,
            I => \N__5233\
        );

    \I__856\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5230\
        );

    \I__855\ : InMux
    port map (
            O => \N__5240\,
            I => \N__5227\
        );

    \I__854\ : InMux
    port map (
            O => \N__5239\,
            I => \N__5224\
        );

    \I__853\ : Span4Mux_v
    port map (
            O => \N__5236\,
            I => \N__5217\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5233\,
            I => \N__5217\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5230\,
            I => \N__5217\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5227\,
            I => \N__5214\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5224\,
            I => \U712_CHIP_RAM.N_166\
        );

    \I__848\ : Odrv4
    port map (
            O => \N__5217\,
            I => \U712_CHIP_RAM.N_166\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__5214\,
            I => \U712_CHIP_RAM.N_166\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__5207\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_7_i_2_cascade_\
        );

    \I__845\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5201\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5201\,
            I => \N__5198\
        );

    \I__843\ : Odrv12
    port map (
            O => \N__5198\,
            I => \U712_CHIP_RAM.N_258\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__5195\,
            I => \U712_CHIP_RAM.N_49_cascade_\
        );

    \I__841\ : InMux
    port map (
            O => \N__5192\,
            I => \N__5188\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__5191\,
            I => \N__5184\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5188\,
            I => \N__5181\
        );

    \I__838\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5178\
        );

    \I__837\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5175\
        );

    \I__836\ : Span4Mux_v
    port map (
            O => \N__5181\,
            I => \N__5172\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__5178\,
            I => \U712_CHIP_RAM.N_206\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5175\,
            I => \U712_CHIP_RAM.N_206\
        );

    \I__833\ : Odrv4
    port map (
            O => \N__5172\,
            I => \U712_CHIP_RAM.N_206\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__5165\,
            I => \N__5162\
        );

    \I__831\ : InMux
    port map (
            O => \N__5162\,
            I => \N__5159\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5159\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_1\
        );

    \I__829\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5150\
        );

    \I__828\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5147\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__5154\,
            I => \N__5144\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__5153\,
            I => \N__5134\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5150\,
            I => \N__5128\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5147\,
            I => \N__5128\
        );

    \I__823\ : InMux
    port map (
            O => \N__5144\,
            I => \N__5123\
        );

    \I__822\ : InMux
    port map (
            O => \N__5143\,
            I => \N__5123\
        );

    \I__821\ : InMux
    port map (
            O => \N__5142\,
            I => \N__5119\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__5141\,
            I => \N__5114\
        );

    \I__819\ : InMux
    port map (
            O => \N__5140\,
            I => \N__5110\
        );

    \I__818\ : InMux
    port map (
            O => \N__5139\,
            I => \N__5105\
        );

    \I__817\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5105\
        );

    \I__816\ : InMux
    port map (
            O => \N__5137\,
            I => \N__5102\
        );

    \I__815\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5097\
        );

    \I__814\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5097\
        );

    \I__813\ : Span4Mux_h
    port map (
            O => \N__5128\,
            I => \N__5092\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5123\,
            I => \N__5092\
        );

    \I__811\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5089\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__5119\,
            I => \N__5086\
        );

    \I__809\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5081\
        );

    \I__808\ : InMux
    port map (
            O => \N__5117\,
            I => \N__5081\
        );

    \I__807\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5076\
        );

    \I__806\ : InMux
    port map (
            O => \N__5113\,
            I => \N__5076\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5110\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5105\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5102\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5097\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__801\ : Odrv4
    port map (
            O => \N__5092\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__5089\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__799\ : Odrv4
    port map (
            O => \N__5086\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5081\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5076\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__796\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5053\
        );

    \I__795\ : InMux
    port map (
            O => \N__5056\,
            I => \N__5050\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__5053\,
            I => \N__5047\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5050\,
            I => \N__5038\
        );

    \I__792\ : Span4Mux_h
    port map (
            O => \N__5047\,
            I => \N__5038\
        );

    \I__791\ : InMux
    port map (
            O => \N__5046\,
            I => \N__5031\
        );

    \I__790\ : InMux
    port map (
            O => \N__5045\,
            I => \N__5031\
        );

    \I__789\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5031\
        );

    \I__788\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5028\
        );

    \I__787\ : Odrv4
    port map (
            O => \N__5038\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5031\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5028\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__784\ : InMux
    port map (
            O => \N__5021\,
            I => \N__5017\
        );

    \I__783\ : InMux
    port map (
            O => \N__5020\,
            I => \N__5014\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5017\,
            I => \N__5011\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5014\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__780\ : Odrv4
    port map (
            O => \N__5011\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__779\ : InMux
    port map (
            O => \N__5006\,
            I => \N__5002\
        );

    \I__778\ : InMux
    port map (
            O => \N__5005\,
            I => \N__4998\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5002\,
            I => \N__4995\
        );

    \I__776\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4992\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4998\,
            I => \N__4987\
        );

    \I__774\ : Span4Mux_h
    port map (
            O => \N__4995\,
            I => \N__4987\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4992\,
            I => \U712_CHIP_RAM.N_167\
        );

    \I__772\ : Odrv4
    port map (
            O => \N__4987\,
            I => \U712_CHIP_RAM.N_167\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__4982\,
            I => \N__4976\
        );

    \I__770\ : InMux
    port map (
            O => \N__4981\,
            I => \N__4972\
        );

    \I__769\ : InMux
    port map (
            O => \N__4980\,
            I => \N__4967\
        );

    \I__768\ : InMux
    port map (
            O => \N__4979\,
            I => \N__4967\
        );

    \I__767\ : InMux
    port map (
            O => \N__4976\,
            I => \N__4964\
        );

    \I__766\ : InMux
    port map (
            O => \N__4975\,
            I => \N__4961\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4972\,
            I => \N__4956\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4967\,
            I => \N__4953\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__4964\,
            I => \N__4948\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4961\,
            I => \N__4948\
        );

    \I__761\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4943\
        );

    \I__760\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4943\
        );

    \I__759\ : Span4Mux_v
    port map (
            O => \N__4956\,
            I => \N__4936\
        );

    \I__758\ : Span4Mux_h
    port map (
            O => \N__4953\,
            I => \N__4936\
        );

    \I__757\ : Span4Mux_v
    port map (
            O => \N__4948\,
            I => \N__4936\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__4943\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__4936\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__754\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4926\
        );

    \I__753\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4920\
        );

    \I__752\ : InMux
    port map (
            O => \N__4929\,
            I => \N__4917\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4926\,
            I => \N__4914\
        );

    \I__750\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4911\
        );

    \I__749\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4908\
        );

    \I__748\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4905\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__4920\,
            I => \N__4902\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4917\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1\
        );

    \I__745\ : Odrv4
    port map (
            O => \N__4914\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__4911\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__4908\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4905\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1\
        );

    \I__741\ : Odrv4
    port map (
            O => \N__4902\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1\
        );

    \I__740\ : InMux
    port map (
            O => \N__4889\,
            I => \N__4879\
        );

    \I__739\ : InMux
    port map (
            O => \N__4888\,
            I => \N__4872\
        );

    \I__738\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4872\
        );

    \I__737\ : InMux
    port map (
            O => \N__4886\,
            I => \N__4872\
        );

    \I__736\ : InMux
    port map (
            O => \N__4885\,
            I => \N__4865\
        );

    \I__735\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4865\
        );

    \I__734\ : InMux
    port map (
            O => \N__4883\,
            I => \N__4865\
        );

    \I__733\ : InMux
    port map (
            O => \N__4882\,
            I => \N__4862\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4879\,
            I => \N__4859\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4872\,
            I => \U712_CHIP_RAM.N_53\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4865\,
            I => \U712_CHIP_RAM.N_53\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__4862\,
            I => \U712_CHIP_RAM.N_53\
        );

    \I__728\ : Odrv4
    port map (
            O => \N__4859\,
            I => \U712_CHIP_RAM.N_53\
        );

    \I__727\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4847\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4847\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__725\ : CascadeMux
    port map (
            O => \N__4844\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_1_cascade_\
        );

    \I__724\ : CEMux
    port map (
            O => \N__4841\,
            I => \N__4837\
        );

    \I__723\ : CEMux
    port map (
            O => \N__4840\,
            I => \N__4834\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4837\,
            I => \N__4830\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4834\,
            I => \N__4827\
        );

    \I__720\ : CEMux
    port map (
            O => \N__4833\,
            I => \N__4824\
        );

    \I__719\ : Span4Mux_h
    port map (
            O => \N__4830\,
            I => \N__4821\
        );

    \I__718\ : Span4Mux_h
    port map (
            O => \N__4827\,
            I => \N__4818\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4824\,
            I => \N__4815\
        );

    \I__716\ : Span4Mux_h
    port map (
            O => \N__4821\,
            I => \N__4812\
        );

    \I__715\ : Span4Mux_h
    port map (
            O => \N__4818\,
            I => \N__4809\
        );

    \I__714\ : Span4Mux_v
    port map (
            O => \N__4815\,
            I => \N__4806\
        );

    \I__713\ : Odrv4
    port map (
            O => \N__4812\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__712\ : Odrv4
    port map (
            O => \N__4809\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__711\ : Odrv4
    port map (
            O => \N__4806\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__4799\,
            I => \U712_CHIP_RAM.N_196_cascade_\
        );

    \I__709\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4789\
        );

    \I__708\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4789\
        );

    \I__707\ : InMux
    port map (
            O => \N__4794\,
            I => \N__4786\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4789\,
            I => \N__4783\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__4786\,
            I => \U712_CHIP_RAM.N_315\
        );

    \I__704\ : Odrv4
    port map (
            O => \N__4783\,
            I => \U712_CHIP_RAM.N_315\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__4778\,
            I => \U712_CHIP_RAM.N_197_i_cascade_\
        );

    \I__702\ : InMux
    port map (
            O => \N__4775\,
            I => \N__4769\
        );

    \I__701\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4769\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4769\,
            I => \N__4766\
        );

    \I__699\ : Odrv4
    port map (
            O => \N__4766\,
            I => \U712_CHIP_RAM.N_233\
        );

    \I__698\ : InMux
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4760\,
            I => \N__4755\
        );

    \I__696\ : InMux
    port map (
            O => \N__4759\,
            I => \N__4750\
        );

    \I__695\ : InMux
    port map (
            O => \N__4758\,
            I => \N__4750\
        );

    \I__694\ : Odrv4
    port map (
            O => \N__4755\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8RZ0\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4750\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8RZ0\
        );

    \I__692\ : InMux
    port map (
            O => \N__4745\,
            I => \N__4741\
        );

    \I__691\ : InMux
    port map (
            O => \N__4744\,
            I => \N__4738\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4741\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__4738\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__688\ : InMux
    port map (
            O => \N__4733\,
            I => \N__4729\
        );

    \I__687\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4726\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4729\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4726\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__4721\,
            I => \N__4717\
        );

    \I__683\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4714\
        );

    \I__682\ : InMux
    port map (
            O => \N__4717\,
            I => \N__4711\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4714\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__4711\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__679\ : InMux
    port map (
            O => \N__4706\,
            I => \N__4702\
        );

    \I__678\ : InMux
    port map (
            O => \N__4705\,
            I => \N__4699\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4702\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__4699\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__675\ : CascadeMux
    port map (
            O => \N__4694\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1_cascade_\
        );

    \I__674\ : CEMux
    port map (
            O => \N__4691\,
            I => \N__4687\
        );

    \I__673\ : CEMux
    port map (
            O => \N__4690\,
            I => \N__4684\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4687\,
            I => \N__4681\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4684\,
            I => \N__4678\
        );

    \I__670\ : Odrv4
    port map (
            O => \N__4681\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\
        );

    \I__669\ : Odrv4
    port map (
            O => \N__4678\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\
        );

    \I__668\ : InMux
    port map (
            O => \N__4673\,
            I => \N__4669\
        );

    \I__667\ : InMux
    port map (
            O => \N__4672\,
            I => \N__4666\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__4669\,
            I => \N__4662\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4666\,
            I => \N__4659\
        );

    \I__664\ : InMux
    port map (
            O => \N__4665\,
            I => \N__4656\
        );

    \I__663\ : Odrv4
    port map (
            O => \N__4662\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__662\ : Odrv4
    port map (
            O => \N__4659\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4656\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__660\ : InMux
    port map (
            O => \N__4649\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__659\ : InMux
    port map (
            O => \N__4646\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__658\ : InMux
    port map (
            O => \N__4643\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__657\ : InMux
    port map (
            O => \N__4640\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__656\ : InMux
    port map (
            O => \N__4637\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__655\ : InMux
    port map (
            O => \N__4634\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__654\ : InMux
    port map (
            O => \N__4631\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__653\ : CascadeMux
    port map (
            O => \N__4628\,
            I => \U712_CHIP_RAM.N_230_cascade_\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__4625\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_0_cascade_\
        );

    \I__651\ : InMux
    port map (
            O => \N__4622\,
            I => \N__4619\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4619\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_1\
        );

    \I__649\ : InMux
    port map (
            O => \N__4616\,
            I => \N__4613\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4613\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_1\
        );

    \I__647\ : InMux
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__4607\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_a3_1_1\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__4604\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_cascade_\
        );

    \I__644\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4598\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4598\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__4595\,
            I => \U712_CHIP_RAM.N_285_cascade_\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__4592\,
            I => \N__4589\
        );

    \I__640\ : InMux
    port map (
            O => \N__4589\,
            I => \N__4586\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4586\,
            I => \N__4583\
        );

    \I__638\ : Odrv4
    port map (
            O => \N__4583\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_1\
        );

    \I__637\ : CascadeMux
    port map (
            O => \N__4580\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_1_cascade_\
        );

    \I__636\ : CascadeMux
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__635\ : InMux
    port map (
            O => \N__4574\,
            I => \N__4571\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__4571\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1\
        );

    \I__633\ : SRMux
    port map (
            O => \N__4568\,
            I => \N__4565\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__631\ : Span4Mux_h
    port map (
            O => \N__4562\,
            I => \N__4559\
        );

    \I__630\ : Odrv4
    port map (
            O => \N__4559\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__629\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4553\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__627\ : Span4Mux_v
    port map (
            O => \N__4550\,
            I => \N__4547\
        );

    \I__626\ : Span4Mux_h
    port map (
            O => \N__4547\,
            I => \N__4544\
        );

    \I__625\ : Sp12to4
    port map (
            O => \N__4544\,
            I => \N__4541\
        );

    \I__624\ : Odrv12
    port map (
            O => \N__4541\,
            I => \A_c_13\
        );

    \I__623\ : CascadeMux
    port map (
            O => \N__4538\,
            I => \N__4535\
        );

    \I__622\ : InMux
    port map (
            O => \N__4535\,
            I => \N__4532\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__4532\,
            I => \N__4529\
        );

    \I__620\ : Span12Mux_v
    port map (
            O => \N__4529\,
            I => \N__4526\
        );

    \I__619\ : Span12Mux_h
    port map (
            O => \N__4526\,
            I => \N__4523\
        );

    \I__618\ : Odrv12
    port map (
            O => \N__4523\,
            I => \A_c_6\
        );

    \I__617\ : InMux
    port map (
            O => \N__4520\,
            I => \N__4517\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__615\ : Span4Mux_h
    port map (
            O => \N__4514\,
            I => \N__4511\
        );

    \I__614\ : Sp12to4
    port map (
            O => \N__4511\,
            I => \N__4508\
        );

    \I__613\ : Span12Mux_v
    port map (
            O => \N__4508\,
            I => \N__4505\
        );

    \I__612\ : Odrv12
    port map (
            O => \N__4505\,
            I => \A_c_15\
        );

    \I__611\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4499\,
            I => \N__4496\
        );

    \I__609\ : Span12Mux_v
    port map (
            O => \N__4496\,
            I => \N__4493\
        );

    \I__608\ : Span12Mux_h
    port map (
            O => \N__4493\,
            I => \N__4490\
        );

    \I__607\ : Odrv12
    port map (
            O => \N__4490\,
            I => \A_c_8\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__4487\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\
        );

    \I__605\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4477\
        );

    \I__604\ : InMux
    port map (
            O => \N__4483\,
            I => \N__4477\
        );

    \I__603\ : InMux
    port map (
            O => \N__4482\,
            I => \N__4474\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4477\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIIGLS1Z0Z_0\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__4474\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIIGLS1Z0Z_0\
        );

    \I__600\ : CascadeMux
    port map (
            O => \N__4469\,
            I => \N__4466\
        );

    \I__599\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4458\
        );

    \I__598\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4458\
        );

    \I__597\ : InMux
    port map (
            O => \N__4464\,
            I => \N__4454\
        );

    \I__596\ : InMux
    port map (
            O => \N__4463\,
            I => \N__4451\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4458\,
            I => \N__4448\
        );

    \I__594\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4445\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4454\,
            I => \N__4440\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4451\,
            I => \N__4440\
        );

    \I__591\ : Odrv4
    port map (
            O => \N__4448\,
            I => \U712_CHIP_RAM.N_176\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__4445\,
            I => \U712_CHIP_RAM.N_176\
        );

    \I__589\ : Odrv4
    port map (
            O => \N__4440\,
            I => \U712_CHIP_RAM.N_176\
        );

    \I__588\ : InMux
    port map (
            O => \N__4433\,
            I => \N__4429\
        );

    \I__587\ : InMux
    port map (
            O => \N__4432\,
            I => \N__4426\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4429\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__4426\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__584\ : CascadeMux
    port map (
            O => \N__4421\,
            I => \U712_CHIP_RAM.N_167_cascade_\
        );

    \I__583\ : CEMux
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__4415\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_9_0_0\
        );

    \I__581\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4409\,
            I => \N__4405\
        );

    \I__579\ : InMux
    port map (
            O => \N__4408\,
            I => \N__4402\
        );

    \I__578\ : Odrv4
    port map (
            O => \N__4405\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__4402\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__576\ : InMux
    port map (
            O => \N__4397\,
            I => \N__4388\
        );

    \I__575\ : InMux
    port map (
            O => \N__4396\,
            I => \N__4388\
        );

    \I__574\ : InMux
    port map (
            O => \N__4395\,
            I => \N__4388\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4388\,
            I => \N__4385\
        );

    \I__572\ : Sp12to4
    port map (
            O => \N__4385\,
            I => \N__4382\
        );

    \I__571\ : Span12Mux_v
    port map (
            O => \N__4382\,
            I => \N__4379\
        );

    \I__570\ : Span12Mux_h
    port map (
            O => \N__4379\,
            I => \N__4376\
        );

    \I__569\ : Odrv12
    port map (
            O => \N__4376\,
            I => \SIZ_c_1\
        );

    \I__568\ : IoInMux
    port map (
            O => \N__4373\,
            I => \N__4370\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4370\,
            I => \N__4367\
        );

    \I__566\ : Span4Mux_s0_v
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__565\ : Sp12to4
    port map (
            O => \N__4364\,
            I => \N__4360\
        );

    \I__564\ : InMux
    port map (
            O => \N__4363\,
            I => \N__4357\
        );

    \I__563\ : Span12Mux_h
    port map (
            O => \N__4360\,
            I => \N__4354\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4357\,
            I => \N__4351\
        );

    \I__561\ : Odrv12
    port map (
            O => \N__4354\,
            I => \CONSTANT_ONE_NET\
        );

    \I__560\ : Odrv4
    port map (
            O => \N__4351\,
            I => \CONSTANT_ONE_NET\
        );

    \I__559\ : InMux
    port map (
            O => \N__4346\,
            I => \N__4343\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__4343\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__557\ : InMux
    port map (
            O => \N__4340\,
            I => \N__4337\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4337\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__4334\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1_cascade_\
        );

    \I__554\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4327\
        );

    \I__553\ : InMux
    port map (
            O => \N__4330\,
            I => \N__4324\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__4327\,
            I => \U712_CHIP_RAM.N_313\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__4324\,
            I => \U712_CHIP_RAM.N_313\
        );

    \I__550\ : InMux
    port map (
            O => \N__4319\,
            I => \N__4316\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4316\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__4313\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_9_0_cascade_\
        );

    \I__547\ : InMux
    port map (
            O => \N__4310\,
            I => \N__4305\
        );

    \I__546\ : InMux
    port map (
            O => \N__4309\,
            I => \N__4300\
        );

    \I__545\ : InMux
    port map (
            O => \N__4308\,
            I => \N__4300\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4305\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0_a3_0\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4300\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0_a3_0\
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__4295\,
            I => \U712_CHIP_RAM.N_232_cascade_\
        );

    \I__541\ : InMux
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4289\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0_a3_1\
        );

    \I__539\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4283\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4283\,
            I => \U712_CHIP_RAM.N_232\
        );

    \I__537\ : InMux
    port map (
            O => \N__4280\,
            I => \N__4276\
        );

    \I__536\ : InMux
    port map (
            O => \N__4279\,
            I => \N__4273\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4276\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__4273\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__533\ : InMux
    port map (
            O => \N__4268\,
            I => \N__4265\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__4265\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0\
        );

    \I__531\ : InMux
    port map (
            O => \N__4262\,
            I => \N__4259\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__4259\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_i_i_a3_0\
        );

    \I__529\ : CascadeMux
    port map (
            O => \N__4256\,
            I => \N__4253\
        );

    \I__528\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4250\,
            I => \N__4247\
        );

    \I__526\ : Odrv4
    port map (
            O => \N__4247\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__525\ : CascadeMux
    port map (
            O => \N__4244\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_cascade_\
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__4241\,
            I => \U712_CHIP_RAM.CLK_EN_e_1_cascade_\
        );

    \I__523\ : IoInMux
    port map (
            O => \N__4238\,
            I => \N__4235\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4235\,
            I => \N__4232\
        );

    \I__521\ : IoSpan4Mux
    port map (
            O => \N__4232\,
            I => \N__4229\
        );

    \I__520\ : Sp12to4
    port map (
            O => \N__4229\,
            I => \N__4226\
        );

    \I__519\ : Span12Mux_s7_h
    port map (
            O => \N__4226\,
            I => \N__4223\
        );

    \I__518\ : Span12Mux_h
    port map (
            O => \N__4223\,
            I => \N__4219\
        );

    \I__517\ : InMux
    port map (
            O => \N__4222\,
            I => \N__4216\
        );

    \I__516\ : Odrv12
    port map (
            O => \N__4219\,
            I => \CLK_EN_c\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4216\,
            I => \CLK_EN_c\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__4211\,
            I => \U712_CHIP_RAM.N_176_cascade_\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__4208\,
            I => \U712_CHIP_RAM.N_166_cascade_\
        );

    \I__512\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4202\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4202\,
            I => \N__4199\
        );

    \I__510\ : Span12Mux_h
    port map (
            O => \N__4199\,
            I => \N__4196\
        );

    \I__509\ : Odrv12
    port map (
            O => \N__4196\,
            I => \A_c_11\
        );

    \I__508\ : InMux
    port map (
            O => \N__4193\,
            I => \N__4190\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__4190\,
            I => \N__4187\
        );

    \I__506\ : Span4Mux_h
    port map (
            O => \N__4187\,
            I => \N__4184\
        );

    \I__505\ : Sp12to4
    port map (
            O => \N__4184\,
            I => \N__4181\
        );

    \I__504\ : Span12Mux_v
    port map (
            O => \N__4181\,
            I => \N__4178\
        );

    \I__503\ : Odrv12
    port map (
            O => \N__4178\,
            I => \A_c_4\
        );

    \I__502\ : InMux
    port map (
            O => \N__4175\,
            I => \N__4172\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__4172\,
            I => \N__4169\
        );

    \I__500\ : Span4Mux_h
    port map (
            O => \N__4169\,
            I => \N__4166\
        );

    \I__499\ : Span4Mux_v
    port map (
            O => \N__4166\,
            I => \N__4163\
        );

    \I__498\ : Sp12to4
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__497\ : Odrv12
    port map (
            O => \N__4160\,
            I => \A_c_9\
        );

    \I__496\ : InMux
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__494\ : Span4Mux_v
    port map (
            O => \N__4151\,
            I => \N__4148\
        );

    \I__493\ : Sp12to4
    port map (
            O => \N__4148\,
            I => \N__4145\
        );

    \I__492\ : Span12Mux_h
    port map (
            O => \N__4145\,
            I => \N__4142\
        );

    \I__491\ : Span12Mux_v
    port map (
            O => \N__4142\,
            I => \N__4139\
        );

    \I__490\ : Odrv12
    port map (
            O => \N__4139\,
            I => \A_c_2\
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__4136\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_1_cascade_\
        );

    \I__488\ : InMux
    port map (
            O => \N__4133\,
            I => \N__4130\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4130\,
            I => \N__4127\
        );

    \I__486\ : Span4Mux_v
    port map (
            O => \N__4127\,
            I => \N__4124\
        );

    \I__485\ : Span4Mux_h
    port map (
            O => \N__4124\,
            I => \N__4121\
        );

    \I__484\ : Sp12to4
    port map (
            O => \N__4121\,
            I => \N__4118\
        );

    \I__483\ : Odrv12
    port map (
            O => \N__4118\,
            I => \A_c_12\
        );

    \I__482\ : InMux
    port map (
            O => \N__4115\,
            I => \N__4112\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4112\,
            I => \N__4109\
        );

    \I__480\ : Span4Mux_v
    port map (
            O => \N__4109\,
            I => \N__4106\
        );

    \I__479\ : Span4Mux_v
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__478\ : Sp12to4
    port map (
            O => \N__4103\,
            I => \N__4100\
        );

    \I__477\ : Odrv12
    port map (
            O => \N__4100\,
            I => \A_c_5\
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__4097\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2_cascade_\
        );

    \I__475\ : InMux
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4091\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_0\
        );

    \I__473\ : InMux
    port map (
            O => \N__4088\,
            I => \N__4085\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4085\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_1_0\
        );

    \I__471\ : CascadeMux
    port map (
            O => \N__4082\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_\
        );

    \I__470\ : InMux
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4076\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_2\
        );

    \I__468\ : InMux
    port map (
            O => \N__4073\,
            I => \N__4070\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__466\ : Span4Mux_h
    port map (
            O => \N__4067\,
            I => \N__4064\
        );

    \I__465\ : Sp12to4
    port map (
            O => \N__4064\,
            I => \N__4061\
        );

    \I__464\ : Span12Mux_v
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__463\ : Odrv12
    port map (
            O => \N__4058\,
            I => \RAMSPACEn_c\
        );

    \I__462\ : InMux
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4052\,
            I => \N__4049\
        );

    \I__460\ : Odrv4
    port map (
            O => \N__4049\,
            I => \U712_CHIP_RAM.un5_DMA_CYCLE_START_0\
        );

    \I__459\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4042\
        );

    \I__458\ : InMux
    port map (
            O => \N__4045\,
            I => \N__4039\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4042\,
            I => \N__4035\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__4039\,
            I => \N__4032\
        );

    \I__455\ : InMux
    port map (
            O => \N__4038\,
            I => \N__4029\
        );

    \I__454\ : Odrv12
    port map (
            O => \N__4035\,
            I => \REG_CYCLEm\
        );

    \I__453\ : Odrv4
    port map (
            O => \N__4032\,
            I => \REG_CYCLEm\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4029\,
            I => \REG_CYCLEm\
        );

    \I__451\ : IoInMux
    port map (
            O => \N__4022\,
            I => \N__4019\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4019\,
            I => \N__4016\
        );

    \I__449\ : Span4Mux_s0_v
    port map (
            O => \N__4016\,
            I => \N__4013\
        );

    \I__448\ : Sp12to4
    port map (
            O => \N__4013\,
            I => \N__4010\
        );

    \I__447\ : Span12Mux_s9_h
    port map (
            O => \N__4010\,
            I => \N__4007\
        );

    \I__446\ : Span12Mux_v
    port map (
            O => \N__4007\,
            I => \N__4004\
        );

    \I__445\ : Odrv12
    port map (
            O => \N__4004\,
            I => \DRDENn_c\
        );

    \I__444\ : InMux
    port map (
            O => \N__4001\,
            I => \N__3998\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__3998\,
            I => \N__3995\
        );

    \I__442\ : Span4Mux_h
    port map (
            O => \N__3995\,
            I => \N__3992\
        );

    \I__441\ : Sp12to4
    port map (
            O => \N__3992\,
            I => \N__3989\
        );

    \I__440\ : Span12Mux_v
    port map (
            O => \N__3989\,
            I => \N__3986\
        );

    \I__439\ : Odrv12
    port map (
            O => \N__3986\,
            I => \A_c_16\
        );

    \I__438\ : InMux
    port map (
            O => \N__3983\,
            I => \N__3980\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__3980\,
            I => \N__3977\
        );

    \I__436\ : Span4Mux_v
    port map (
            O => \N__3977\,
            I => \N__3974\
        );

    \I__435\ : Span4Mux_v
    port map (
            O => \N__3974\,
            I => \N__3971\
        );

    \I__434\ : Sp12to4
    port map (
            O => \N__3971\,
            I => \N__3968\
        );

    \I__433\ : Span12Mux_h
    port map (
            O => \N__3968\,
            I => \N__3965\
        );

    \I__432\ : Odrv12
    port map (
            O => \N__3965\,
            I => \A_c_18\
        );

    \I__431\ : InMux
    port map (
            O => \N__3962\,
            I => \N__3958\
        );

    \I__430\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3955\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3958\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3955\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__427\ : InMux
    port map (
            O => \N__3950\,
            I => \N__3947\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__3947\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__3944\,
            I => \N__3940\
        );

    \I__424\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3937\
        );

    \I__423\ : InMux
    port map (
            O => \N__3940\,
            I => \N__3934\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3937\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3934\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__420\ : InMux
    port map (
            O => \N__3929\,
            I => \N__3926\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3926\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__418\ : IoInMux
    port map (
            O => \N__3923\,
            I => \N__3920\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3920\,
            I => \N__3917\
        );

    \I__416\ : Span12Mux_s4_v
    port map (
            O => \N__3917\,
            I => \N__3913\
        );

    \I__415\ : InMux
    port map (
            O => \N__3916\,
            I => \N__3910\
        );

    \I__414\ : Odrv12
    port map (
            O => \N__3913\,
            I => \DBDIR_c\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__3910\,
            I => \DBDIR_c\
        );

    \I__412\ : InMux
    port map (
            O => \N__3905\,
            I => \N__3902\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__3902\,
            I => \N__3899\
        );

    \I__410\ : Span4Mux_v
    port map (
            O => \N__3899\,
            I => \N__3896\
        );

    \I__409\ : Odrv4
    port map (
            O => \N__3896\,
            I => \TACK_EN_i_ess\
        );

    \I__408\ : IoInMux
    port map (
            O => \N__3893\,
            I => \N__3890\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__3890\,
            I => \N__3887\
        );

    \I__406\ : Span12Mux_s5_v
    port map (
            O => \N__3887\,
            I => \N__3884\
        );

    \I__405\ : Odrv12
    port map (
            O => \N__3884\,
            I => \VBENn_c\
        );

    \I__404\ : InMux
    port map (
            O => \N__3881\,
            I => \N__3878\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__3878\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1\
        );

    \I__402\ : CascadeMux
    port map (
            O => \N__3875\,
            I => \N__3869\
        );

    \I__401\ : InMux
    port map (
            O => \N__3874\,
            I => \N__3866\
        );

    \I__400\ : InMux
    port map (
            O => \N__3873\,
            I => \N__3859\
        );

    \I__399\ : InMux
    port map (
            O => \N__3872\,
            I => \N__3859\
        );

    \I__398\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3859\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__3866\,
            I => \N__3856\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3859\,
            I => \N__3853\
        );

    \I__395\ : Span12Mux_v
    port map (
            O => \N__3856\,
            I => \N__3850\
        );

    \I__394\ : Span12Mux_h
    port map (
            O => \N__3853\,
            I => \N__3847\
        );

    \I__393\ : Span12Mux_h
    port map (
            O => \N__3850\,
            I => \N__3842\
        );

    \I__392\ : Span12Mux_v
    port map (
            O => \N__3847\,
            I => \N__3842\
        );

    \I__391\ : Odrv12
    port map (
            O => \N__3842\,
            I => \CLK40_PLL_i\
        );

    \I__390\ : InMux
    port map (
            O => \N__3839\,
            I => \N__3835\
        );

    \I__389\ : InMux
    port map (
            O => \N__3838\,
            I => \N__3832\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3835\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__3832\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__386\ : InMux
    port map (
            O => \N__3827\,
            I => \N__3823\
        );

    \I__385\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3820\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3823\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3820\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__382\ : InMux
    port map (
            O => \N__3815\,
            I => \bfn_7_7_0_\
        );

    \I__381\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3808\
        );

    \I__380\ : InMux
    port map (
            O => \N__3811\,
            I => \N__3805\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__3808\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3805\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__377\ : InMux
    port map (
            O => \N__3800\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__376\ : InMux
    port map (
            O => \N__3797\,
            I => \N__3793\
        );

    \I__375\ : InMux
    port map (
            O => \N__3796\,
            I => \N__3790\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3793\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__3790\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__372\ : InMux
    port map (
            O => \N__3785\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__371\ : InMux
    port map (
            O => \N__3782\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__370\ : CascadeMux
    port map (
            O => \N__3779\,
            I => \N__3775\
        );

    \I__369\ : InMux
    port map (
            O => \N__3778\,
            I => \N__3772\
        );

    \I__368\ : InMux
    port map (
            O => \N__3775\,
            I => \N__3769\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__3772\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__3769\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__365\ : InMux
    port map (
            O => \N__3764\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__364\ : InMux
    port map (
            O => \N__3761\,
            I => \N__3757\
        );

    \I__363\ : InMux
    port map (
            O => \N__3760\,
            I => \N__3754\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__3757\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__3754\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__360\ : InMux
    port map (
            O => \N__3749\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__359\ : InMux
    port map (
            O => \N__3746\,
            I => \N__3742\
        );

    \I__358\ : InMux
    port map (
            O => \N__3745\,
            I => \N__3739\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__3742\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__3739\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__355\ : InMux
    port map (
            O => \N__3734\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__354\ : InMux
    port map (
            O => \N__3731\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__353\ : IoInMux
    port map (
            O => \N__3728\,
            I => \N__3725\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__3725\,
            I => \N__3722\
        );

    \I__351\ : Span4Mux_s2_v
    port map (
            O => \N__3722\,
            I => \N__3719\
        );

    \I__350\ : Span4Mux_v
    port map (
            O => \N__3719\,
            I => \N__3716\
        );

    \I__349\ : Span4Mux_h
    port map (
            O => \N__3716\,
            I => \N__3713\
        );

    \I__348\ : Odrv4
    port map (
            O => \N__3713\,
            I => \CLK80_PLL_i_i\
        );

    \I__347\ : InMux
    port map (
            O => \N__3710\,
            I => \N__3707\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__3707\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\
        );

    \I__345\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3697\
        );

    \I__344\ : InMux
    port map (
            O => \N__3703\,
            I => \N__3697\
        );

    \I__343\ : InMux
    port map (
            O => \N__3702\,
            I => \N__3694\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3697\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__3694\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__340\ : IoInMux
    port map (
            O => \N__3689\,
            I => \N__3686\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__3686\,
            I => \N__3683\
        );

    \I__338\ : Span4Mux_s3_h
    port map (
            O => \N__3683\,
            I => \N__3680\
        );

    \I__337\ : Span4Mux_h
    port map (
            O => \N__3680\,
            I => \N__3677\
        );

    \I__336\ : Sp12to4
    port map (
            O => \N__3677\,
            I => \N__3674\
        );

    \I__335\ : Span12Mux_v
    port map (
            O => \N__3674\,
            I => \N__3670\
        );

    \I__334\ : InMux
    port map (
            O => \N__3673\,
            I => \N__3667\
        );

    \I__333\ : Odrv12
    port map (
            O => \N__3670\,
            I => \TACK_OUTn\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__3667\,
            I => \TACK_OUTn\
        );

    \I__331\ : InMux
    port map (
            O => \N__3662\,
            I => \N__3650\
        );

    \I__330\ : InMux
    port map (
            O => \N__3661\,
            I => \N__3650\
        );

    \I__329\ : InMux
    port map (
            O => \N__3660\,
            I => \N__3650\
        );

    \I__328\ : InMux
    port map (
            O => \N__3659\,
            I => \N__3650\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__3650\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__326\ : IoInMux
    port map (
            O => \N__3647\,
            I => \N__3644\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__3644\,
            I => \N__3641\
        );

    \I__324\ : Odrv12
    port map (
            O => \N__3641\,
            I => \CLK40_PLL_i_i\
        );

    \I__323\ : IoInMux
    port map (
            O => \N__3638\,
            I => \N__3635\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__3635\,
            I => \N__3632\
        );

    \I__321\ : Span4Mux_s3_h
    port map (
            O => \N__3632\,
            I => \N__3629\
        );

    \I__320\ : Span4Mux_v
    port map (
            O => \N__3629\,
            I => \N__3626\
        );

    \I__319\ : Span4Mux_v
    port map (
            O => \N__3626\,
            I => \N__3623\
        );

    \I__318\ : Odrv4
    port map (
            O => \N__3623\,
            I => \N_981_i\
        );

    \I__317\ : IoInMux
    port map (
            O => \N__3620\,
            I => \N__3617\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__3617\,
            I => \N__3614\
        );

    \I__315\ : Span4Mux_s0_v
    port map (
            O => \N__3614\,
            I => \N__3611\
        );

    \I__314\ : Span4Mux_v
    port map (
            O => \N__3611\,
            I => \N__3608\
        );

    \I__313\ : Sp12to4
    port map (
            O => \N__3608\,
            I => \N__3605\
        );

    \I__312\ : Span12Mux_h
    port map (
            O => \N__3605\,
            I => \N__3602\
        );

    \I__311\ : Span12Mux_v
    port map (
            O => \N__3602\,
            I => \N__3599\
        );

    \I__310\ : Odrv12
    port map (
            O => \N__3599\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__8473\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__8475\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__8476\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__8471\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__8472\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__8474\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8354\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7208\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7253\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLK40_OUT_obuf_RNO_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3874\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3905\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_981_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8840\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__3796\,
            in1 => \N__3811\,
            in2 => \N__3779\,
            in3 => \N__3826\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3745\,
            in2 => \_gnd_net_\,
            in3 => \N__3760\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3702\,
            in2 => \_gnd_net_\,
            in3 => \N__3838\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000110000"
        )
    port map (
            in0 => \N__3710\,
            in1 => \N__3659\,
            in2 => \N__6788\,
            in3 => \N__6540\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8836\,
            ce => 'H',
            sr => \N__9254\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3704\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8836\,
            ce => 'H',
            sr => \N__9254\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3839\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8836\,
            ce => 'H',
            sr => \N__9254\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110001000"
        )
    port map (
            in0 => \N__3662\,
            in1 => \N__3872\,
            in2 => \N__6542\,
            in3 => \N__6766\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8836\,
            ce => 'H',
            sr => \N__9254\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110100010"
        )
    port map (
            in0 => \N__3673\,
            in1 => \N__3661\,
            in2 => \N__3875\,
            in3 => \N__3703\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8836\,
            ce => 'H',
            sr => \N__9254\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__3660\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3873\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8836\,
            ce => 'H',
            sr => \N__9254\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3827\,
            in2 => \_gnd_net_\,
            in3 => \N__3815\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__8470\,
            ce => 'H',
            sr => \N__4568\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3812\,
            in2 => \_gnd_net_\,
            in3 => \N__3800\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__8470\,
            ce => 'H',
            sr => \N__4568\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3797\,
            in2 => \_gnd_net_\,
            in3 => \N__3785\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__8470\,
            ce => 'H',
            sr => \N__4568\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3962\,
            in2 => \_gnd_net_\,
            in3 => \N__3782\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__8470\,
            ce => 'H',
            sr => \N__4568\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3778\,
            in2 => \_gnd_net_\,
            in3 => \N__3764\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__8470\,
            ce => 'H',
            sr => \N__4568\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3761\,
            in2 => \_gnd_net_\,
            in3 => \N__3749\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__8470\,
            ce => 'H',
            sr => \N__4568\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3746\,
            in2 => \_gnd_net_\,
            in3 => \N__3734\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__8470\,
            ce => 'H',
            sr => \N__4568\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3943\,
            in2 => \_gnd_net_\,
            in3 => \N__3731\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8470\,
            ce => 'H',
            sr => \N__4568\
        );

    \U712_CHIP_RAM.REFRESH_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111111011"
        )
    port map (
            in0 => \N__3961\,
            in1 => \N__3950\,
            in2 => \N__3944\,
            in3 => \N__3929\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8824\,
            ce => 'H',
            sr => \N__9265\
        );

    \U712_CHIP_RAM.DBDIR_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__6445\,
            in1 => \N__3916\,
            in2 => \_gnd_net_\,
            in3 => \N__4280\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8829\,
            ce => 'H',
            sr => \N__9260\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__8429\,
            in1 => \N__6765\,
            in2 => \_gnd_net_\,
            in3 => \N__6541\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8835\,
            ce => \N__6743\,
            sr => \N__9244\
        );

    \U712_BUFFERS.un1_VBENn_0_a3_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4046\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7896\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000101011"
        )
    port map (
            in0 => \N__6060\,
            in1 => \N__6188\,
            in2 => \N__6323\,
            in3 => \N__3881\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000111"
        )
    port map (
            in0 => \N__4959\,
            in1 => \N__5143\,
            in2 => \N__6728\,
            in3 => \N__6380\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000001100"
        )
    port map (
            in0 => \N__6381\,
            in1 => \N__8433\,
            in2 => \N__5154\,
            in3 => \N__4960\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_i_i_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__4079\,
            in1 => \N__5315\,
            in2 => \N__6396\,
            in3 => \N__4055\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8825\,
            ce => 'H',
            sr => \N__9255\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4930\,
            in1 => \N__6376\,
            in2 => \_gnd_net_\,
            in3 => \N__5133\,
            lcout => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011111110000"
        )
    port map (
            in0 => \N__4310\,
            in1 => \N__4673\,
            in2 => \N__4082\,
            in3 => \N__5316\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8825\,
            ce => 'H',
            sr => \N__9255\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6181\,
            in1 => \N__6061\,
            in2 => \N__5153\,
            in3 => \N__6316\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_2_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4412\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8830\,
            ce => 'H',
            sr => \N__9245\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010100"
        )
    port map (
            in0 => \N__7564\,
            in1 => \N__7021\,
            in2 => \N__5933\,
            in3 => \N__7051\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8830\,
            ce => 'H',
            sr => \N__9245\
        );

    \U712_CHIP_RAM.DBENn_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110001011101110"
        )
    port map (
            in0 => \N__5619\,
            in1 => \N__4268\,
            in2 => \N__6089\,
            in3 => \N__8534\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8830\,
            ce => 'H',
            sr => \N__9245\
        );

    \U712_REG_SM.REG_CYCLE_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101110"
        )
    port map (
            in0 => \N__7489\,
            in1 => \N__4038\,
            in2 => \N__7022\,
            in3 => \N__7511\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8833\,
            ce => 'H',
            sr => \N__9235\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__4073\,
            in1 => \N__7824\,
            in2 => \N__7616\,
            in3 => \N__4433\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8833\,
            ce => 'H',
            sr => \N__9235\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4408\,
            in2 => \_gnd_net_\,
            in3 => \N__5021\,
            lcout => \U712_CHIP_RAM.un5_DMA_CYCLE_START_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_0_a3_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4045\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4001\,
            in1 => \N__3983\,
            in2 => \_gnd_net_\,
            in3 => \N__7432\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7396\,
            in1 => \N__4205\,
            in2 => \_gnd_net_\,
            in3 => \N__4193\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4363\,
            in2 => \_gnd_net_\,
            in3 => \N__6077\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4175\,
            in1 => \N__4157\,
            in2 => \_gnd_net_\,
            in3 => \N__7395\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5971\,
            in2 => \_gnd_net_\,
            in3 => \N__4094\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111011"
        )
    port map (
            in0 => \N__4483\,
            in1 => \N__4465\,
            in2 => \N__4136\,
            in3 => \N__6321\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8817\,
            ce => \N__4691\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4133\,
            in1 => \N__4115\,
            in2 => \_gnd_net_\,
            in3 => \N__7391\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6054\,
            in1 => \N__4463\,
            in2 => \_gnd_net_\,
            in3 => \N__5240\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__6320\,
            in1 => \N__6055\,
            in2 => \N__4097\,
            in3 => \N__5156\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__5972\,
            in1 => \N__4088\,
            in2 => \N__4469\,
            in3 => \N__4484\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8817\,
            ce => \N__4691\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__4262\,
            in1 => \N__4929\,
            in2 => \N__4256\,
            in3 => \N__4889\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8820\,
            ce => \N__4833\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4763\,
            in1 => \N__6305\,
            in2 => \N__5191\,
            in3 => \N__5057\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_a3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6267\,
            in1 => \N__6175\,
            in2 => \_gnd_net_\,
            in3 => \N__4457\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__6611\,
            in1 => \N__4222\,
            in2 => \N__4244\,
            in3 => \N__6044\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CLK_EN_e_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__5056\,
            in1 => \N__4331\,
            in2 => \N__4241\,
            in3 => \N__6206\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8822\,
            ce => 'H',
            sr => \N__9246\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6691\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5122\,
            lcout => \U712_CHIP_RAM.N_176\,
            ltout => \U712_CHIP_RAM.N_176_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_4_0_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000111011"
        )
    port map (
            in0 => \N__6266\,
            in1 => \N__5137\,
            in2 => \N__4211\,
            in3 => \N__5239\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6157\,
            in2 => \_gnd_net_\,
            in3 => \N__6265\,
            lcout => \U712_CHIP_RAM.N_166\,
            ltout => \U712_CHIP_RAM.N_166_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6043\,
            in1 => \N__6692\,
            in2 => \N__4208\,
            in3 => \N__6610\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIVLD65_0_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4975\,
            in1 => \N__6375\,
            in2 => \N__4334\,
            in3 => \N__5005\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIH7LR1_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010010000000"
        )
    port map (
            in0 => \N__6695\,
            in1 => \N__4330\,
            in2 => \N__6297\,
            in3 => \N__5043\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR9AQ_3_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5113\,
            in2 => \_gnd_net_\,
            in3 => \N__6151\,
            lcout => \U712_CHIP_RAM.N_313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__4665\,
            in1 => \N__4309\,
            in2 => \N__5141\,
            in3 => \N__4319\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9286\,
            in1 => \_gnd_net_\,
            in2 => \N__4313\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_9_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6084\,
            in2 => \N__6627\,
            in3 => \N__4308\,
            lcout => \U712_CHIP_RAM.N_232\,
            ltout => \U712_CHIP_RAM.N_232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__4794\,
            in1 => \N__8443\,
            in2 => \N__4295\,
            in3 => \N__4924\,
            lcout => \U712_CHIP_RAM.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__6696\,
            in1 => \N__4292\,
            in2 => \N__6628\,
            in3 => \N__5140\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8826\,
            ce => 'H',
            sr => \N__9236\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4286\,
            in2 => \_gnd_net_\,
            in3 => \N__4279\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4432\,
            in2 => \_gnd_net_\,
            in3 => \N__6493\,
            lcout => \U712_CHIP_RAM.N_167\,
            ltout => \U712_CHIP_RAM.N_167_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__4981\,
            in1 => \N__6401\,
            in2 => \N__4421\,
            in3 => \N__4931\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8831\,
            ce => \N__4418\,
            sr => \N__9232\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5020\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8834\,
            ce => 'H',
            sr => \N__9228\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__7884\,
            in1 => \N__8276\,
            in2 => \_gnd_net_\,
            in3 => \N__4397\,
            lcout => \U712_BYTE_ENABLE.N_265\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__8313\,
            in1 => \N__5452\,
            in2 => \N__7914\,
            in3 => \N__4396\,
            lcout => \U712_BYTE_ENABLE.N_268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__8312\,
            in1 => \N__5451\,
            in2 => \N__7913\,
            in3 => \N__4395\,
            lcout => \U712_BYTE_ENABLE.N_272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__7912\,
            in1 => \N__4346\,
            in2 => \N__7454\,
            in3 => \N__8939\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__7910\,
            in1 => \N__4340\,
            in2 => \N__7431\,
            in3 => \N__8585\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIIGLS1_0_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__8444\,
            in1 => \N__6078\,
            in2 => \_gnd_net_\,
            in3 => \N__5242\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNIIGLS1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8050\,
            in1 => \N__7366\,
            in2 => \N__8187\,
            in3 => \N__8132\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_2_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__8133\,
            in1 => \N__8051\,
            in2 => \_gnd_net_\,
            in3 => \N__7386\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__4556\,
            in1 => \_gnd_net_\,
            in2 => \N__4538\,
            in3 => \N__7387\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4520\,
            in1 => \N__4502\,
            in2 => \_gnd_net_\,
            in3 => \N__7367\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__7368\,
            in1 => \N__7911\,
            in2 => \N__4487\,
            in3 => \N__9038\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6177\,
            in1 => \N__6056\,
            in2 => \_gnd_net_\,
            in3 => \N__6718\,
            lcout => \U712_CHIP_RAM.N_258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101011"
        )
    port map (
            in0 => \N__4482\,
            in1 => \N__4464\,
            in2 => \N__6322\,
            in3 => \N__4622\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8814\,
            ce => \N__4690\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6041\,
            in2 => \_gnd_net_\,
            in3 => \N__6176\,
            lcout => \U712_CHIP_RAM.N_206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6042\,
            in1 => \N__5241\,
            in2 => \_gnd_net_\,
            in3 => \N__5155\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_230_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__6719\,
            in1 => \N__5187\,
            in2 => \N__4628\,
            in3 => \N__6312\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__5964\,
            in1 => \_gnd_net_\,
            in2 => \N__4625\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIGGM16_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__4980\,
            in1 => \N__4923\,
            in2 => \N__4592\,
            in3 => \N__6403\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__8436\,
            in1 => \N__4775\,
            in2 => \N__4577\,
            in3 => \N__4796\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4672\,
            in1 => \N__4616\,
            in2 => \_gnd_net_\,
            in3 => \N__8437\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__4610\,
            in1 => \N__6714\,
            in2 => \N__4604\,
            in3 => \N__6629\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_285_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4601\,
            in2 => \N__4595\,
            in3 => \N__8131\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHHIB1_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8438\,
            in1 => \N__5006\,
            in2 => \_gnd_net_\,
            in3 => \N__5142\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_1\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIGNOI5_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4979\,
            in1 => \N__6402\,
            in2 => \N__4580\,
            in3 => \N__6202\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITE99E_3_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__8439\,
            in1 => \N__4774\,
            in2 => \N__4694\,
            in3 => \N__4795\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6053\,
            in2 => \_gnd_net_\,
            in3 => \N__6615\,
            lcout => \U712_CHIP_RAM.N_314\,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4886\,
            in1 => \N__6707\,
            in2 => \_gnd_net_\,
            in3 => \N__4649\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__8821\,
            ce => \N__4840\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6295\,
            in2 => \_gnd_net_\,
            in3 => \N__4646\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4887\,
            in1 => \N__6185\,
            in2 => \_gnd_net_\,
            in3 => \N__4643\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__8821\,
            ce => \N__4840\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4883\,
            in1 => \N__4706\,
            in2 => \_gnd_net_\,
            in3 => \N__4640\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__8821\,
            ce => \N__4840\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4888\,
            in1 => \N__4733\,
            in2 => \_gnd_net_\,
            in3 => \N__4637\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__8821\,
            ce => \N__4840\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4884\,
            in1 => \N__4720\,
            in2 => \_gnd_net_\,
            in3 => \N__4634\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__8821\,
            ce => \N__4840\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__4745\,
            in1 => \N__4885\,
            in2 => \_gnd_net_\,
            in3 => \N__4631\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8821\,
            ce => \N__4840\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIVLD65_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110100000000"
        )
    port map (
            in0 => \N__5001\,
            in1 => \N__6404\,
            in2 => \N__4982\,
            in3 => \N__4925\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_1\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__4882\,
            in1 => \N__4850\,
            in2 => \N__4844\,
            in3 => \N__4759\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8823\,
            ce => \N__4841\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000001000"
        )
    port map (
            in0 => \N__5118\,
            in1 => \N__6694\,
            in2 => \N__6187\,
            in3 => \N__6269\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_196_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6079\,
            in2 => \N__4799\,
            in3 => \N__6613\,
            lcout => \U712_CHIP_RAM.N_315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6693\,
            in2 => \_gnd_net_\,
            in3 => \N__6268\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_197_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__6161\,
            in1 => \N__4758\,
            in2 => \N__4778\,
            in3 => \N__6614\,
            lcout => \U712_CHIP_RAM.N_233\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5117\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8435\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8RZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4744\,
            in1 => \N__4732\,
            in2 => \N__4721\,
            in3 => \N__4705\,
            lcout => \U712_CHIP_RAM.N_165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_6_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5044\,
            in2 => \_gnd_net_\,
            in3 => \N__6720\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_219_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111010101"
        )
    port map (
            in0 => \N__5138\,
            in1 => \N__6186\,
            in2 => \N__5249\,
            in3 => \N__6296\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_7_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__5246\,
            in1 => \N__5963\,
            in2 => \N__5207\,
            in3 => \N__5204\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111001010"
        )
    port map (
            in0 => \N__6098\,
            in1 => \N__6556\,
            in2 => \N__5195\,
            in3 => \N__6563\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8827\,
            ce => 'H',
            sr => \N__9229\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_5_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5045\,
            in1 => \N__5192\,
            in2 => \N__6298\,
            in3 => \N__7811\,
            lcout => \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__6332\,
            in1 => \N__5046\,
            in2 => \N__5165\,
            in3 => \N__5139\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8827\,
            ce => 'H',
            sr => \N__9229\
        );

    \DBR_SYNC_1_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6962\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8832\,
            ce => 'H',
            sr => \N__9222\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5526\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5390\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8832\,
            ce => 'H',
            sr => \N__9222\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0_0_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__5334\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5634\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0_0_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5635\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5335\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_185_i_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__5402\,
            in1 => \N__5415\,
            in2 => \N__5539\,
            in3 => \N__5603\,
            lcout => \N_185_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5458\,
            in1 => \N__8326\,
            in2 => \_gnd_net_\,
            in3 => \N__7885\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_270_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_186_i_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__5416\,
            in1 => \N__5488\,
            in2 => \N__5573\,
            in3 => \N__5389\,
            lcout => \N_186_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_187_i_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__5417\,
            in1 => \N__5546\,
            in2 => \N__5540\,
            in3 => \N__5489\,
            lcout => \N_187_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__5459\,
            in1 => \N__8327\,
            in2 => \_gnd_net_\,
            in3 => \N__7886\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_266_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_184_i_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__5414\,
            in1 => \N__5401\,
            in2 => \N__5393\,
            in3 => \N__5388\,
            lcout => \N_184_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_i_m2_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__6481\,
            in1 => \N__6444\,
            in2 => \_gnd_net_\,
            in3 => \N__5342\,
            lcout => \DRDDIR_i_m2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__7306\,
            in1 => \N__8573\,
            in2 => \N__6884\,
            in3 => \N__5276\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8806\,
            ce => \N__8724\,
            sr => \N__9261\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__7307\,
            in1 => \N__6881\,
            in2 => \N__9410\,
            in3 => \N__5747\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8806\,
            ce => \N__8724\,
            sr => \N__9261\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__7299\,
            in1 => \N__7274\,
            in2 => \N__6882\,
            in3 => \N__5720\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8808\,
            ce => \N__8703\,
            sr => \N__9256\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__7920\,
            in1 => \N__5690\,
            in2 => \N__7464\,
            in3 => \N__9092\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__7298\,
            in1 => \N__6871\,
            in2 => \N__5684\,
            in3 => \N__7265\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8808\,
            ce => \N__8703\,
            sr => \N__9256\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110111011"
        )
    port map (
            in0 => \N__8669\,
            in1 => \N__7956\,
            in2 => \N__5915\,
            in3 => \N__7888\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111101"
        )
    port map (
            in0 => \N__8126\,
            in1 => \N__8064\,
            in2 => \N__7445\,
            in3 => \N__8181\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9287\,
            in1 => \_gnd_net_\,
            in2 => \N__5657\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_2_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8063\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8127\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__7890\,
            in1 => \N__5654\,
            in2 => \N__7446\,
            in3 => \N__8630\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__7889\,
            in1 => \N__5911\,
            in2 => \N__7965\,
            in3 => \N__8668\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011111111"
        )
    port map (
            in0 => \N__8978\,
            in1 => \N__6859\,
            in2 => \N__7919\,
            in3 => \N__7449\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010000"
        )
    port map (
            in0 => \N__7448\,
            in1 => \N__7902\,
            in2 => \N__6877\,
            in3 => \N__8977\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5888\,
            in1 => \N__5867\,
            in2 => \_gnd_net_\,
            in3 => \N__7450\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__7451\,
            in1 => \N__7903\,
            in2 => \N__5849\,
            in3 => \N__9026\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5846\,
            in2 => \N__5840\,
            in3 => \N__5837\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8815\,
            ce => \N__8704\,
            sr => \N__9237\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5813\,
            in1 => \N__5804\,
            in2 => \_gnd_net_\,
            in3 => \N__5753\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8815\,
            ce => \N__8704\,
            sr => \N__9237\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5774\,
            in1 => \N__7898\,
            in2 => \_gnd_net_\,
            in3 => \N__8594\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6876\,
            in2 => \N__5756\,
            in3 => \N__7452\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6482\,
            in1 => \N__6449\,
            in2 => \_gnd_net_\,
            in3 => \N__6397\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_1_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6697\,
            in1 => \N__6273\,
            in2 => \N__6088\,
            in3 => \N__6612\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7897\,
            in2 => \N__6191\,
            in3 => \N__6171\,
            lcout => \U712_CHIP_RAM.N_248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__6080\,
            in1 => \N__6701\,
            in2 => \_gnd_net_\,
            in3 => \N__6616\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_0_2_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__7218\,
            in1 => \N__7088\,
            in2 => \N__7073\,
            in3 => \N__7166\,
            lcout => \U712_REG_SM.N_171\,
            ltout => \U712_REG_SM.N_171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__7112\,
            in1 => \_gnd_net_\,
            in2 => \N__5939\,
            in3 => \N__7140\,
            lcout => \U712_REG_SM.N_205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIFFTG1_2_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7220\,
            in1 => \N__7138\,
            in2 => \N__7175\,
            in3 => \N__7110\,
            lcout => OPEN,
            ltout => \U712_REG_SM.DS_EN_0_sqmuxa_0_a2_0_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7090\,
            in1 => \N__7071\,
            in2 => \N__5936\,
            in3 => \N__5932\,
            lcout => \U712_REG_SM.DS_EN_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7089\,
            in1 => \N__7219\,
            in2 => \N__7174\,
            in3 => \N__7070\,
            lcout => \U712_REG_SM.N_199\,
            ltout => \U712_REG_SM.N_199_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7111\,
            in2 => \N__6791\,
            in3 => \N__7139\,
            lcout => \U712_REG_SM.N_210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__8394\,
            in1 => \N__6787\,
            in2 => \N__6770\,
            in3 => \N__6528\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_208_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6746\,
            in3 => \N__9285\,
            lcout => \U712_CYCLE_TERM.N_208_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__6734\,
            in1 => \N__6727\,
            in2 => \_gnd_net_\,
            in3 => \N__6623\,
            lcout => \U712_CHIP_RAM.N_249\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6973\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6557\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__7109\,
            in1 => \N__7741\,
            in2 => \N__6515\,
            in3 => \N__7148\,
            lcout => \U712_REG_SM.STATE_COUNT_RNITQLC2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__7108\,
            in1 => \N__6503\,
            in2 => \_gnd_net_\,
            in3 => \N__7147\,
            lcout => \U712_REG_SM.N_174\,
            ltout => \U712_REG_SM.N_174_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIBM0G2_2_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__6961\,
            in1 => \_gnd_net_\,
            in2 => \N__6497\,
            in3 => \N__6494\,
            lcout => \U712_REG_SM.N_202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000000000"
        )
    port map (
            in0 => \N__7010\,
            in1 => \N__7033\,
            in2 => \N__6992\,
            in3 => \N__7052\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8828\,
            ce => 'H',
            sr => \N__9217\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__7034\,
            in1 => \N__6988\,
            in2 => \N__7490\,
            in3 => \N__7510\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8828\,
            ce => 'H',
            sr => \N__9217\
        );

    \U712_REG_SM.REG_TACK_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111010"
        )
    port map (
            in0 => \N__7032\,
            in1 => \N__7011\,
            in2 => \N__6977\,
            in3 => \N__6987\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8828\,
            ce => 'H',
            sr => \N__9217\
        );

    \DBR_SYNC_0_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8517\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8828\,
            ce => 'H',
            sr => \N__9217\
        );

    \U712_CHIP_RAM.CASn_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7466\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8802\,
            ce => 'H',
            sr => \N__9264\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8071\,
            in1 => \N__7453\,
            in2 => \N__8144\,
            in3 => \N__8194\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8803\,
            ce => \N__8725\,
            sr => \N__9253\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__7921\,
            in1 => \N__6914\,
            in2 => \N__7465\,
            in3 => \N__9050\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__7296\,
            in1 => \N__6872\,
            in2 => \N__6905\,
            in3 => \N__9443\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8805\,
            ce => \N__8711\,
            sr => \N__9243\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__8675\,
            in1 => \N__7297\,
            in2 => \N__6883\,
            in3 => \N__6821\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8805\,
            ce => \N__8711\,
            sr => \N__9243\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7887\,
            in2 => \_gnd_net_\,
            in3 => \N__7447\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8618\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9388\,
            ce => \N__9351\,
            sr => \N__9231\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8657\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9388\,
            ce => \N__9351\,
            sr => \N__9231\
        );

    \U712_REG_SM.C3_SYNC_0_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7252\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8813\,
            ce => 'H',
            sr => \N__9227\
        );

    \U712_REG_SM.C1_SYNC_2_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7072\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8816\,
            ce => 'H',
            sr => \N__9221\
        );

    \U712_REG_SM.C1_SYNC_0_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7207\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8816\,
            ce => 'H',
            sr => \N__9221\
        );

    \U712_REG_SM.C3_SYNC_1_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7173\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8816\,
            ce => 'H',
            sr => \N__9221\
        );

    \U712_REG_SM.C3_SYNC_2_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7141\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8816\,
            ce => 'H',
            sr => \N__9221\
        );

    \U712_REG_SM.C1_SYNC_1_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7091\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8816\,
            ce => 'H',
            sr => \N__9221\
        );

    \U712_REG_SM.REG_CYCLE_GO_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__7662\,
            in1 => \N__7578\,
            in2 => \N__7730\,
            in3 => \N__7627\,
            lcout => \U712_REG_SM.REG_CYCLE_GOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8819\,
            ce => 'H',
            sr => \N__9216\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__7580\,
            in1 => \N__7742\,
            in2 => \N__7729\,
            in3 => \N__7663\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8819\,
            ce => 'H',
            sr => \N__9216\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__7725\,
            in1 => \N__7577\,
            in2 => \_gnd_net_\,
            in3 => \N__7560\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8819\,
            ce => 'H',
            sr => \N__9216\
        );

    \U712_REG_SM.REGENn_1_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__7559\,
            in1 => \N__7677\,
            in2 => \_gnd_net_\,
            in3 => \N__7661\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8819\,
            ce => 'H',
            sr => \N__9216\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__7664\,
            in1 => \N__7536\,
            in2 => \_gnd_net_\,
            in3 => \N__7524\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8819\,
            ce => 'H',
            sr => \N__9216\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000111011"
        )
    port map (
            in0 => \N__7579\,
            in1 => \N__7649\,
            in2 => \N__7628\,
            in3 => \N__7615\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8819\,
            ce => 'H',
            sr => \N__9216\
        );

    \U712_REG_SM.DS_EN_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001010"
        )
    port map (
            in0 => \N__8227\,
            in1 => \N__7525\,
            in2 => \N__7565\,
            in3 => \N__7538\,
            lcout => \DS_ENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8819\,
            ce => 'H',
            sr => \N__9216\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111000000000"
        )
    port map (
            in0 => \N__7537\,
            in1 => \N__7488\,
            in2 => \N__7526\,
            in3 => \N__7506\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8819\,
            ce => 'H',
            sr => \N__9216\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__8518\,
            in1 => \N__9283\,
            in2 => \_gnd_net_\,
            in3 => \N__8480\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8434\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__8236\,
            in1 => \N__8324\,
            in2 => \_gnd_net_\,
            in3 => \N__8268\,
            lcout => \N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011111111"
        )
    port map (
            in0 => \N__8325\,
            in1 => \_gnd_net_\,
            in2 => \N__8275\,
            in3 => \N__8237\,
            lcout => \N_113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CRCSn_LC_13_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8198\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8801\,
            ce => 'H',
            sr => \N__9267\
        );

    \U712_CHIP_RAM.WEn_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8140\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8804\,
            ce => 'H',
            sr => \N__9266\
        );

    \U712_CHIP_RAM.RASn_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8072\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8807\,
            ce => 'H',
            sr => \N__9262\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__8009\,
            in1 => \N__7967\,
            in2 => \N__7922\,
            in3 => \N__8852\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8809\,
            ce => \N__8729\,
            sr => \N__9257\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__7966\,
            in1 => \N__7943\,
            in2 => \N__9017\,
            in3 => \N__7918\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8809\,
            ce => \N__8729\,
            sr => \N__9257\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9080\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9387\,
            ce => \N__9353\,
            sr => \N__9247\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9116\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9387\,
            ce => \N__9353\,
            sr => \N__9247\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8653\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__8922\,
            sr => \N__9238\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8617\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__8920\,
            sr => \N__9233\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9002\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__8920\,
            sr => \N__9233\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8558\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9385\,
            ce => \N__9341\,
            sr => \N__9230\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8557\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__8904\,
            sr => \N__9223\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__8519\,
            in1 => \N__9284\,
            in2 => \_gnd_net_\,
            in3 => \N__9395\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9112\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__8927\,
            sr => \N__9258\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9076\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__8927\,
            sr => \N__9258\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9431\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__8923\,
            sr => \N__9248\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9470\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__8923\,
            sr => \N__9248\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8963\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9386\,
            ce => \N__9352\,
            sr => \N__9239\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8998\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9386\,
            ce => \N__9352\,
            sr => \N__9239\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8962\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__8921\,
            sr => \N__9234\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8870\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9391\,
            ce => \N__9355\,
            sr => \N__9263\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9469\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9390\,
            ce => \N__9359\,
            sr => \N__9259\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9427\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9389\,
            ce => \N__9354\,
            sr => \N__9249\
        );
end \INTERFACE\;

module U109_CYCLE_TERMINATION (

    output TACKn

);

assign TACKn = 1'bz;

endmodule

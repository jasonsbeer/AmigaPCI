// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 9 2025 18:43:01

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U111_TOP" view "INTERFACE"

module U111_TOP (
    D_UU_AMIGA,
    D_LM_AMIGA,
    D_UM_AMIGA,
    D_LL_AMIGA,
    D_LM_040,
    D_UM_040,
    D_LL_040,
    D_UU_040,
    A_AMIGA,
    A_040,
    SIZ,
    TSn,
    RESETn,
    CLKRAMA,
    PORTSIZE,
    TEA_CPUn,
    LBENn,
    CLK40B,
    TBI_CPUn,
    TAn,
    CPUBGn,
    BUFENn,
    RnW,
    CLK80_CPU,
    BUFDIR,
    TCI_CPUn,
    TS_CPUn,
    CLKRAMB,
    CLK40A,
    DMAn,
    CLK40C,
    CLK40_IN,
    TACKn,
    BGn);

    inout [7:0] D_UU_AMIGA;
    inout [7:0] D_LM_AMIGA;
    inout [7:0] D_UM_AMIGA;
    inout [7:0] D_LL_AMIGA;
    inout [7:0] D_LM_040;
    inout [7:0] D_UM_040;
    inout [7:0] D_LL_040;
    inout [7:0] D_UU_040;
    output [1:0] A_AMIGA;
    input [1:0] A_040;
    input [1:0] SIZ;
    output TSn;
    input RESETn;
    output CLKRAMA;
    input PORTSIZE;
    output TEA_CPUn;
    input LBENn;
    output CLK40B;
    output TBI_CPUn;
    inout TAn;
    output CPUBGn;
    output BUFENn;
    input RnW;
    output CLK80_CPU;
    output BUFDIR;
    output TCI_CPUn;
    input TS_CPUn;
    output CLKRAMB;
    output CLK40A;
    output DMAn;
    output CLK40C;
    input CLK40_IN;
    inout TACKn;
    input BGn;

    wire N__8184;
    wire N__8168;
    wire N__8167;
    wire N__8166;
    wire N__8159;
    wire N__8158;
    wire N__8157;
    wire N__8150;
    wire N__8149;
    wire N__8148;
    wire N__8141;
    wire N__8140;
    wire N__8139;
    wire N__8132;
    wire N__8131;
    wire N__8130;
    wire N__8123;
    wire N__8122;
    wire N__8121;
    wire N__8114;
    wire N__8113;
    wire N__8112;
    wire N__8105;
    wire N__8104;
    wire N__8103;
    wire N__8096;
    wire N__8095;
    wire N__8094;
    wire N__8087;
    wire N__8086;
    wire N__8085;
    wire N__8078;
    wire N__8077;
    wire N__8076;
    wire N__8069;
    wire N__8068;
    wire N__8067;
    wire N__8060;
    wire N__8059;
    wire N__8058;
    wire N__8051;
    wire N__8050;
    wire N__8049;
    wire N__8042;
    wire N__8041;
    wire N__8040;
    wire N__8033;
    wire N__8032;
    wire N__8031;
    wire N__8024;
    wire N__8023;
    wire N__8022;
    wire N__8015;
    wire N__8014;
    wire N__8013;
    wire N__8006;
    wire N__8005;
    wire N__8004;
    wire N__7997;
    wire N__7996;
    wire N__7995;
    wire N__7988;
    wire N__7987;
    wire N__7986;
    wire N__7979;
    wire N__7978;
    wire N__7977;
    wire N__7970;
    wire N__7969;
    wire N__7968;
    wire N__7961;
    wire N__7960;
    wire N__7959;
    wire N__7952;
    wire N__7951;
    wire N__7950;
    wire N__7943;
    wire N__7942;
    wire N__7941;
    wire N__7934;
    wire N__7933;
    wire N__7932;
    wire N__7925;
    wire N__7924;
    wire N__7923;
    wire N__7916;
    wire N__7915;
    wire N__7914;
    wire N__7907;
    wire N__7906;
    wire N__7905;
    wire N__7898;
    wire N__7897;
    wire N__7896;
    wire N__7889;
    wire N__7888;
    wire N__7887;
    wire N__7880;
    wire N__7879;
    wire N__7878;
    wire N__7871;
    wire N__7870;
    wire N__7869;
    wire N__7862;
    wire N__7861;
    wire N__7860;
    wire N__7853;
    wire N__7852;
    wire N__7851;
    wire N__7844;
    wire N__7843;
    wire N__7842;
    wire N__7835;
    wire N__7834;
    wire N__7833;
    wire N__7826;
    wire N__7825;
    wire N__7824;
    wire N__7817;
    wire N__7816;
    wire N__7815;
    wire N__7808;
    wire N__7807;
    wire N__7806;
    wire N__7799;
    wire N__7798;
    wire N__7797;
    wire N__7790;
    wire N__7789;
    wire N__7788;
    wire N__7781;
    wire N__7780;
    wire N__7779;
    wire N__7772;
    wire N__7771;
    wire N__7770;
    wire N__7763;
    wire N__7762;
    wire N__7761;
    wire N__7754;
    wire N__7753;
    wire N__7752;
    wire N__7745;
    wire N__7744;
    wire N__7743;
    wire N__7736;
    wire N__7735;
    wire N__7734;
    wire N__7727;
    wire N__7726;
    wire N__7725;
    wire N__7718;
    wire N__7717;
    wire N__7716;
    wire N__7709;
    wire N__7708;
    wire N__7707;
    wire N__7700;
    wire N__7699;
    wire N__7698;
    wire N__7691;
    wire N__7690;
    wire N__7689;
    wire N__7682;
    wire N__7681;
    wire N__7680;
    wire N__7673;
    wire N__7672;
    wire N__7671;
    wire N__7664;
    wire N__7663;
    wire N__7662;
    wire N__7655;
    wire N__7654;
    wire N__7653;
    wire N__7646;
    wire N__7645;
    wire N__7644;
    wire N__7637;
    wire N__7636;
    wire N__7635;
    wire N__7628;
    wire N__7627;
    wire N__7626;
    wire N__7619;
    wire N__7618;
    wire N__7617;
    wire N__7610;
    wire N__7609;
    wire N__7608;
    wire N__7601;
    wire N__7600;
    wire N__7599;
    wire N__7592;
    wire N__7591;
    wire N__7590;
    wire N__7583;
    wire N__7582;
    wire N__7581;
    wire N__7574;
    wire N__7573;
    wire N__7572;
    wire N__7565;
    wire N__7564;
    wire N__7563;
    wire N__7556;
    wire N__7555;
    wire N__7554;
    wire N__7547;
    wire N__7546;
    wire N__7545;
    wire N__7538;
    wire N__7537;
    wire N__7536;
    wire N__7529;
    wire N__7528;
    wire N__7527;
    wire N__7520;
    wire N__7519;
    wire N__7518;
    wire N__7511;
    wire N__7510;
    wire N__7509;
    wire N__7502;
    wire N__7501;
    wire N__7500;
    wire N__7493;
    wire N__7492;
    wire N__7491;
    wire N__7484;
    wire N__7483;
    wire N__7482;
    wire N__7475;
    wire N__7474;
    wire N__7473;
    wire N__7466;
    wire N__7465;
    wire N__7464;
    wire N__7457;
    wire N__7456;
    wire N__7455;
    wire N__7448;
    wire N__7447;
    wire N__7446;
    wire N__7439;
    wire N__7438;
    wire N__7437;
    wire N__7430;
    wire N__7429;
    wire N__7428;
    wire N__7421;
    wire N__7420;
    wire N__7419;
    wire N__7412;
    wire N__7411;
    wire N__7410;
    wire N__7403;
    wire N__7402;
    wire N__7401;
    wire N__7394;
    wire N__7393;
    wire N__7392;
    wire N__7385;
    wire N__7384;
    wire N__7383;
    wire N__7376;
    wire N__7375;
    wire N__7374;
    wire N__7367;
    wire N__7366;
    wire N__7365;
    wire N__7358;
    wire N__7357;
    wire N__7356;
    wire N__7349;
    wire N__7348;
    wire N__7347;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7321;
    wire N__7320;
    wire N__7319;
    wire N__7316;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7302;
    wire N__7299;
    wire N__7296;
    wire N__7293;
    wire N__7290;
    wire N__7287;
    wire N__7284;
    wire N__7281;
    wire N__7278;
    wire N__7273;
    wire N__7272;
    wire N__7267;
    wire N__7264;
    wire N__7263;
    wire N__7262;
    wire N__7261;
    wire N__7260;
    wire N__7259;
    wire N__7258;
    wire N__7257;
    wire N__7254;
    wire N__7251;
    wire N__7250;
    wire N__7249;
    wire N__7248;
    wire N__7243;
    wire N__7234;
    wire N__7233;
    wire N__7232;
    wire N__7231;
    wire N__7230;
    wire N__7229;
    wire N__7228;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7216;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7200;
    wire N__7195;
    wire N__7190;
    wire N__7189;
    wire N__7188;
    wire N__7185;
    wire N__7180;
    wire N__7177;
    wire N__7170;
    wire N__7165;
    wire N__7162;
    wire N__7159;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7120;
    wire N__7119;
    wire N__7116;
    wire N__7113;
    wire N__7112;
    wire N__7109;
    wire N__7106;
    wire N__7103;
    wire N__7100;
    wire N__7095;
    wire N__7092;
    wire N__7089;
    wire N__7086;
    wire N__7083;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7044;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7036;
    wire N__7033;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7017;
    wire N__7014;
    wire N__7011;
    wire N__7006;
    wire N__7005;
    wire N__7004;
    wire N__7003;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6991;
    wire N__6982;
    wire N__6979;
    wire N__6976;
    wire N__6975;
    wire N__6974;
    wire N__6971;
    wire N__6968;
    wire N__6965;
    wire N__6960;
    wire N__6957;
    wire N__6954;
    wire N__6951;
    wire N__6948;
    wire N__6945;
    wire N__6942;
    wire N__6939;
    wire N__6936;
    wire N__6931;
    wire N__6928;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6906;
    wire N__6905;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6888;
    wire N__6885;
    wire N__6882;
    wire N__6877;
    wire N__6874;
    wire N__6871;
    wire N__6868;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6856;
    wire N__6853;
    wire N__6850;
    wire N__6847;
    wire N__6844;
    wire N__6841;
    wire N__6838;
    wire N__6837;
    wire N__6834;
    wire N__6831;
    wire N__6826;
    wire N__6825;
    wire N__6822;
    wire N__6819;
    wire N__6814;
    wire N__6811;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6799;
    wire N__6796;
    wire N__6793;
    wire N__6790;
    wire N__6787;
    wire N__6784;
    wire N__6781;
    wire N__6778;
    wire N__6775;
    wire N__6772;
    wire N__6771;
    wire N__6768;
    wire N__6765;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6755;
    wire N__6752;
    wire N__6749;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6723;
    wire N__6718;
    wire N__6715;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6694;
    wire N__6693;
    wire N__6690;
    wire N__6687;
    wire N__6684;
    wire N__6681;
    wire N__6680;
    wire N__6675;
    wire N__6672;
    wire N__6667;
    wire N__6664;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6630;
    wire N__6629;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6617;
    wire N__6612;
    wire N__6609;
    wire N__6606;
    wire N__6603;
    wire N__6600;
    wire N__6597;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6561;
    wire N__6558;
    wire N__6555;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6545;
    wire N__6540;
    wire N__6537;
    wire N__6534;
    wire N__6531;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6502;
    wire N__6499;
    wire N__6496;
    wire N__6493;
    wire N__6490;
    wire N__6487;
    wire N__6484;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6460;
    wire N__6459;
    wire N__6458;
    wire N__6455;
    wire N__6452;
    wire N__6449;
    wire N__6446;
    wire N__6443;
    wire N__6440;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6411;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6360;
    wire N__6359;
    wire N__6356;
    wire N__6353;
    wire N__6350;
    wire N__6347;
    wire N__6342;
    wire N__6339;
    wire N__6336;
    wire N__6331;
    wire N__6328;
    wire N__6325;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6303;
    wire N__6302;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6290;
    wire N__6283;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6261;
    wire N__6258;
    wire N__6253;
    wire N__6250;
    wire N__6249;
    wire N__6248;
    wire N__6247;
    wire N__6246;
    wire N__6243;
    wire N__6242;
    wire N__6241;
    wire N__6240;
    wire N__6239;
    wire N__6236;
    wire N__6233;
    wire N__6228;
    wire N__6225;
    wire N__6218;
    wire N__6215;
    wire N__6202;
    wire N__6201;
    wire N__6200;
    wire N__6199;
    wire N__6198;
    wire N__6197;
    wire N__6194;
    wire N__6193;
    wire N__6192;
    wire N__6191;
    wire N__6188;
    wire N__6183;
    wire N__6178;
    wire N__6175;
    wire N__6170;
    wire N__6167;
    wire N__6154;
    wire N__6153;
    wire N__6152;
    wire N__6149;
    wire N__6148;
    wire N__6147;
    wire N__6144;
    wire N__6141;
    wire N__6138;
    wire N__6137;
    wire N__6134;
    wire N__6131;
    wire N__6130;
    wire N__6129;
    wire N__6122;
    wire N__6117;
    wire N__6114;
    wire N__6109;
    wire N__6106;
    wire N__6103;
    wire N__6098;
    wire N__6095;
    wire N__6094;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6080;
    wire N__6075;
    wire N__6072;
    wire N__6069;
    wire N__6066;
    wire N__6063;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6045;
    wire N__6042;
    wire N__6041;
    wire N__6038;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6020;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5992;
    wire N__5989;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5977;
    wire N__5974;
    wire N__5973;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5943;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5904;
    wire N__5903;
    wire N__5900;
    wire N__5897;
    wire N__5894;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5878;
    wire N__5875;
    wire N__5872;
    wire N__5871;
    wire N__5868;
    wire N__5867;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5850;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5831;
    wire N__5828;
    wire N__5825;
    wire N__5822;
    wire N__5819;
    wire N__5814;
    wire N__5811;
    wire N__5806;
    wire N__5801;
    wire N__5796;
    wire N__5793;
    wire N__5788;
    wire N__5785;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5767;
    wire N__5766;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5754;
    wire N__5753;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5736;
    wire N__5733;
    wire N__5730;
    wire N__5725;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5704;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5692;
    wire N__5689;
    wire N__5688;
    wire N__5687;
    wire N__5686;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5673;
    wire N__5670;
    wire N__5667;
    wire N__5664;
    wire N__5661;
    wire N__5650;
    wire N__5647;
    wire N__5644;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5625;
    wire N__5622;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5554;
    wire N__5551;
    wire N__5548;
    wire N__5547;
    wire N__5544;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5478;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5457;
    wire N__5456;
    wire N__5453;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5440;
    wire N__5439;
    wire N__5430;
    wire N__5427;
    wire N__5426;
    wire N__5425;
    wire N__5424;
    wire N__5423;
    wire N__5422;
    wire N__5421;
    wire N__5420;
    wire N__5419;
    wire N__5418;
    wire N__5417;
    wire N__5416;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5385;
    wire N__5384;
    wire N__5383;
    wire N__5382;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5357;
    wire N__5354;
    wire N__5353;
    wire N__5352;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5331;
    wire N__5330;
    wire N__5323;
    wire N__5322;
    wire N__5317;
    wire N__5314;
    wire N__5313;
    wire N__5310;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5279;
    wire N__5276;
    wire N__5275;
    wire N__5274;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5264;
    wire N__5259;
    wire N__5254;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5236;
    wire N__5233;
    wire N__5230;
    wire N__5225;
    wire N__5224;
    wire N__5217;
    wire N__5214;
    wire N__5209;
    wire N__5206;
    wire N__5201;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5185;
    wire N__5182;
    wire N__5181;
    wire N__5180;
    wire N__5177;
    wire N__5176;
    wire N__5175;
    wire N__5172;
    wire N__5167;
    wire N__5162;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5146;
    wire N__5143;
    wire N__5140;
    wire N__5139;
    wire N__5138;
    wire N__5135;
    wire N__5130;
    wire N__5127;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5101;
    wire N__5098;
    wire N__5095;
    wire N__5092;
    wire N__5089;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5020;
    wire N__5017;
    wire N__5014;
    wire N__5011;
    wire N__5008;
    wire N__5005;
    wire N__5002;
    wire N__4999;
    wire N__4996;
    wire N__4993;
    wire N__4990;
    wire N__4987;
    wire N__4984;
    wire N__4981;
    wire N__4980;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4933;
    wire N__4930;
    wire N__4927;
    wire N__4924;
    wire N__4921;
    wire N__4918;
    wire N__4915;
    wire N__4912;
    wire N__4909;
    wire N__4906;
    wire N__4903;
    wire N__4900;
    wire N__4897;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4882;
    wire N__4881;
    wire N__4880;
    wire N__4879;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4871;
    wire N__4870;
    wire N__4869;
    wire N__4864;
    wire N__4861;
    wire N__4860;
    wire N__4859;
    wire N__4858;
    wire N__4857;
    wire N__4856;
    wire N__4855;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4836;
    wire N__4831;
    wire N__4830;
    wire N__4829;
    wire N__4824;
    wire N__4821;
    wire N__4820;
    wire N__4819;
    wire N__4818;
    wire N__4817;
    wire N__4816;
    wire N__4815;
    wire N__4814;
    wire N__4813;
    wire N__4812;
    wire N__4809;
    wire N__4808;
    wire N__4807;
    wire N__4800;
    wire N__4797;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4770;
    wire N__4765;
    wire N__4762;
    wire N__4761;
    wire N__4760;
    wire N__4759;
    wire N__4754;
    wire N__4751;
    wire N__4746;
    wire N__4743;
    wire N__4734;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4712;
    wire N__4709;
    wire N__4708;
    wire N__4705;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4687;
    wire N__4680;
    wire N__4677;
    wire N__4674;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4650;
    wire N__4647;
    wire N__4644;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4609;
    wire N__4606;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4573;
    wire N__4570;
    wire N__4567;
    wire N__4564;
    wire N__4561;
    wire N__4558;
    wire N__4555;
    wire N__4552;
    wire N__4549;
    wire N__4546;
    wire N__4543;
    wire N__4540;
    wire N__4537;
    wire N__4534;
    wire N__4531;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4521;
    wire N__4520;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4467;
    wire N__4462;
    wire N__4459;
    wire N__4458;
    wire N__4455;
    wire N__4454;
    wire N__4453;
    wire N__4452;
    wire N__4451;
    wire N__4450;
    wire N__4449;
    wire N__4448;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4399;
    wire N__4396;
    wire N__4393;
    wire N__4390;
    wire N__4387;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4375;
    wire N__4372;
    wire N__4369;
    wire N__4366;
    wire N__4363;
    wire N__4360;
    wire N__4357;
    wire N__4354;
    wire N__4351;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4302;
    wire N__4299;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4270;
    wire N__4267;
    wire N__4264;
    wire N__4261;
    wire N__4258;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4222;
    wire N__4219;
    wire N__4216;
    wire N__4215;
    wire N__4212;
    wire N__4209;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4197;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4122;
    wire N__4119;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4105;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4093;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4075;
    wire N__4072;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4060;
    wire N__4057;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4038;
    wire N__4035;
    wire N__4032;
    wire N__4029;
    wire N__4026;
    wire N__4021;
    wire N__4018;
    wire N__4015;
    wire N__4012;
    wire N__4009;
    wire N__4006;
    wire N__4003;
    wire N__4000;
    wire N__3997;
    wire N__3994;
    wire N__3991;
    wire N__3988;
    wire N__3985;
    wire N__3982;
    wire N__3979;
    wire N__3976;
    wire N__3973;
    wire N__3970;
    wire N__3967;
    wire N__3964;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3952;
    wire N__3949;
    wire N__3946;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3934;
    wire N__3931;
    wire N__3928;
    wire N__3925;
    wire N__3922;
    wire N__3919;
    wire N__3916;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3898;
    wire N__3897;
    wire N__3894;
    wire N__3891;
    wire N__3888;
    wire N__3885;
    wire N__3882;
    wire N__3879;
    wire N__3876;
    wire N__3873;
    wire N__3870;
    wire N__3865;
    wire N__3862;
    wire N__3859;
    wire N__3856;
    wire N__3853;
    wire N__3850;
    wire N__3847;
    wire N__3844;
    wire N__3841;
    wire N__3838;
    wire N__3835;
    wire N__3832;
    wire N__3829;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3817;
    wire N__3814;
    wire N__3811;
    wire N__3808;
    wire N__3805;
    wire N__3802;
    wire N__3799;
    wire N__3796;
    wire N__3793;
    wire N__3792;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3760;
    wire N__3757;
    wire N__3754;
    wire N__3751;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3736;
    wire N__3733;
    wire N__3730;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3717;
    wire N__3714;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3694;
    wire N__3691;
    wire N__3688;
    wire N__3685;
    wire N__3682;
    wire N__3679;
    wire N__3676;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3664;
    wire N__3661;
    wire N__3658;
    wire N__3655;
    wire N__3652;
    wire N__3649;
    wire N__3646;
    wire N__3643;
    wire N__3640;
    wire N__3637;
    wire N__3636;
    wire N__3633;
    wire N__3630;
    wire N__3627;
    wire N__3624;
    wire N__3621;
    wire N__3618;
    wire N__3615;
    wire N__3610;
    wire N__3607;
    wire N__3604;
    wire N__3601;
    wire N__3598;
    wire N__3595;
    wire N__3592;
    wire N__3589;
    wire N__3586;
    wire N__3583;
    wire N__3580;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3568;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3550;
    wire N__3547;
    wire N__3544;
    wire N__3541;
    wire N__3538;
    wire N__3535;
    wire N__3532;
    wire N__3529;
    wire N__3526;
    wire N__3523;
    wire N__3520;
    wire N__3517;
    wire N__3514;
    wire N__3511;
    wire N__3508;
    wire N__3505;
    wire N__3502;
    wire N__3499;
    wire N__3496;
    wire N__3493;
    wire N__3490;
    wire N__3487;
    wire N__3484;
    wire N__3481;
    wire N__3478;
    wire N__3475;
    wire N__3472;
    wire N__3469;
    wire N__3466;
    wire N__3463;
    wire N__3460;
    wire N__3457;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3445;
    wire N__3442;
    wire N__3439;
    wire N__3436;
    wire N__3433;
    wire N__3430;
    wire N__3427;
    wire N__3426;
    wire N__3423;
    wire N__3420;
    wire N__3417;
    wire N__3414;
    wire N__3411;
    wire N__3408;
    wire N__3405;
    wire N__3402;
    wire N__3399;
    wire N__3396;
    wire N__3391;
    wire N__3388;
    wire N__3385;
    wire N__3382;
    wire N__3379;
    wire N__3376;
    wire N__3373;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3361;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3337;
    wire N__3334;
    wire N__3331;
    wire N__3328;
    wire N__3325;
    wire N__3322;
    wire N__3319;
    wire N__3316;
    wire N__3313;
    wire N__3310;
    wire N__3307;
    wire N__3304;
    wire N__3301;
    wire N__3298;
    wire N__3295;
    wire N__3292;
    wire N__3289;
    wire N__3286;
    wire N__3283;
    wire N__3280;
    wire N__3277;
    wire N__3274;
    wire N__3271;
    wire N__3268;
    wire N__3265;
    wire N__3262;
    wire N__3259;
    wire N__3256;
    wire N__3253;
    wire N__3250;
    wire N__3247;
    wire N__3244;
    wire N__3241;
    wire N__3238;
    wire N__3235;
    wire N__3232;
    wire N__3229;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3190;
    wire N__3187;
    wire N__3184;
    wire N__3181;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3171;
    wire N__3168;
    wire N__3165;
    wire N__3162;
    wire N__3159;
    wire N__3156;
    wire N__3153;
    wire N__3150;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3121;
    wire N__3118;
    wire N__3117;
    wire N__3114;
    wire N__3111;
    wire N__3108;
    wire N__3105;
    wire N__3102;
    wire N__3099;
    wire N__3096;
    wire N__3093;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3070;
    wire N__3067;
    wire N__3064;
    wire N__3061;
    wire N__3058;
    wire N__3055;
    wire N__3052;
    wire N__3049;
    wire N__3046;
    wire N__3043;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3031;
    wire N__3028;
    wire N__3025;
    wire N__3022;
    wire N__3019;
    wire N__3016;
    wire N__3013;
    wire N__3010;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__2998;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2980;
    wire N__2979;
    wire N__2976;
    wire N__2973;
    wire N__2970;
    wire N__2967;
    wire N__2964;
    wire N__2961;
    wire N__2958;
    wire N__2955;
    wire N__2952;
    wire N__2949;
    wire N__2946;
    wire N__2943;
    wire N__2938;
    wire N__2935;
    wire N__2932;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2920;
    wire N__2917;
    wire N__2914;
    wire N__2911;
    wire N__2908;
    wire N__2905;
    wire N__2902;
    wire N__2899;
    wire N__2896;
    wire N__2893;
    wire N__2892;
    wire N__2891;
    wire N__2888;
    wire N__2883;
    wire N__2882;
    wire N__2879;
    wire N__2876;
    wire N__2873;
    wire N__2870;
    wire N__2867;
    wire N__2864;
    wire N__2859;
    wire N__2856;
    wire N__2853;
    wire N__2850;
    wire N__2847;
    wire N__2842;
    wire N__2839;
    wire N__2836;
    wire N__2833;
    wire N__2830;
    wire N__2827;
    wire N__2824;
    wire N__2821;
    wire N__2818;
    wire N__2815;
    wire N__2814;
    wire N__2811;
    wire N__2808;
    wire N__2805;
    wire N__2802;
    wire N__2799;
    wire N__2796;
    wire N__2791;
    wire N__2788;
    wire N__2785;
    wire N__2782;
    wire N__2779;
    wire N__2776;
    wire N__2773;
    wire N__2770;
    wire N__2767;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2755;
    wire N__2752;
    wire N__2749;
    wire N__2746;
    wire N__2745;
    wire N__2742;
    wire N__2739;
    wire N__2736;
    wire N__2733;
    wire N__2730;
    wire N__2727;
    wire N__2724;
    wire N__2721;
    wire N__2718;
    wire N__2715;
    wire N__2712;
    wire N__2709;
    wire N__2706;
    wire N__2701;
    wire N__2698;
    wire N__2695;
    wire N__2692;
    wire N__2689;
    wire N__2686;
    wire N__2683;
    wire N__2680;
    wire N__2677;
    wire N__2674;
    wire N__2671;
    wire N__2668;
    wire N__2665;
    wire N__2662;
    wire N__2659;
    wire N__2656;
    wire N__2653;
    wire N__2650;
    wire N__2647;
    wire N__2644;
    wire N__2641;
    wire N__2638;
    wire N__2635;
    wire N__2632;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2620;
    wire N__2617;
    wire N__2614;
    wire N__2611;
    wire N__2608;
    wire N__2605;
    wire N__2602;
    wire N__2599;
    wire N__2596;
    wire N__2593;
    wire N__2590;
    wire N__2587;
    wire N__2584;
    wire N__2581;
    wire N__2578;
    wire N__2575;
    wire N__2574;
    wire N__2573;
    wire N__2572;
    wire N__2569;
    wire N__2566;
    wire N__2563;
    wire N__2560;
    wire N__2559;
    wire N__2558;
    wire N__2549;
    wire N__2546;
    wire N__2543;
    wire N__2542;
    wire N__2535;
    wire N__2532;
    wire N__2531;
    wire N__2530;
    wire N__2529;
    wire N__2526;
    wire N__2523;
    wire N__2520;
    wire N__2517;
    wire N__2514;
    wire N__2513;
    wire N__2512;
    wire N__2511;
    wire N__2510;
    wire N__2509;
    wire N__2508;
    wire N__2507;
    wire N__2496;
    wire N__2493;
    wire N__2490;
    wire N__2489;
    wire N__2488;
    wire N__2485;
    wire N__2482;
    wire N__2479;
    wire N__2476;
    wire N__2475;
    wire N__2474;
    wire N__2473;
    wire N__2472;
    wire N__2469;
    wire N__2468;
    wire N__2467;
    wire N__2460;
    wire N__2457;
    wire N__2454;
    wire N__2453;
    wire N__2452;
    wire N__2451;
    wire N__2450;
    wire N__2449;
    wire N__2440;
    wire N__2437;
    wire N__2434;
    wire N__2431;
    wire N__2428;
    wire N__2425;
    wire N__2422;
    wire N__2419;
    wire N__2412;
    wire N__2409;
    wire N__2406;
    wire N__2403;
    wire N__2400;
    wire N__2397;
    wire N__2396;
    wire N__2395;
    wire N__2386;
    wire N__2371;
    wire N__2366;
    wire N__2363;
    wire N__2360;
    wire N__2357;
    wire N__2354;
    wire N__2351;
    wire N__2348;
    wire N__2345;
    wire N__2340;
    wire N__2337;
    wire N__2334;
    wire N__2331;
    wire N__2326;
    wire N__2323;
    wire N__2320;
    wire VCCG0;
    wire GNDG0;
    wire TAn_in;
    wire A_040_c_1;
    wire A_040_c_0;
    wire A_AMIGA_c_0;
    wire RnW_c_i;
    wire D_LL_040_in_2;
    wire D_UM_040_in_2;
    wire un1_D_UM_040_2;
    wire D_LM_AMIGA_in_5;
    wire un1_D_LM_AMIGA_5;
    wire D_LM_AMIGA_in_6;
    wire un1_D_LM_AMIGA_6;
    wire D_LL_040_in_3;
    wire D_UM_040_in_3;
    wire un1_D_UM_040_3;
    wire CONSTANT_ONE_NET;
    wire D_UU_040_in_6;
    wire D_LM_040_in_6;
    wire un1_D_UU_040_6;
    wire D_UU_040_in_0;
    wire D_LM_040_in_0;
    wire un1_D_UU_040_0;
    wire D_LM_AMIGA_in_3;
    wire un1_D_LM_AMIGA_3;
    wire D_LM_AMIGA_in_2;
    wire un1_D_LM_AMIGA_2;
    wire D_LL_040_in_7;
    wire D_UM_040_in_7;
    wire un1_D_UM_040_7;
    wire D_LL_AMIGA_in_0;
    wire un1_D_LL_AMIGA_0;
    wire LBENn_c_i_0;
    wire TSn_c;
    wire \INVU111_CYCLE_SM.TSnC_net ;
    wire D_LL_AMIGA_in_5;
    wire un1_D_LL_AMIGA_5;
    wire D_LM_AMIGA_in_4;
    wire un1_D_LM_AMIGA_4;
    wire D_UM_040_in_6;
    wire D_LL_040_in_6;
    wire un1_D_UM_040_6;
    wire D_LL_040_in_1;
    wire D_UM_040_in_1;
    wire un1_D_UM_040_1;
    wire LBENn_c_i;
    wire D_LM_040_in_1;
    wire D_UU_040_in_1;
    wire un1_D_UU_040_1;
    wire D_LM_040_in_4;
    wire D_UU_040_in_4;
    wire un1_D_UU_040_4;
    wire D_UU_040_in_2;
    wire D_LM_040_in_2;
    wire un1_D_UU_040_2;
    wire D_LL_AMIGA_in_2;
    wire un1_D_LL_AMIGA_2;
    wire D_LL_AMIGA_in_4;
    wire un1_D_LL_AMIGA_4;
    wire D_LL_AMIGA_in_6;
    wire un1_D_LL_AMIGA_6;
    wire D_LM_AMIGA_in_0;
    wire un1_D_LM_AMIGA_0;
    wire D_LL_AMIGA_in_7;
    wire un1_D_LL_AMIGA_7;
    wire D_LL_040_in_0;
    wire D_UM_040_in_0;
    wire un1_D_UM_040_0;
    wire D_UM_040_in_4;
    wire D_LL_040_in_4;
    wire un1_D_UM_040_4;
    wire D_LM_040_in_5;
    wire D_UU_040_in_5;
    wire un1_D_UU_040_5;
    wire D_LM_040_in_7;
    wire D_UU_040_in_7;
    wire un1_D_UU_040_7;
    wire D_LL_AMIGA_in_3;
    wire un1_D_LL_AMIGA_3;
    wire D_LL_AMIGA_in_1;
    wire un1_D_LL_AMIGA_1;
    wire A_AMIGA_c_1;
    wire D_LM_AMIGA_in_1;
    wire \U111_CYCLE_SM.FLIP_cascade_ ;
    wire un1_D_LM_AMIGA_1;
    wire GB_BUFFER_CLK40_THRU_CO;
    wire CLK80;
    wire GB_BUFFER_CLK80_THRU_CO;
    wire \U111_CYCLE_SM.A_OUT_0_cascade_ ;
    wire \U111_CYCLE_SM.A_OUTZ0 ;
    wire \U111_CYCLE_SM.N_75_0_cascade_ ;
    wire \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net ;
    wire \U111_CYCLE_SM.TS_ENZ0 ;
    wire \U111_CYCLE_SM.un3_LW_CYCLE_START ;
    wire \INVU111_CYCLE_SM.TA_ENC_net ;
    wire \U111_CYCLE_SM.RESETn_c_i ;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire PORTSIZE_c;
    wire \U111_CYCLE_SM.LW_TRANS_0 ;
    wire D_LM_AMIGA_in_7;
    wire un1_D_LM_AMIGA_7;
    wire D_LL_040_in_5;
    wire D_UM_040_in_5;
    wire un1_D_UM_040_5;
    wire D_UU_040_in_3;
    wire \U111_CYCLE_SM.FLIP ;
    wire D_LM_040_in_3;
    wire un1_D_UU_040_3;
    wire U111_CYCLE_SM_TBI_CPUn_0_i;
    wire \U111_CYCLE_SM.TS_EN_5 ;
    wire BGn_c;
    wire CPU_READ_EN_i;
    wire \INVU111_CYCLE_SM.CYCLE_STATE_1C_net ;
    wire \U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0_cascade_ ;
    wire \U111_CYCLE_SM.LW_CYCLE_STARTZ0 ;
    wire \U111_CYCLE_SM.N_97_cascade_ ;
    wire \INVU111_CYCLE_SM.LW_CYCLEC_net ;
    wire \U111_CYCLE_SM.LW_CYCLE_0 ;
    wire \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net ;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ;
    wire D_UU_AMIGA_in_1;
    wire un1_D_UU_AMIGA_1;
    wire \U111_CYCLE_SM.TA_ENZ0 ;
    wire LBENn_c;
    wire TAn_1_i;
    wire D_UM_AMIGA_in_1;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ;
    wire un1_D_UM_AMIGA_1;
    wire TS_CPUn_c;
    wire CLK40;
    wire \U111_CYCLE_SM.TS_EN_2_0 ;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ;
    wire D_UU_AMIGA_in_7;
    wire un1_D_UU_AMIGA_7;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ;
    wire D_UU_AMIGA_in_2;
    wire un1_D_UU_AMIGA_2;
    wire un1_D_UM_AMIGA_0;
    wire un1_D_UM_AMIGA_2;
    wire un1_D_UM_AMIGA_6;
    wire D_UM_AMIGA_in_0;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ;
    wire D_UM_AMIGA_in_6;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ;
    wire D_UM_AMIGA_in_2;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net ;
    wire TACKn_in;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ;
    wire RESETn_c;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_ ;
    wire RnW_c;
    wire \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa ;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ;
    wire D_UM_AMIGA_in_5;
    wire un1_D_UM_AMIGA_5;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ;
    wire D_UU_AMIGA_in_3;
    wire un1_D_UU_AMIGA_3;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ;
    wire D_UU_AMIGA_in_4;
    wire un1_D_UU_AMIGA_4;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ;
    wire D_UU_AMIGA_in_6;
    wire un1_D_UU_AMIGA_6;
    wire D_UM_AMIGA_in_3;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ;
    wire un1_D_UM_AMIGA_3;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net ;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ;
    wire \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0 ;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ;
    wire D_UM_AMIGA_in_7;
    wire un1_D_UM_AMIGA_7;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ;
    wire D_UU_AMIGA_in_0;
    wire un1_D_UU_AMIGA_0;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ;
    wire D_UU_AMIGA_in_5;
    wire un1_D_UU_AMIGA_5;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ;
    wire D_UM_AMIGA_in_4;
    wire \U111_CYCLE_SM.LW_CYCLEZ0 ;
    wire un1_D_UM_AMIGA_4;
    wire _gnd_net_;

    defparam pll_pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll_pll.TEST_MODE=1'b0;
    defparam pll_pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll_pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll_pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll_pll.FILTER_RANGE=3'b011;
    defparam pll_pll.FEEDBACK_PATH="SIMPLE";
    defparam pll_pll.FDA_RELATIVE=4'b0000;
    defparam pll_pll.FDA_FEEDBACK=4'b0000;
    defparam pll_pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll_pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll_pll.DIVR=4'b0000;
    defparam pll_pll.DIVQ=3'b011;
    defparam pll_pll.DIVF=7'b0001111;
    defparam pll_pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40_2F pll_pll (
            .SCLK(),
            .PLLOUTGLOBALA(CLK80),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALB(CLK40),
            .SDI(),
            .PLLOUTCOREA(),
            .BYPASS(),
            .RESETB(N__2891),
            .PLLOUTCOREB(),
            .LOCK(),
            .SDO(),
            .EXTFEEDBACK(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__8184));
    IO_PAD pll_iopad (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__8184),
            .PACKAGEPIN(CLK40_IN));
    IO_PAD LBENn_ibuf_iopad (
            .OE(N__8168),
            .DIN(N__8167),
            .DOUT(N__8166),
            .PACKAGEPIN(LBENn));
    defparam LBENn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam LBENn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO LBENn_ibuf_preio (
            .PADOEN(N__8168),
            .PADOUT(N__8167),
            .PADIN(N__8166),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(LBENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_3_iopad (
            .OE(N__8159),
            .DIN(N__8158),
            .DOUT(N__8157),
            .PACKAGEPIN(D_UM_040[3]));
    defparam D_UM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_3_preio (
            .PADOEN(N__8159),
            .PADOUT(N__8158),
            .PADIN(N__8157),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5417),
            .DIN0(D_UM_040_in_3),
            .DOUT0(N__7066),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TAn_iobuf_iopad.PULLUP=1'b1;
    IO_PAD TAn_iobuf_iopad (
            .OE(N__8150),
            .DIN(N__8149),
            .DOUT(N__8148),
            .PACKAGEPIN(TAn));
    defparam TAn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TAn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TAn_iobuf_preio (
            .PADOEN(N__8150),
            .PADOUT(N__8149),
            .PADIN(N__8148),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5788),
            .DIN0(TAn_in),
            .DOUT0(N__6316),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_1_iopad (
            .OE(N__8141),
            .DIN(N__8140),
            .DOUT(N__8139),
            .PACKAGEPIN(D_LL_AMIGA[1]));
    defparam D_LL_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_1_preio (
            .PADOEN(N__8141),
            .PADOUT(N__8140),
            .PADIN(N__8139),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2572),
            .DIN0(D_LL_AMIGA_in_1),
            .DOUT0(N__3898),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_5_iopad (
            .OE(N__8132),
            .DIN(N__8131),
            .DOUT(N__8130),
            .PACKAGEPIN(D_UU_AMIGA[5]));
    defparam D_UU_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_5_preio (
            .PADOEN(N__8132),
            .PADOUT(N__8131),
            .PADIN(N__8130),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2396),
            .DIN0(D_UU_AMIGA_in_5),
            .DOUT0(N__4084),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_6_iopad (
            .OE(N__8123),
            .DIN(N__8122),
            .DOUT(N__8121),
            .PACKAGEPIN(D_UU_040[6]));
    defparam D_UU_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_6_preio (
            .PADOEN(N__8123),
            .PADOUT(N__8122),
            .PADIN(N__8121),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5385),
            .DIN0(D_UU_040_in_6),
            .DOUT0(N__6520),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam CPUBGn_obuf_iopad.PULLUP=1'b1;
    IO_PAD CPUBGn_obuf_iopad (
            .OE(N__8114),
            .DIN(N__8113),
            .DOUT(N__8112),
            .PACKAGEPIN(CPUBGn));
    defparam CPUBGn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUBGn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CPUBGn_obuf_preio (
            .PADOEN(N__8114),
            .PADOUT(N__8113),
            .PADIN(N__8112),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_7_iopad (
            .OE(N__8105),
            .DIN(N__8104),
            .DOUT(N__8103),
            .PACKAGEPIN(D_LL_040[7]));
    defparam D_LL_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_7_preio (
            .PADOEN(N__8105),
            .PADOUT(N__8104),
            .PADIN(N__8103),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5423),
            .DIN0(D_LL_040_in_7),
            .DOUT0(N__4336),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_4_iopad (
            .OE(N__8096),
            .DIN(N__8095),
            .DOUT(N__8094),
            .PACKAGEPIN(D_LL_AMIGA[4]));
    defparam D_LL_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_4_preio (
            .PADOEN(N__8096),
            .PADOUT(N__8095),
            .PADIN(N__8094),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2449),
            .DIN0(D_LL_AMIGA_in_4),
            .DOUT0(N__4215),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_3_iopad (
            .OE(N__8087),
            .DIN(N__8086),
            .DOUT(N__8085),
            .PACKAGEPIN(D_UM_AMIGA[3]));
    defparam D_UM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_3_preio (
            .PADOEN(N__8087),
            .PADOUT(N__8086),
            .PADIN(N__8085),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2468),
            .DIN0(D_UM_AMIGA_in_3),
            .DOUT0(N__2917),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_3_iopad (
            .OE(N__8078),
            .DIN(N__8077),
            .DOUT(N__8076),
            .PACKAGEPIN(D_UU_040[3]));
    defparam D_UU_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_3_preio (
            .PADOEN(N__8078),
            .PADOUT(N__8077),
            .PADIN(N__8076),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5419),
            .DIN0(D_UU_040_in_3),
            .DOUT0(N__6655),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TEA_CPUn_obuf_iopad.PULLUP=1'b1;
    IO_PAD TEA_CPUn_obuf_iopad (
            .OE(N__8069),
            .DIN(N__8068),
            .DOUT(N__8067),
            .PACKAGEPIN(TEA_CPUn));
    defparam TEA_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TEA_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TEA_CPUn_obuf_preio (
            .PADOEN(N__8069),
            .PADOUT(N__8068),
            .PADIN(N__8067),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2892),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_1_iopad (
            .OE(N__8060),
            .DIN(N__8059),
            .DOUT(N__8058),
            .PACKAGEPIN(A_040[1]));
    defparam A_040_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_1_preio (
            .PADOEN(N__8060),
            .PADOUT(N__8059),
            .PADIN(N__8058),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_3_iopad (
            .OE(N__8051),
            .DIN(N__8050),
            .DOUT(N__8049),
            .PACKAGEPIN(D_LM_AMIGA[3]));
    defparam D_LM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_3_preio (
            .PADOEN(N__8051),
            .PADOUT(N__8050),
            .PADIN(N__8049),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2531),
            .DIN0(D_LM_AMIGA_in_3),
            .DOUT0(N__4657),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_0_iopad (
            .OE(N__8042),
            .DIN(N__8041),
            .DOUT(N__8040),
            .PACKAGEPIN(D_LM_040[0]));
    defparam D_LM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_0_preio (
            .PADOEN(N__8042),
            .PADOUT(N__8041),
            .PADIN(N__8040),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5424),
            .DIN0(D_LM_040_in_0),
            .DOUT0(N__4372),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_6_iopad (
            .OE(N__8033),
            .DIN(N__8032),
            .DOUT(N__8031),
            .PACKAGEPIN(D_UM_AMIGA[6]));
    defparam D_UM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_6_preio (
            .PADOEN(N__8033),
            .PADOUT(N__8032),
            .PADIN(N__8031),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2395),
            .DIN0(D_UM_AMIGA_in_6),
            .DOUT0(N__3142),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_4_iopad (
            .OE(N__8024),
            .DIN(N__8023),
            .DOUT(N__8022),
            .PACKAGEPIN(D_LM_AMIGA[4]));
    defparam D_LM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_4_preio (
            .PADOEN(N__8024),
            .PADOUT(N__8023),
            .PADIN(N__8022),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2512),
            .DIN0(D_LM_AMIGA_in_4),
            .DOUT0(N__3727),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_1_iopad (
            .OE(N__8015),
            .DIN(N__8014),
            .DOUT(N__8013),
            .PACKAGEPIN(A_AMIGA[1]));
    defparam A_AMIGA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_1_preio (
            .PADOEN(N__8015),
            .PADOUT(N__8014),
            .PADIN(N__8013),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3915),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_7_iopad (
            .OE(N__8006),
            .DIN(N__8005),
            .DOUT(N__8004),
            .PACKAGEPIN(D_LM_040[7]));
    defparam D_LM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_7_preio (
            .PADOEN(N__8006),
            .PADOUT(N__8005),
            .PADIN(N__8004),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5322),
            .DIN0(D_LM_040_in_7),
            .DOUT0(N__5002),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_4_iopad (
            .OE(N__7997),
            .DIN(N__7996),
            .DOUT(N__7995),
            .PACKAGEPIN(D_UM_040[4]));
    defparam D_UM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_4_preio (
            .PADOEN(N__7997),
            .PADOUT(N__7996),
            .PADIN(N__7995),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5420),
            .DIN0(D_UM_040_in_4),
            .DOUT0(N__7144),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_obuf_iopad (
            .OE(N__7988),
            .DIN(N__7987),
            .DOUT(N__7986),
            .PACKAGEPIN(CLK40B));
    defparam CLK40B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_obuf_preio (
            .PADOEN(N__7988),
            .PADOUT(N__7987),
            .PADIN(N__7986),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4521),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_0_iopad (
            .OE(N__7979),
            .DIN(N__7978),
            .DOUT(N__7977),
            .PACKAGEPIN(D_UU_AMIGA[0]));
    defparam D_UU_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_0_preio (
            .PADOEN(N__7979),
            .PADOUT(N__7978),
            .PADIN(N__7977),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2475),
            .DIN0(D_UU_AMIGA_in_0),
            .DOUT0(N__2698),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_1_iopad (
            .OE(N__7970),
            .DIN(N__7969),
            .DOUT(N__7968),
            .PACKAGEPIN(D_UM_040[1]));
    defparam D_UM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_1_preio (
            .PADOEN(N__7970),
            .PADOUT(N__7969),
            .PADIN(N__7968),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5352),
            .DIN0(D_UM_040_in_1),
            .DOUT0(N__5719),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_4_iopad (
            .OE(N__7961),
            .DIN(N__7960),
            .DOUT(N__7959),
            .PACKAGEPIN(D_LL_040[4]));
    defparam D_LL_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_4_preio (
            .PADOEN(N__7961),
            .PADOUT(N__7960),
            .PADIN(N__7959),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5461),
            .DIN0(D_LL_040_in_4),
            .DOUT0(N__3538),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_7_iopad (
            .OE(N__7952),
            .DIN(N__7951),
            .DOUT(N__7950),
            .PACKAGEPIN(D_LL_AMIGA[7]));
    defparam D_LL_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_7_preio (
            .PADOEN(N__7952),
            .PADOUT(N__7951),
            .PADIN(N__7950),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2450),
            .DIN0(D_LL_AMIGA_in_7),
            .DOUT0(N__3430),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_7_iopad (
            .OE(N__7943),
            .DIN(N__7942),
            .DOUT(N__7941),
            .PACKAGEPIN(D_UU_AMIGA[7]));
    defparam D_UU_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_7_preio (
            .PADOEN(N__7943),
            .PADOUT(N__7942),
            .PADIN(N__7941),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2509),
            .DIN0(D_UU_AMIGA_in_7),
            .DOUT0(N__4003),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFDIR_obuf_iopad (
            .OE(N__7934),
            .DIN(N__7933),
            .DOUT(N__7932),
            .PACKAGEPIN(BUFDIR));
    defparam BUFDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFDIR_obuf_preio (
            .PADOEN(N__7934),
            .PADOUT(N__7933),
            .PADIN(N__7932),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6052),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_5_iopad (
            .OE(N__7925),
            .DIN(N__7924),
            .DOUT(N__7923),
            .PACKAGEPIN(D_LM_AMIGA[5]));
    defparam D_LM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_5_preio (
            .PADOEN(N__7925),
            .PADOUT(N__7924),
            .PADIN(N__7923),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2488),
            .DIN0(D_LM_AMIGA_in_5),
            .DOUT0(N__4153),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_4_iopad (
            .OE(N__7916),
            .DIN(N__7915),
            .DOUT(N__7914),
            .PACKAGEPIN(D_UU_040[4]));
    defparam D_UU_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_4_preio (
            .PADOEN(N__7916),
            .PADOUT(N__7915),
            .PADIN(N__7914),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5381),
            .DIN0(D_UU_040_in_4),
            .DOUT0(N__6592),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SIZ_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__7907),
            .DIN(N__7906),
            .DOUT(N__7905),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__7907),
            .PADOUT(N__7906),
            .PADIN(N__7905),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_6_iopad (
            .OE(N__7898),
            .DIN(N__7897),
            .DOUT(N__7896),
            .PACKAGEPIN(D_LM_040[6]));
    defparam D_LM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_6_preio (
            .PADOEN(N__7898),
            .PADOUT(N__7897),
            .PADIN(N__7896),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5264),
            .DIN0(D_LM_040_in_6),
            .DOUT0(N__2995),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_5_iopad (
            .OE(N__7889),
            .DIN(N__7888),
            .DOUT(N__7887),
            .PACKAGEPIN(D_UM_040[5]));
    defparam D_UM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_5_preio (
            .PADOEN(N__7889),
            .PADOUT(N__7888),
            .PADIN(N__7887),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5274),
            .DIN0(D_UM_040_in_5),
            .DOUT0(N__6718),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TS_CPUn_ibuf_iopad (
            .OE(N__7880),
            .DIN(N__7879),
            .DOUT(N__7878),
            .PACKAGEPIN(TS_CPUn));
    defparam TS_CPUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TS_CPUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TS_CPUn_ibuf_preio (
            .PADOEN(N__7880),
            .PADOUT(N__7879),
            .PADIN(N__7878),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TS_CPUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_1_iopad (
            .OE(N__7871),
            .DIN(N__7870),
            .DOUT(N__7869),
            .PACKAGEPIN(D_LL_040[1]));
    defparam D_LL_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_1_preio (
            .PADOEN(N__7871),
            .PADOUT(N__7870),
            .PADIN(N__7869),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5452),
            .DIN0(D_LL_040_in_1),
            .DOUT0(N__3934),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_3_iopad (
            .OE(N__7862),
            .DIN(N__7861),
            .DOUT(N__7860),
            .PACKAGEPIN(D_LL_AMIGA[3]));
    defparam D_LL_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_3_preio (
            .PADOEN(N__7862),
            .PADOUT(N__7861),
            .PADIN(N__7860),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2573),
            .DIN0(D_LL_AMIGA_in_3),
            .DOUT0(N__2979),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_5_iopad (
            .OE(N__7853),
            .DIN(N__7852),
            .DOUT(N__7851),
            .PACKAGEPIN(D_UM_AMIGA[5]));
    defparam D_UM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_5_preio (
            .PADOEN(N__7853),
            .PADOUT(N__7852),
            .PADIN(N__7851),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2508),
            .DIN0(D_UM_AMIGA_in_5),
            .DOUT0(N__4915),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_1_iopad (
            .OE(N__7844),
            .DIN(N__7843),
            .DOUT(N__7842),
            .PACKAGEPIN(D_UU_040[1]));
    defparam D_UU_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_1_preio (
            .PADOEN(N__7844),
            .PADOUT(N__7843),
            .PADIN(N__7842),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5418),
            .DIN0(D_UU_040_in_1),
            .DOUT0(N__5932),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_3_iopad (
            .OE(N__7835),
            .DIN(N__7834),
            .DOUT(N__7833),
            .PACKAGEPIN(D_UU_AMIGA[3]));
    defparam D_UU_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_3_preio (
            .PADOEN(N__7835),
            .PADOUT(N__7834),
            .PADIN(N__7833),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2511),
            .DIN0(D_UU_AMIGA_in_3),
            .DOUT0(N__4609),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_1_iopad (
            .OE(N__7826),
            .DIN(N__7825),
            .DOUT(N__7824),
            .PACKAGEPIN(D_LM_AMIGA[1]));
    defparam D_LM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_1_preio (
            .PADOEN(N__7826),
            .PADOUT(N__7825),
            .PADIN(N__7824),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2542),
            .DIN0(D_LM_AMIGA_in_1),
            .DOUT0(N__3799),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_2_iopad (
            .OE(N__7817),
            .DIN(N__7816),
            .DOUT(N__7815),
            .PACKAGEPIN(D_LM_040[2]));
    defparam D_LM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_2_preio (
            .PADOEN(N__7817),
            .PADOUT(N__7816),
            .PADIN(N__7815),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5422),
            .DIN0(D_LM_040_in_2),
            .DOUT0(N__3445),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_5_iopad (
            .OE(N__7808),
            .DIN(N__7807),
            .DOUT(N__7806),
            .PACKAGEPIN(D_LL_040[5]));
    defparam D_LL_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_5_preio (
            .PADOEN(N__7808),
            .PADOUT(N__7807),
            .PADIN(N__7806),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5425),
            .DIN0(D_LL_040_in_5),
            .DOUT0(N__3262),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_6_iopad (
            .OE(N__7799),
            .DIN(N__7798),
            .DOUT(N__7797),
            .PACKAGEPIN(D_LL_AMIGA[6]));
    defparam D_LL_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_6_preio (
            .PADOEN(N__7799),
            .PADOUT(N__7798),
            .PADIN(N__7797),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2558),
            .DIN0(D_LL_AMIGA_in_6),
            .DOUT0(N__3187),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_6_iopad (
            .OE(N__7790),
            .DIN(N__7789),
            .DOUT(N__7788),
            .PACKAGEPIN(D_UU_AMIGA[6]));
    defparam D_UU_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_6_preio (
            .PADOEN(N__7790),
            .PADOUT(N__7789),
            .PADIN(N__7788),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2510),
            .DIN0(D_UU_AMIGA_in_6),
            .DOUT0(N__2785),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_1_iopad (
            .OE(N__7781),
            .DIN(N__7780),
            .DOUT(N__7779),
            .PACKAGEPIN(D_UM_AMIGA[1]));
    defparam D_UM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_1_preio (
            .PADOEN(N__7781),
            .PADOUT(N__7780),
            .PADIN(N__7779),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2489),
            .DIN0(D_UM_AMIGA_in_1),
            .DOUT0(N__3838),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_5_iopad (
            .OE(N__7772),
            .DIN(N__7771),
            .DOUT(N__7770),
            .PACKAGEPIN(D_UU_040[5]));
    defparam D_UU_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_5_preio (
            .PADOEN(N__7772),
            .PADOUT(N__7771),
            .PADIN(N__7770),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5275),
            .DIN0(D_UU_040_in_5),
            .DOUT0(N__6799),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_iobuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__7763),
            .DIN(N__7762),
            .DOUT(N__7761),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__7763),
            .PADOUT(N__7762),
            .PADIN(N__7761),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3301),
            .DIN0(TACKn_in),
            .DOUT0(N__2644),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMA_obuf_iopad (
            .OE(N__7754),
            .DIN(N__7753),
            .DOUT(N__7752),
            .PACKAGEPIN(CLKRAMA));
    defparam CLKRAMA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMA_obuf_preio (
            .PADOEN(N__7754),
            .PADOUT(N__7753),
            .PADIN(N__7752),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4525),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_2_iopad (
            .OE(N__7745),
            .DIN(N__7744),
            .DOUT(N__7743),
            .PACKAGEPIN(D_UM_040[2]));
    defparam D_UM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_2_preio (
            .PADOEN(N__7745),
            .PADOUT(N__7744),
            .PADIN(N__7743),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5313),
            .DIN0(D_UM_040_in_2),
            .DOUT0(N__6499),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_2_iopad (
            .OE(N__7736),
            .DIN(N__7735),
            .DOUT(N__7734),
            .PACKAGEPIN(D_LL_040[2]));
    defparam D_LL_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_2_preio (
            .PADOEN(N__7736),
            .PADOUT(N__7735),
            .PADIN(N__7734),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5439),
            .DIN0(D_LL_040_in_2),
            .DOUT0(N__3568),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TCI_CPUn_obuf_iopad.PULLUP=1'b1;
    IO_PAD TCI_CPUn_obuf_iopad (
            .OE(N__7727),
            .DIN(N__7726),
            .DOUT(N__7725),
            .PACKAGEPIN(TCI_CPUn));
    defparam TCI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TCI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TCI_CPUn_obuf_preio (
            .PADOEN(N__7727),
            .PADOUT(N__7726),
            .PADIN(N__7725),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2882),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMB_obuf_iopad (
            .OE(N__7718),
            .DIN(N__7717),
            .DOUT(N__7716),
            .PACKAGEPIN(CLKRAMB));
    defparam CLKRAMB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMB_obuf_preio (
            .PADOEN(N__7718),
            .PADOUT(N__7717),
            .PADIN(N__7716),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4426),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_2_iopad (
            .OE(N__7709),
            .DIN(N__7708),
            .DOUT(N__7707),
            .PACKAGEPIN(D_LL_AMIGA[2]));
    defparam D_LL_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_2_preio (
            .PADOEN(N__7709),
            .PADOUT(N__7708),
            .PADIN(N__7707),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2574),
            .DIN0(D_LL_AMIGA_in_2),
            .DOUT0(N__3121),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_4_iopad (
            .OE(N__7700),
            .DIN(N__7699),
            .DOUT(N__7698),
            .PACKAGEPIN(D_UM_AMIGA[4]));
    defparam D_UM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_4_preio (
            .PADOEN(N__7700),
            .PADOUT(N__7699),
            .PADIN(N__7698),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2472),
            .DIN0(D_UM_AMIGA_in_4),
            .DOUT0(N__4168),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_2_iopad (
            .OE(N__7691),
            .DIN(N__7690),
            .DOUT(N__7689),
            .PACKAGEPIN(D_UU_AMIGA[2]));
    defparam D_UU_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_2_preio (
            .PADOEN(N__7691),
            .PADOUT(N__7690),
            .PADIN(N__7689),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2474),
            .DIN0(D_UU_AMIGA_in_2),
            .DOUT0(N__3604),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__7682),
            .DIN(N__7681),
            .DOUT(N__7680),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__7682),
            .PADOUT(N__7681),
            .PADIN(N__7680),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3820),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_6_iopad (
            .OE(N__7673),
            .DIN(N__7672),
            .DOUT(N__7671),
            .PACKAGEPIN(D_LM_AMIGA[6]));
    defparam D_LM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_6_preio (
            .PADOEN(N__7673),
            .PADOUT(N__7672),
            .PADIN(N__7671),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2453),
            .DIN0(D_LM_AMIGA_in_6),
            .DOUT0(N__2821),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam RnW_ibuf_iopad.PULLUP=1'b1;
    IO_PAD RnW_ibuf_iopad (
            .OE(N__7664),
            .DIN(N__7663),
            .DOUT(N__7662),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__7664),
            .PADOUT(N__7663),
            .PADIN(N__7662),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_5_iopad (
            .OE(N__7655),
            .DIN(N__7654),
            .DOUT(N__7653),
            .PACKAGEPIN(D_LM_040[5]));
    defparam D_LM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_5_preio (
            .PADOEN(N__7655),
            .PADOUT(N__7654),
            .PADIN(N__7653),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5331),
            .DIN0(D_LM_040_in_5),
            .DOUT0(N__3037),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_6_iopad (
            .OE(N__7646),
            .DIN(N__7645),
            .DOUT(N__7644),
            .PACKAGEPIN(D_UM_040[6]));
    defparam D_UM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_6_preio (
            .PADOEN(N__7646),
            .PADOUT(N__7645),
            .PADIN(N__7644),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5224),
            .DIN0(D_UM_040_in_6),
            .DOUT0(N__6481),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMAn_obuf_iopad (
            .OE(N__7637),
            .DIN(N__7636),
            .DOUT(N__7635),
            .PACKAGEPIN(DMAn));
    defparam DMAn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMAn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMAn_obuf_preio (
            .PADOEN(N__7637),
            .PADOUT(N__7636),
            .PADIN(N__7635),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2896),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_6_iopad (
            .OE(N__7628),
            .DIN(N__7627),
            .DOUT(N__7626),
            .PACKAGEPIN(D_LL_040[6]));
    defparam D_LL_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_6_preio (
            .PADOEN(N__7628),
            .PADOUT(N__7627),
            .PADIN(N__7626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5426),
            .DIN0(D_LL_040_in_6),
            .DOUT0(N__3502),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_5_iopad (
            .OE(N__7619),
            .DIN(N__7618),
            .DOUT(N__7617),
            .PACKAGEPIN(D_LL_AMIGA[5]));
    defparam D_LL_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_5_preio (
            .PADOEN(N__7619),
            .PADOUT(N__7618),
            .PADIN(N__7617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2559),
            .DIN0(D_LL_AMIGA_in_5),
            .DOUT0(N__4984),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_0_iopad (
            .OE(N__7610),
            .DIN(N__7609),
            .DOUT(N__7608),
            .PACKAGEPIN(D_UM_AMIGA[0]));
    defparam D_UM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_0_preio (
            .PADOEN(N__7610),
            .PADOUT(N__7609),
            .PADIN(N__7608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2530),
            .DIN0(D_UM_AMIGA_in_0),
            .DOUT0(N__4258),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_2_iopad (
            .OE(N__7601),
            .DIN(N__7600),
            .DOUT(N__7599),
            .PACKAGEPIN(D_UU_040[2]));
    defparam D_UU_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_2_preio (
            .PADOEN(N__7601),
            .PADOUT(N__7600),
            .PADIN(N__7599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5382),
            .DIN0(D_UU_040_in_2),
            .DOUT0(N__5512),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_2_iopad (
            .OE(N__7592),
            .DIN(N__7591),
            .DOUT(N__7590),
            .PACKAGEPIN(D_LM_AMIGA[2]));
    defparam D_LM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_2_preio (
            .PADOEN(N__7592),
            .PADOUT(N__7591),
            .PADIN(N__7590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2529),
            .DIN0(D_LM_AMIGA_in_2),
            .DOUT0(N__3636),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK80_CPU_obuf_iopad (
            .OE(N__7583),
            .DIN(N__7582),
            .DOUT(N__7581),
            .PACKAGEPIN(CLK80_CPU));
    defparam CLK80_CPU_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK80_CPU_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK80_CPU_obuf_preio (
            .PADOEN(N__7583),
            .PADOUT(N__7582),
            .PADIN(N__7581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4422),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_3_iopad (
            .OE(N__7574),
            .DIN(N__7573),
            .DOUT(N__7572),
            .PACKAGEPIN(D_LL_040[3]));
    defparam D_LL_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_3_preio (
            .PADOEN(N__7574),
            .PADOUT(N__7573),
            .PADIN(N__7572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5456),
            .DIN0(D_LL_040_in_3),
            .DOUT0(N__3970),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_1_iopad (
            .OE(N__7565),
            .DIN(N__7564),
            .DOUT(N__7563),
            .PACKAGEPIN(D_LM_040[1]));
    defparam D_LM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_1_preio (
            .PADOEN(N__7565),
            .PADOUT(N__7564),
            .PADIN(N__7563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5421),
            .DIN0(D_LM_040_in_1),
            .DOUT0(N__4543),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TSn_obuf_iopad.PULLUP=1'b1;
    IO_PAD TSn_obuf_iopad (
            .OE(N__7556),
            .DIN(N__7555),
            .DOUT(N__7554),
            .PACKAGEPIN(TSn));
    defparam TSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TSn_obuf_preio (
            .PADOEN(N__7556),
            .PADOUT(N__7555),
            .PADIN(N__7554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3292),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_7_iopad (
            .OE(N__7547),
            .DIN(N__7546),
            .DOUT(N__7545),
            .PACKAGEPIN(D_UM_AMIGA[7]));
    defparam D_UM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_7_preio (
            .PADOEN(N__7547),
            .PADOUT(N__7546),
            .PADIN(N__7545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2507),
            .DIN0(D_UM_AMIGA_in_7),
            .DOUT0(N__3364),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_7_iopad (
            .OE(N__7538),
            .DIN(N__7537),
            .DOUT(N__7536),
            .PACKAGEPIN(D_LM_AMIGA[7]));
    defparam D_LM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_7_preio (
            .PADOEN(N__7538),
            .PADOUT(N__7537),
            .PADIN(N__7536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2452),
            .DIN0(D_LM_AMIGA_in_7),
            .DOUT0(N__4063),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PORTSIZE_ibuf_iopad.PULLUP=1'b1;
    IO_PAD PORTSIZE_ibuf_iopad (
            .OE(N__7529),
            .DIN(N__7528),
            .DOUT(N__7527),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PORTSIZE_ibuf_preio (
            .PADOEN(N__7529),
            .PADOUT(N__7528),
            .PADIN(N__7527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PORTSIZE_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_0_iopad (
            .OE(N__7520),
            .DIN(N__7519),
            .DOUT(N__7518),
            .PACKAGEPIN(A_AMIGA[0]));
    defparam A_AMIGA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_0_preio (
            .PADOEN(N__7520),
            .PADOUT(N__7519),
            .PADIN(N__7518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2593),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_4_iopad (
            .OE(N__7511),
            .DIN(N__7510),
            .DOUT(N__7509),
            .PACKAGEPIN(D_LM_040[4]));
    defparam D_LM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_4_preio (
            .PADOEN(N__7511),
            .PADOUT(N__7510),
            .PADIN(N__7509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5353),
            .DIN0(D_LM_040_in_4),
            .DOUT0(N__3223),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_7_iopad (
            .OE(N__7502),
            .DIN(N__7501),
            .DOUT(N__7500),
            .PACKAGEPIN(D_UM_040[7]));
    defparam D_UM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_7_preio (
            .PADOEN(N__7502),
            .PADOUT(N__7501),
            .PADIN(N__7500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5416),
            .DIN0(D_UM_040_in_7),
            .DOUT0(N__6931),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__7493),
            .DIN(N__7492),
            .DOUT(N__7491),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__7493),
            .PADOUT(N__7492),
            .PADIN(N__7491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_1_iopad (
            .OE(N__7484),
            .DIN(N__7483),
            .DOUT(N__7482),
            .PACKAGEPIN(D_UU_AMIGA[1]));
    defparam D_UU_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_1_preio (
            .PADOEN(N__7484),
            .PADOUT(N__7483),
            .PADIN(N__7482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2467),
            .DIN0(D_UU_AMIGA_in_1),
            .DOUT0(N__3742),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__7475),
            .DIN(N__7474),
            .DOUT(N__7473),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__7475),
            .PADOUT(N__7474),
            .PADIN(N__7473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4520),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_0_iopad (
            .OE(N__7466),
            .DIN(N__7465),
            .DOUT(N__7464),
            .PACKAGEPIN(D_UM_040[0]));
    defparam D_UM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_0_preio (
            .PADOEN(N__7466),
            .PADOUT(N__7465),
            .PADIN(N__7464),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5330),
            .DIN0(D_UM_040_in_0),
            .DOUT0(N__5500),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_0_iopad (
            .OE(N__7457),
            .DIN(N__7456),
            .DOUT(N__7455),
            .PACKAGEPIN(D_LL_AMIGA[0]));
    defparam D_LL_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_0_preio (
            .PADOEN(N__7457),
            .PADOUT(N__7456),
            .PADIN(N__7455),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2578),
            .DIN0(D_LL_AMIGA_in_0),
            .DOUT0(N__4315),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_4_iopad (
            .OE(N__7448),
            .DIN(N__7447),
            .DOUT(N__7446),
            .PACKAGEPIN(D_UU_AMIGA[4]));
    defparam D_UU_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_4_preio (
            .PADOEN(N__7448),
            .PADOUT(N__7447),
            .PADIN(N__7446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2473),
            .DIN0(D_UU_AMIGA_in_4),
            .DOUT0(N__3673),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_7_iopad (
            .OE(N__7439),
            .DIN(N__7438),
            .DOUT(N__7437),
            .PACKAGEPIN(D_UU_040[7]));
    defparam D_UU_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_7_preio (
            .PADOEN(N__7439),
            .PADOUT(N__7438),
            .PADIN(N__7437),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5384),
            .DIN0(D_UU_040_in_7),
            .DOUT0(N__5578),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SIZ_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__7430),
            .DIN(N__7429),
            .DOUT(N__7428),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__7430),
            .PADOUT(N__7429),
            .PADIN(N__7428),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam BGn_ibuf_iopad.PULLUP=1'b1;
    IO_PAD BGn_ibuf_iopad (
            .OE(N__7421),
            .DIN(N__7420),
            .DOUT(N__7419),
            .PACKAGEPIN(BGn));
    defparam BGn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BGn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BGn_ibuf_preio (
            .PADOEN(N__7421),
            .PADOUT(N__7420),
            .PADIN(N__7419),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BGn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_0_iopad (
            .OE(N__7412),
            .DIN(N__7411),
            .DOUT(N__7410),
            .PACKAGEPIN(D_LL_040[0]));
    defparam D_LL_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_0_preio (
            .PADOEN(N__7412),
            .PADOUT(N__7411),
            .PADIN(N__7410),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5457),
            .DIN0(D_LL_040_in_0),
            .DOUT0(N__3325),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_2_iopad (
            .OE(N__7403),
            .DIN(N__7402),
            .DOUT(N__7401),
            .PACKAGEPIN(D_UM_AMIGA[2]));
    defparam D_UM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_2_preio (
            .PADOEN(N__7403),
            .PADOUT(N__7402),
            .PADIN(N__7401),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2513),
            .DIN0(D_UM_AMIGA_in_2),
            .DOUT0(N__3070),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_0_iopad (
            .OE(N__7394),
            .DIN(N__7393),
            .DOUT(N__7392),
            .PACKAGEPIN(D_UU_040[0]));
    defparam D_UU_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_0_preio (
            .PADOEN(N__7394),
            .PADOUT(N__7393),
            .PADIN(N__7392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5383),
            .DIN0(D_UU_040_in_0),
            .DOUT0(N__6868),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_0_iopad (
            .OE(N__7385),
            .DIN(N__7384),
            .DOUT(N__7383),
            .PACKAGEPIN(A_040[0]));
    defparam A_040_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_0_preio (
            .PADOEN(N__7385),
            .PADOUT(N__7384),
            .PADIN(N__7383),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_0_iopad (
            .OE(N__7376),
            .DIN(N__7375),
            .DOUT(N__7374),
            .PACKAGEPIN(D_LM_AMIGA[0]));
    defparam D_LM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_0_preio (
            .PADOEN(N__7376),
            .PADOUT(N__7375),
            .PADIN(N__7374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2451),
            .DIN0(D_LM_AMIGA_in_0),
            .DOUT0(N__2746),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBI_CPUn_obuf_iopad (
            .OE(N__7367),
            .DIN(N__7366),
            .DOUT(N__7365),
            .PACKAGEPIN(TBI_CPUn));
    defparam TBI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TBI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TBI_CPUn_obuf_preio (
            .PADOEN(N__7367),
            .PADOUT(N__7366),
            .PADIN(N__7365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4585),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40A_obuf_iopad (
            .OE(N__7358),
            .DIN(N__7357),
            .DOUT(N__7356),
            .PACKAGEPIN(CLK40A));
    defparam CLK40A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40A_obuf_preio (
            .PADOEN(N__7358),
            .PADOUT(N__7357),
            .PADIN(N__7356),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4519),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_3_iopad (
            .OE(N__7349),
            .DIN(N__7348),
            .DOUT(N__7347),
            .PACKAGEPIN(D_LM_040[3]));
    defparam D_LM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_3_preio (
            .PADOEN(N__7349),
            .PADOUT(N__7348),
            .PADIN(N__7347),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5392),
            .DIN0(D_LM_040_in_3),
            .DOUT0(N__2665),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1874 (
            .O(N__7330),
            .I(N__7327));
    LocalMux I__1873 (
            .O(N__7327),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ));
    InMux I__1872 (
            .O(N__7324),
            .I(N__7321));
    LocalMux I__1871 (
            .O(N__7321),
            .I(N__7316));
    InMux I__1870 (
            .O(N__7320),
            .I(N__7313));
    InMux I__1869 (
            .O(N__7319),
            .I(N__7310));
    Span4Mux_v I__1868 (
            .O(N__7316),
            .I(N__7307));
    LocalMux I__1867 (
            .O(N__7313),
            .I(N__7302));
    LocalMux I__1866 (
            .O(N__7310),
            .I(N__7302));
    Span4Mux_v I__1865 (
            .O(N__7307),
            .I(N__7299));
    Span4Mux_v I__1864 (
            .O(N__7302),
            .I(N__7296));
    Sp12to4 I__1863 (
            .O(N__7299),
            .I(N__7293));
    Span4Mux_v I__1862 (
            .O(N__7296),
            .I(N__7290));
    Span12Mux_h I__1861 (
            .O(N__7293),
            .I(N__7287));
    Sp12to4 I__1860 (
            .O(N__7290),
            .I(N__7284));
    Span12Mux_v I__1859 (
            .O(N__7287),
            .I(N__7281));
    Span12Mux_h I__1858 (
            .O(N__7284),
            .I(N__7278));
    Odrv12 I__1857 (
            .O(N__7281),
            .I(D_UM_AMIGA_in_4));
    Odrv12 I__1856 (
            .O(N__7278),
            .I(D_UM_AMIGA_in_4));
    InMux I__1855 (
            .O(N__7273),
            .I(N__7267));
    InMux I__1854 (
            .O(N__7272),
            .I(N__7267));
    LocalMux I__1853 (
            .O(N__7267),
            .I(N__7264));
    Span4Mux_v I__1852 (
            .O(N__7264),
            .I(N__7254));
    InMux I__1851 (
            .O(N__7263),
            .I(N__7251));
    InMux I__1850 (
            .O(N__7262),
            .I(N__7243));
    InMux I__1849 (
            .O(N__7261),
            .I(N__7243));
    InMux I__1848 (
            .O(N__7260),
            .I(N__7234));
    InMux I__1847 (
            .O(N__7259),
            .I(N__7234));
    InMux I__1846 (
            .O(N__7258),
            .I(N__7234));
    InMux I__1845 (
            .O(N__7257),
            .I(N__7234));
    Sp12to4 I__1844 (
            .O(N__7254),
            .I(N__7224));
    LocalMux I__1843 (
            .O(N__7251),
            .I(N__7221));
    InMux I__1842 (
            .O(N__7250),
            .I(N__7216));
    InMux I__1841 (
            .O(N__7249),
            .I(N__7216));
    InMux I__1840 (
            .O(N__7248),
            .I(N__7213));
    LocalMux I__1839 (
            .O(N__7243),
            .I(N__7210));
    LocalMux I__1838 (
            .O(N__7234),
            .I(N__7207));
    InMux I__1837 (
            .O(N__7233),
            .I(N__7200));
    InMux I__1836 (
            .O(N__7232),
            .I(N__7200));
    InMux I__1835 (
            .O(N__7231),
            .I(N__7200));
    InMux I__1834 (
            .O(N__7230),
            .I(N__7195));
    InMux I__1833 (
            .O(N__7229),
            .I(N__7195));
    InMux I__1832 (
            .O(N__7228),
            .I(N__7190));
    InMux I__1831 (
            .O(N__7227),
            .I(N__7190));
    Span12Mux_h I__1830 (
            .O(N__7224),
            .I(N__7185));
    Span4Mux_h I__1829 (
            .O(N__7221),
            .I(N__7180));
    LocalMux I__1828 (
            .O(N__7216),
            .I(N__7180));
    LocalMux I__1827 (
            .O(N__7213),
            .I(N__7177));
    Span4Mux_v I__1826 (
            .O(N__7210),
            .I(N__7170));
    Span4Mux_h I__1825 (
            .O(N__7207),
            .I(N__7170));
    LocalMux I__1824 (
            .O(N__7200),
            .I(N__7170));
    LocalMux I__1823 (
            .O(N__7195),
            .I(N__7165));
    LocalMux I__1822 (
            .O(N__7190),
            .I(N__7165));
    InMux I__1821 (
            .O(N__7189),
            .I(N__7162));
    InMux I__1820 (
            .O(N__7188),
            .I(N__7159));
    Odrv12 I__1819 (
            .O(N__7185),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    Odrv4 I__1818 (
            .O(N__7180),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    Odrv4 I__1817 (
            .O(N__7177),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    Odrv4 I__1816 (
            .O(N__7170),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    Odrv12 I__1815 (
            .O(N__7165),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    LocalMux I__1814 (
            .O(N__7162),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    LocalMux I__1813 (
            .O(N__7159),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    IoInMux I__1812 (
            .O(N__7144),
            .I(N__7141));
    LocalMux I__1811 (
            .O(N__7141),
            .I(N__7138));
    IoSpan4Mux I__1810 (
            .O(N__7138),
            .I(N__7135));
    Span4Mux_s3_v I__1809 (
            .O(N__7135),
            .I(N__7132));
    Sp12to4 I__1808 (
            .O(N__7132),
            .I(N__7129));
    Span12Mux_h I__1807 (
            .O(N__7129),
            .I(N__7126));
    Odrv12 I__1806 (
            .O(N__7126),
            .I(un1_D_UM_AMIGA_4));
    InMux I__1805 (
            .O(N__7123),
            .I(N__7120));
    LocalMux I__1804 (
            .O(N__7120),
            .I(N__7116));
    InMux I__1803 (
            .O(N__7119),
            .I(N__7113));
    Span4Mux_v I__1802 (
            .O(N__7116),
            .I(N__7109));
    LocalMux I__1801 (
            .O(N__7113),
            .I(N__7106));
    InMux I__1800 (
            .O(N__7112),
            .I(N__7103));
    Span4Mux_v I__1799 (
            .O(N__7109),
            .I(N__7100));
    Span4Mux_v I__1798 (
            .O(N__7106),
            .I(N__7095));
    LocalMux I__1797 (
            .O(N__7103),
            .I(N__7095));
    Sp12to4 I__1796 (
            .O(N__7100),
            .I(N__7092));
    Span4Mux_v I__1795 (
            .O(N__7095),
            .I(N__7089));
    Span12Mux_h I__1794 (
            .O(N__7092),
            .I(N__7086));
    Sp12to4 I__1793 (
            .O(N__7089),
            .I(N__7083));
    Span12Mux_v I__1792 (
            .O(N__7086),
            .I(N__7078));
    Span12Mux_h I__1791 (
            .O(N__7083),
            .I(N__7078));
    Odrv12 I__1790 (
            .O(N__7078),
            .I(D_UM_AMIGA_in_3));
    InMux I__1789 (
            .O(N__7075),
            .I(N__7072));
    LocalMux I__1788 (
            .O(N__7072),
            .I(N__7069));
    Odrv12 I__1787 (
            .O(N__7069),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ));
    IoInMux I__1786 (
            .O(N__7066),
            .I(N__7063));
    LocalMux I__1785 (
            .O(N__7063),
            .I(N__7060));
    IoSpan4Mux I__1784 (
            .O(N__7060),
            .I(N__7057));
    IoSpan4Mux I__1783 (
            .O(N__7057),
            .I(N__7054));
    Span4Mux_s2_h I__1782 (
            .O(N__7054),
            .I(N__7051));
    Sp12to4 I__1781 (
            .O(N__7051),
            .I(N__7048));
    Odrv12 I__1780 (
            .O(N__7048),
            .I(un1_D_UM_AMIGA_3));
    CEMux I__1779 (
            .O(N__7045),
            .I(N__7040));
    CEMux I__1778 (
            .O(N__7044),
            .I(N__7037));
    CEMux I__1777 (
            .O(N__7043),
            .I(N__7033));
    LocalMux I__1776 (
            .O(N__7040),
            .I(N__7028));
    LocalMux I__1775 (
            .O(N__7037),
            .I(N__7028));
    CEMux I__1774 (
            .O(N__7036),
            .I(N__7025));
    LocalMux I__1773 (
            .O(N__7033),
            .I(N__7022));
    Span4Mux_v I__1772 (
            .O(N__7028),
            .I(N__7017));
    LocalMux I__1771 (
            .O(N__7025),
            .I(N__7017));
    Span4Mux_h I__1770 (
            .O(N__7022),
            .I(N__7014));
    Span4Mux_h I__1769 (
            .O(N__7017),
            .I(N__7011));
    Odrv4 I__1768 (
            .O(N__7014),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    Odrv4 I__1767 (
            .O(N__7011),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    SRMux I__1766 (
            .O(N__7006),
            .I(N__7000));
    SRMux I__1765 (
            .O(N__7005),
            .I(N__6997));
    SRMux I__1764 (
            .O(N__7004),
            .I(N__6994));
    SRMux I__1763 (
            .O(N__7003),
            .I(N__6991));
    LocalMux I__1762 (
            .O(N__7000),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0 ));
    LocalMux I__1761 (
            .O(N__6997),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0 ));
    LocalMux I__1760 (
            .O(N__6994),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0 ));
    LocalMux I__1759 (
            .O(N__6991),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0 ));
    InMux I__1758 (
            .O(N__6982),
            .I(N__6979));
    LocalMux I__1757 (
            .O(N__6979),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ));
    InMux I__1756 (
            .O(N__6976),
            .I(N__6971));
    InMux I__1755 (
            .O(N__6975),
            .I(N__6968));
    InMux I__1754 (
            .O(N__6974),
            .I(N__6965));
    LocalMux I__1753 (
            .O(N__6971),
            .I(N__6960));
    LocalMux I__1752 (
            .O(N__6968),
            .I(N__6960));
    LocalMux I__1751 (
            .O(N__6965),
            .I(N__6957));
    Span4Mux_v I__1750 (
            .O(N__6960),
            .I(N__6954));
    Span12Mux_v I__1749 (
            .O(N__6957),
            .I(N__6951));
    Span4Mux_v I__1748 (
            .O(N__6954),
            .I(N__6948));
    Span12Mux_h I__1747 (
            .O(N__6951),
            .I(N__6945));
    Sp12to4 I__1746 (
            .O(N__6948),
            .I(N__6942));
    Span12Mux_v I__1745 (
            .O(N__6945),
            .I(N__6939));
    Span12Mux_h I__1744 (
            .O(N__6942),
            .I(N__6936));
    Odrv12 I__1743 (
            .O(N__6939),
            .I(D_UM_AMIGA_in_7));
    Odrv12 I__1742 (
            .O(N__6936),
            .I(D_UM_AMIGA_in_7));
    IoInMux I__1741 (
            .O(N__6931),
            .I(N__6928));
    LocalMux I__1740 (
            .O(N__6928),
            .I(N__6925));
    Sp12to4 I__1739 (
            .O(N__6925),
            .I(N__6922));
    Span12Mux_h I__1738 (
            .O(N__6922),
            .I(N__6919));
    Odrv12 I__1737 (
            .O(N__6919),
            .I(un1_D_UM_AMIGA_7));
    InMux I__1736 (
            .O(N__6916),
            .I(N__6913));
    LocalMux I__1735 (
            .O(N__6913),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ));
    InMux I__1734 (
            .O(N__6910),
            .I(N__6907));
    LocalMux I__1733 (
            .O(N__6907),
            .I(N__6902));
    InMux I__1732 (
            .O(N__6906),
            .I(N__6899));
    InMux I__1731 (
            .O(N__6905),
            .I(N__6896));
    Span4Mux_v I__1730 (
            .O(N__6902),
            .I(N__6893));
    LocalMux I__1729 (
            .O(N__6899),
            .I(N__6888));
    LocalMux I__1728 (
            .O(N__6896),
            .I(N__6888));
    Span4Mux_v I__1727 (
            .O(N__6893),
            .I(N__6885));
    Span4Mux_v I__1726 (
            .O(N__6888),
            .I(N__6882));
    Span4Mux_v I__1725 (
            .O(N__6885),
            .I(N__6877));
    Span4Mux_h I__1724 (
            .O(N__6882),
            .I(N__6877));
    Sp12to4 I__1723 (
            .O(N__6877),
            .I(N__6874));
    Span12Mux_h I__1722 (
            .O(N__6874),
            .I(N__6871));
    Odrv12 I__1721 (
            .O(N__6871),
            .I(D_UU_AMIGA_in_0));
    IoInMux I__1720 (
            .O(N__6868),
            .I(N__6865));
    LocalMux I__1719 (
            .O(N__6865),
            .I(N__6862));
    Span4Mux_s3_v I__1718 (
            .O(N__6862),
            .I(N__6859));
    Span4Mux_h I__1717 (
            .O(N__6859),
            .I(N__6856));
    Span4Mux_h I__1716 (
            .O(N__6856),
            .I(N__6853));
    Span4Mux_v I__1715 (
            .O(N__6853),
            .I(N__6850));
    Odrv4 I__1714 (
            .O(N__6850),
            .I(un1_D_UU_AMIGA_0));
    InMux I__1713 (
            .O(N__6847),
            .I(N__6844));
    LocalMux I__1712 (
            .O(N__6844),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ));
    InMux I__1711 (
            .O(N__6841),
            .I(N__6838));
    LocalMux I__1710 (
            .O(N__6838),
            .I(N__6834));
    InMux I__1709 (
            .O(N__6837),
            .I(N__6831));
    Span4Mux_v I__1708 (
            .O(N__6834),
            .I(N__6826));
    LocalMux I__1707 (
            .O(N__6831),
            .I(N__6826));
    Span4Mux_h I__1706 (
            .O(N__6826),
            .I(N__6822));
    InMux I__1705 (
            .O(N__6825),
            .I(N__6819));
    Span4Mux_h I__1704 (
            .O(N__6822),
            .I(N__6814));
    LocalMux I__1703 (
            .O(N__6819),
            .I(N__6814));
    Span4Mux_v I__1702 (
            .O(N__6814),
            .I(N__6811));
    Sp12to4 I__1701 (
            .O(N__6811),
            .I(N__6808));
    Span12Mux_h I__1700 (
            .O(N__6808),
            .I(N__6805));
    Span12Mux_v I__1699 (
            .O(N__6805),
            .I(N__6802));
    Odrv12 I__1698 (
            .O(N__6802),
            .I(D_UU_AMIGA_in_5));
    IoInMux I__1697 (
            .O(N__6799),
            .I(N__6796));
    LocalMux I__1696 (
            .O(N__6796),
            .I(N__6793));
    Span4Mux_s3_v I__1695 (
            .O(N__6793),
            .I(N__6790));
    Span4Mux_v I__1694 (
            .O(N__6790),
            .I(N__6787));
    Sp12to4 I__1693 (
            .O(N__6787),
            .I(N__6784));
    Span12Mux_h I__1692 (
            .O(N__6784),
            .I(N__6781));
    Odrv12 I__1691 (
            .O(N__6781),
            .I(un1_D_UU_AMIGA_5));
    InMux I__1690 (
            .O(N__6778),
            .I(N__6775));
    LocalMux I__1689 (
            .O(N__6775),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ));
    InMux I__1688 (
            .O(N__6772),
            .I(N__6768));
    InMux I__1687 (
            .O(N__6771),
            .I(N__6765));
    LocalMux I__1686 (
            .O(N__6768),
            .I(N__6761));
    LocalMux I__1685 (
            .O(N__6765),
            .I(N__6758));
    InMux I__1684 (
            .O(N__6764),
            .I(N__6755));
    Span4Mux_v I__1683 (
            .O(N__6761),
            .I(N__6752));
    Span4Mux_v I__1682 (
            .O(N__6758),
            .I(N__6749));
    LocalMux I__1681 (
            .O(N__6755),
            .I(N__6746));
    Sp12to4 I__1680 (
            .O(N__6752),
            .I(N__6743));
    Sp12to4 I__1679 (
            .O(N__6749),
            .I(N__6740));
    Span12Mux_h I__1678 (
            .O(N__6746),
            .I(N__6737));
    Span12Mux_h I__1677 (
            .O(N__6743),
            .I(N__6734));
    Span12Mux_h I__1676 (
            .O(N__6740),
            .I(N__6731));
    Span12Mux_h I__1675 (
            .O(N__6737),
            .I(N__6728));
    Span12Mux_v I__1674 (
            .O(N__6734),
            .I(N__6723));
    Span12Mux_h I__1673 (
            .O(N__6731),
            .I(N__6723));
    Odrv12 I__1672 (
            .O(N__6728),
            .I(D_UM_AMIGA_in_5));
    Odrv12 I__1671 (
            .O(N__6723),
            .I(D_UM_AMIGA_in_5));
    IoInMux I__1670 (
            .O(N__6718),
            .I(N__6715));
    LocalMux I__1669 (
            .O(N__6715),
            .I(N__6712));
    Span4Mux_s2_v I__1668 (
            .O(N__6712),
            .I(N__6709));
    Sp12to4 I__1667 (
            .O(N__6709),
            .I(N__6706));
    Span12Mux_h I__1666 (
            .O(N__6706),
            .I(N__6703));
    Odrv12 I__1665 (
            .O(N__6703),
            .I(un1_D_UM_AMIGA_5));
    InMux I__1664 (
            .O(N__6700),
            .I(N__6697));
    LocalMux I__1663 (
            .O(N__6697),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ));
    InMux I__1662 (
            .O(N__6694),
            .I(N__6690));
    InMux I__1661 (
            .O(N__6693),
            .I(N__6687));
    LocalMux I__1660 (
            .O(N__6690),
            .I(N__6684));
    LocalMux I__1659 (
            .O(N__6687),
            .I(N__6681));
    Span4Mux_h I__1658 (
            .O(N__6684),
            .I(N__6675));
    Span4Mux_v I__1657 (
            .O(N__6681),
            .I(N__6675));
    InMux I__1656 (
            .O(N__6680),
            .I(N__6672));
    Span4Mux_h I__1655 (
            .O(N__6675),
            .I(N__6667));
    LocalMux I__1654 (
            .O(N__6672),
            .I(N__6667));
    Sp12to4 I__1653 (
            .O(N__6667),
            .I(N__6664));
    Span12Mux_v I__1652 (
            .O(N__6664),
            .I(N__6661));
    Span12Mux_h I__1651 (
            .O(N__6661),
            .I(N__6658));
    Odrv12 I__1650 (
            .O(N__6658),
            .I(D_UU_AMIGA_in_3));
    IoInMux I__1649 (
            .O(N__6655),
            .I(N__6652));
    LocalMux I__1648 (
            .O(N__6652),
            .I(N__6649));
    Span12Mux_s0_v I__1647 (
            .O(N__6649),
            .I(N__6646));
    Span12Mux_h I__1646 (
            .O(N__6646),
            .I(N__6643));
    Odrv12 I__1645 (
            .O(N__6643),
            .I(un1_D_UU_AMIGA_3));
    InMux I__1644 (
            .O(N__6640),
            .I(N__6637));
    LocalMux I__1643 (
            .O(N__6637),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ));
    InMux I__1642 (
            .O(N__6634),
            .I(N__6631));
    LocalMux I__1641 (
            .O(N__6631),
            .I(N__6626));
    InMux I__1640 (
            .O(N__6630),
            .I(N__6623));
    InMux I__1639 (
            .O(N__6629),
            .I(N__6620));
    Span4Mux_v I__1638 (
            .O(N__6626),
            .I(N__6617));
    LocalMux I__1637 (
            .O(N__6623),
            .I(N__6612));
    LocalMux I__1636 (
            .O(N__6620),
            .I(N__6612));
    Sp12to4 I__1635 (
            .O(N__6617),
            .I(N__6609));
    Span12Mux_v I__1634 (
            .O(N__6612),
            .I(N__6606));
    Span12Mux_h I__1633 (
            .O(N__6609),
            .I(N__6603));
    Span12Mux_h I__1632 (
            .O(N__6606),
            .I(N__6600));
    Span12Mux_v I__1631 (
            .O(N__6603),
            .I(N__6597));
    Odrv12 I__1630 (
            .O(N__6600),
            .I(D_UU_AMIGA_in_4));
    Odrv12 I__1629 (
            .O(N__6597),
            .I(D_UU_AMIGA_in_4));
    IoInMux I__1628 (
            .O(N__6592),
            .I(N__6589));
    LocalMux I__1627 (
            .O(N__6589),
            .I(N__6586));
    Span4Mux_s2_v I__1626 (
            .O(N__6586),
            .I(N__6583));
    Span4Mux_h I__1625 (
            .O(N__6583),
            .I(N__6580));
    Span4Mux_v I__1624 (
            .O(N__6580),
            .I(N__6577));
    Span4Mux_v I__1623 (
            .O(N__6577),
            .I(N__6574));
    Odrv4 I__1622 (
            .O(N__6574),
            .I(un1_D_UU_AMIGA_4));
    InMux I__1621 (
            .O(N__6571),
            .I(N__6568));
    LocalMux I__1620 (
            .O(N__6568),
            .I(N__6565));
    Odrv4 I__1619 (
            .O(N__6565),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ));
    InMux I__1618 (
            .O(N__6562),
            .I(N__6558));
    InMux I__1617 (
            .O(N__6561),
            .I(N__6555));
    LocalMux I__1616 (
            .O(N__6558),
            .I(N__6551));
    LocalMux I__1615 (
            .O(N__6555),
            .I(N__6548));
    InMux I__1614 (
            .O(N__6554),
            .I(N__6545));
    Span4Mux_v I__1613 (
            .O(N__6551),
            .I(N__6540));
    Span4Mux_v I__1612 (
            .O(N__6548),
            .I(N__6540));
    LocalMux I__1611 (
            .O(N__6545),
            .I(N__6537));
    Span4Mux_h I__1610 (
            .O(N__6540),
            .I(N__6534));
    Span4Mux_v I__1609 (
            .O(N__6537),
            .I(N__6531));
    Sp12to4 I__1608 (
            .O(N__6534),
            .I(N__6526));
    Sp12to4 I__1607 (
            .O(N__6531),
            .I(N__6526));
    Span12Mux_h I__1606 (
            .O(N__6526),
            .I(N__6523));
    Odrv12 I__1605 (
            .O(N__6523),
            .I(D_UU_AMIGA_in_6));
    IoInMux I__1604 (
            .O(N__6520),
            .I(N__6517));
    LocalMux I__1603 (
            .O(N__6517),
            .I(N__6514));
    Span4Mux_s2_v I__1602 (
            .O(N__6514),
            .I(N__6511));
    Span4Mux_h I__1601 (
            .O(N__6511),
            .I(N__6508));
    Sp12to4 I__1600 (
            .O(N__6508),
            .I(N__6505));
    Span12Mux_s8_v I__1599 (
            .O(N__6505),
            .I(N__6502));
    Odrv12 I__1598 (
            .O(N__6502),
            .I(un1_D_UU_AMIGA_6));
    IoInMux I__1597 (
            .O(N__6499),
            .I(N__6496));
    LocalMux I__1596 (
            .O(N__6496),
            .I(N__6493));
    Span4Mux_s2_h I__1595 (
            .O(N__6493),
            .I(N__6490));
    Sp12to4 I__1594 (
            .O(N__6490),
            .I(N__6487));
    Span12Mux_v I__1593 (
            .O(N__6487),
            .I(N__6484));
    Odrv12 I__1592 (
            .O(N__6484),
            .I(un1_D_UM_AMIGA_2));
    IoInMux I__1591 (
            .O(N__6481),
            .I(N__6478));
    LocalMux I__1590 (
            .O(N__6478),
            .I(N__6475));
    Sp12to4 I__1589 (
            .O(N__6475),
            .I(N__6472));
    Span12Mux_h I__1588 (
            .O(N__6472),
            .I(N__6469));
    Odrv12 I__1587 (
            .O(N__6469),
            .I(un1_D_UM_AMIGA_6));
    InMux I__1586 (
            .O(N__6466),
            .I(N__6463));
    LocalMux I__1585 (
            .O(N__6463),
            .I(N__6460));
    Span4Mux_v I__1584 (
            .O(N__6460),
            .I(N__6455));
    InMux I__1583 (
            .O(N__6459),
            .I(N__6452));
    InMux I__1582 (
            .O(N__6458),
            .I(N__6449));
    Span4Mux_v I__1581 (
            .O(N__6455),
            .I(N__6446));
    LocalMux I__1580 (
            .O(N__6452),
            .I(N__6443));
    LocalMux I__1579 (
            .O(N__6449),
            .I(N__6440));
    Span4Mux_v I__1578 (
            .O(N__6446),
            .I(N__6433));
    Span4Mux_v I__1577 (
            .O(N__6443),
            .I(N__6433));
    Span4Mux_v I__1576 (
            .O(N__6440),
            .I(N__6433));
    Sp12to4 I__1575 (
            .O(N__6433),
            .I(N__6430));
    Span12Mux_h I__1574 (
            .O(N__6430),
            .I(N__6427));
    Odrv12 I__1573 (
            .O(N__6427),
            .I(D_UM_AMIGA_in_0));
    InMux I__1572 (
            .O(N__6424),
            .I(N__6421));
    LocalMux I__1571 (
            .O(N__6421),
            .I(N__6418));
    Odrv4 I__1570 (
            .O(N__6418),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ));
    InMux I__1569 (
            .O(N__6415),
            .I(N__6412));
    LocalMux I__1568 (
            .O(N__6412),
            .I(N__6408));
    InMux I__1567 (
            .O(N__6411),
            .I(N__6405));
    Span4Mux_v I__1566 (
            .O(N__6408),
            .I(N__6402));
    LocalMux I__1565 (
            .O(N__6405),
            .I(N__6398));
    Span4Mux_v I__1564 (
            .O(N__6402),
            .I(N__6395));
    InMux I__1563 (
            .O(N__6401),
            .I(N__6392));
    Span4Mux_v I__1562 (
            .O(N__6398),
            .I(N__6389));
    Sp12to4 I__1561 (
            .O(N__6395),
            .I(N__6382));
    LocalMux I__1560 (
            .O(N__6392),
            .I(N__6382));
    Sp12to4 I__1559 (
            .O(N__6389),
            .I(N__6382));
    Span12Mux_h I__1558 (
            .O(N__6382),
            .I(N__6379));
    Span12Mux_v I__1557 (
            .O(N__6379),
            .I(N__6376));
    Odrv12 I__1556 (
            .O(N__6376),
            .I(D_UM_AMIGA_in_6));
    InMux I__1555 (
            .O(N__6373),
            .I(N__6370));
    LocalMux I__1554 (
            .O(N__6370),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ));
    InMux I__1553 (
            .O(N__6367),
            .I(N__6364));
    LocalMux I__1552 (
            .O(N__6364),
            .I(N__6361));
    Span4Mux_v I__1551 (
            .O(N__6361),
            .I(N__6356));
    InMux I__1550 (
            .O(N__6360),
            .I(N__6353));
    InMux I__1549 (
            .O(N__6359),
            .I(N__6350));
    Span4Mux_v I__1548 (
            .O(N__6356),
            .I(N__6347));
    LocalMux I__1547 (
            .O(N__6353),
            .I(N__6342));
    LocalMux I__1546 (
            .O(N__6350),
            .I(N__6342));
    Span4Mux_v I__1545 (
            .O(N__6347),
            .I(N__6339));
    Span4Mux_v I__1544 (
            .O(N__6342),
            .I(N__6336));
    Sp12to4 I__1543 (
            .O(N__6339),
            .I(N__6331));
    Sp12to4 I__1542 (
            .O(N__6336),
            .I(N__6331));
    Span12Mux_h I__1541 (
            .O(N__6331),
            .I(N__6328));
    Odrv12 I__1540 (
            .O(N__6328),
            .I(D_UM_AMIGA_in_2));
    InMux I__1539 (
            .O(N__6325),
            .I(N__6322));
    LocalMux I__1538 (
            .O(N__6322),
            .I(N__6319));
    Odrv4 I__1537 (
            .O(N__6319),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ));
    IoInMux I__1536 (
            .O(N__6316),
            .I(N__6313));
    LocalMux I__1535 (
            .O(N__6313),
            .I(N__6310));
    IoSpan4Mux I__1534 (
            .O(N__6310),
            .I(N__6307));
    Span4Mux_s3_v I__1533 (
            .O(N__6307),
            .I(N__6304));
    Span4Mux_v I__1532 (
            .O(N__6304),
            .I(N__6298));
    InMux I__1531 (
            .O(N__6303),
            .I(N__6295));
    InMux I__1530 (
            .O(N__6302),
            .I(N__6290));
    InMux I__1529 (
            .O(N__6301),
            .I(N__6290));
    Span4Mux_v I__1528 (
            .O(N__6298),
            .I(N__6283));
    LocalMux I__1527 (
            .O(N__6295),
            .I(N__6283));
    LocalMux I__1526 (
            .O(N__6290),
            .I(N__6283));
    Span4Mux_v I__1525 (
            .O(N__6283),
            .I(N__6279));
    InMux I__1524 (
            .O(N__6282),
            .I(N__6276));
    Span4Mux_h I__1523 (
            .O(N__6279),
            .I(N__6272));
    LocalMux I__1522 (
            .O(N__6276),
            .I(N__6269));
    InMux I__1521 (
            .O(N__6275),
            .I(N__6266));
    Sp12to4 I__1520 (
            .O(N__6272),
            .I(N__6261));
    Span12Mux_h I__1519 (
            .O(N__6269),
            .I(N__6261));
    LocalMux I__1518 (
            .O(N__6266),
            .I(N__6258));
    Span12Mux_v I__1517 (
            .O(N__6261),
            .I(N__6253));
    Span12Mux_h I__1516 (
            .O(N__6258),
            .I(N__6253));
    Odrv12 I__1515 (
            .O(N__6253),
            .I(TACKn_in));
    CascadeMux I__1514 (
            .O(N__6250),
            .I(N__6243));
    InMux I__1513 (
            .O(N__6249),
            .I(N__6236));
    InMux I__1512 (
            .O(N__6248),
            .I(N__6233));
    InMux I__1511 (
            .O(N__6247),
            .I(N__6228));
    InMux I__1510 (
            .O(N__6246),
            .I(N__6228));
    InMux I__1509 (
            .O(N__6243),
            .I(N__6225));
    InMux I__1508 (
            .O(N__6242),
            .I(N__6218));
    InMux I__1507 (
            .O(N__6241),
            .I(N__6218));
    InMux I__1506 (
            .O(N__6240),
            .I(N__6218));
    InMux I__1505 (
            .O(N__6239),
            .I(N__6215));
    LocalMux I__1504 (
            .O(N__6236),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1503 (
            .O(N__6233),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1502 (
            .O(N__6228),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1501 (
            .O(N__6225),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1500 (
            .O(N__6218),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1499 (
            .O(N__6215),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    CascadeMux I__1498 (
            .O(N__6202),
            .I(N__6194));
    InMux I__1497 (
            .O(N__6201),
            .I(N__6188));
    InMux I__1496 (
            .O(N__6200),
            .I(N__6183));
    InMux I__1495 (
            .O(N__6199),
            .I(N__6183));
    InMux I__1494 (
            .O(N__6198),
            .I(N__6178));
    InMux I__1493 (
            .O(N__6197),
            .I(N__6178));
    InMux I__1492 (
            .O(N__6194),
            .I(N__6175));
    InMux I__1491 (
            .O(N__6193),
            .I(N__6170));
    InMux I__1490 (
            .O(N__6192),
            .I(N__6170));
    InMux I__1489 (
            .O(N__6191),
            .I(N__6167));
    LocalMux I__1488 (
            .O(N__6188),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1487 (
            .O(N__6183),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1486 (
            .O(N__6178),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1485 (
            .O(N__6175),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1484 (
            .O(N__6170),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1483 (
            .O(N__6167),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    CascadeMux I__1482 (
            .O(N__6154),
            .I(N__6149));
    InMux I__1481 (
            .O(N__6153),
            .I(N__6144));
    InMux I__1480 (
            .O(N__6152),
            .I(N__6141));
    InMux I__1479 (
            .O(N__6149),
            .I(N__6138));
    CascadeMux I__1478 (
            .O(N__6148),
            .I(N__6134));
    InMux I__1477 (
            .O(N__6147),
            .I(N__6131));
    LocalMux I__1476 (
            .O(N__6144),
            .I(N__6122));
    LocalMux I__1475 (
            .O(N__6141),
            .I(N__6122));
    LocalMux I__1474 (
            .O(N__6138),
            .I(N__6122));
    InMux I__1473 (
            .O(N__6137),
            .I(N__6117));
    InMux I__1472 (
            .O(N__6134),
            .I(N__6117));
    LocalMux I__1471 (
            .O(N__6131),
            .I(N__6114));
    InMux I__1470 (
            .O(N__6130),
            .I(N__6109));
    InMux I__1469 (
            .O(N__6129),
            .I(N__6109));
    Span4Mux_v I__1468 (
            .O(N__6122),
            .I(N__6106));
    LocalMux I__1467 (
            .O(N__6117),
            .I(N__6103));
    Span4Mux_h I__1466 (
            .O(N__6114),
            .I(N__6098));
    LocalMux I__1465 (
            .O(N__6109),
            .I(N__6098));
    Span4Mux_v I__1464 (
            .O(N__6106),
            .I(N__6095));
    Span4Mux_v I__1463 (
            .O(N__6103),
            .I(N__6089));
    Span4Mux_v I__1462 (
            .O(N__6098),
            .I(N__6089));
    Span4Mux_h I__1461 (
            .O(N__6095),
            .I(N__6086));
    InMux I__1460 (
            .O(N__6094),
            .I(N__6083));
    Span4Mux_h I__1459 (
            .O(N__6089),
            .I(N__6080));
    Span4Mux_v I__1458 (
            .O(N__6086),
            .I(N__6075));
    LocalMux I__1457 (
            .O(N__6083),
            .I(N__6075));
    Sp12to4 I__1456 (
            .O(N__6080),
            .I(N__6072));
    Span4Mux_v I__1455 (
            .O(N__6075),
            .I(N__6069));
    Span12Mux_s11_h I__1454 (
            .O(N__6072),
            .I(N__6066));
    Span4Mux_h I__1453 (
            .O(N__6069),
            .I(N__6063));
    Span12Mux_v I__1452 (
            .O(N__6066),
            .I(N__6058));
    Sp12to4 I__1451 (
            .O(N__6063),
            .I(N__6058));
    Odrv12 I__1450 (
            .O(N__6058),
            .I(RESETn_c));
    CascadeMux I__1449 (
            .O(N__6055),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_ ));
    IoInMux I__1448 (
            .O(N__6052),
            .I(N__6049));
    LocalMux I__1447 (
            .O(N__6049),
            .I(N__6046));
    Span4Mux_s3_v I__1446 (
            .O(N__6046),
            .I(N__6042));
    InMux I__1445 (
            .O(N__6045),
            .I(N__6038));
    Span4Mux_h I__1444 (
            .O(N__6042),
            .I(N__6034));
    InMux I__1443 (
            .O(N__6041),
            .I(N__6031));
    LocalMux I__1442 (
            .O(N__6038),
            .I(N__6028));
    InMux I__1441 (
            .O(N__6037),
            .I(N__6025));
    Span4Mux_v I__1440 (
            .O(N__6034),
            .I(N__6020));
    LocalMux I__1439 (
            .O(N__6031),
            .I(N__6020));
    Span4Mux_h I__1438 (
            .O(N__6028),
            .I(N__6015));
    LocalMux I__1437 (
            .O(N__6025),
            .I(N__6015));
    Span4Mux_v I__1436 (
            .O(N__6020),
            .I(N__6012));
    Sp12to4 I__1435 (
            .O(N__6015),
            .I(N__6009));
    Sp12to4 I__1434 (
            .O(N__6012),
            .I(N__6006));
    Span12Mux_s11_v I__1433 (
            .O(N__6009),
            .I(N__6003));
    Span12Mux_h I__1432 (
            .O(N__6006),
            .I(N__6000));
    Span12Mux_h I__1431 (
            .O(N__6003),
            .I(N__5997));
    Odrv12 I__1430 (
            .O(N__6000),
            .I(RnW_c));
    Odrv12 I__1429 (
            .O(N__5997),
            .I(RnW_c));
    CascadeMux I__1428 (
            .O(N__5992),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0_cascade_ ));
    InMux I__1427 (
            .O(N__5989),
            .I(N__5986));
    LocalMux I__1426 (
            .O(N__5986),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa ));
    InMux I__1425 (
            .O(N__5983),
            .I(N__5980));
    LocalMux I__1424 (
            .O(N__5980),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ));
    InMux I__1423 (
            .O(N__5977),
            .I(N__5974));
    LocalMux I__1422 (
            .O(N__5974),
            .I(N__5969));
    InMux I__1421 (
            .O(N__5973),
            .I(N__5966));
    InMux I__1420 (
            .O(N__5972),
            .I(N__5963));
    Span4Mux_v I__1419 (
            .O(N__5969),
            .I(N__5960));
    LocalMux I__1418 (
            .O(N__5966),
            .I(N__5955));
    LocalMux I__1417 (
            .O(N__5963),
            .I(N__5955));
    Span4Mux_v I__1416 (
            .O(N__5960),
            .I(N__5952));
    Span4Mux_v I__1415 (
            .O(N__5955),
            .I(N__5949));
    Span4Mux_v I__1414 (
            .O(N__5952),
            .I(N__5946));
    Span4Mux_v I__1413 (
            .O(N__5949),
            .I(N__5943));
    Sp12to4 I__1412 (
            .O(N__5946),
            .I(N__5938));
    Sp12to4 I__1411 (
            .O(N__5943),
            .I(N__5938));
    Span12Mux_h I__1410 (
            .O(N__5938),
            .I(N__5935));
    Odrv12 I__1409 (
            .O(N__5935),
            .I(D_UU_AMIGA_in_1));
    IoInMux I__1408 (
            .O(N__5932),
            .I(N__5929));
    LocalMux I__1407 (
            .O(N__5929),
            .I(N__5926));
    IoSpan4Mux I__1406 (
            .O(N__5926),
            .I(N__5923));
    Span4Mux_s3_h I__1405 (
            .O(N__5923),
            .I(N__5920));
    Sp12to4 I__1404 (
            .O(N__5920),
            .I(N__5917));
    Span12Mux_h I__1403 (
            .O(N__5917),
            .I(N__5914));
    Odrv12 I__1402 (
            .O(N__5914),
            .I(un1_D_UU_AMIGA_1));
    InMux I__1401 (
            .O(N__5911),
            .I(N__5908));
    LocalMux I__1400 (
            .O(N__5908),
            .I(N__5905));
    Sp12to4 I__1399 (
            .O(N__5905),
            .I(N__5900));
    InMux I__1398 (
            .O(N__5904),
            .I(N__5897));
    CascadeMux I__1397 (
            .O(N__5903),
            .I(N__5894));
    Span12Mux_v I__1396 (
            .O(N__5900),
            .I(N__5891));
    LocalMux I__1395 (
            .O(N__5897),
            .I(N__5888));
    InMux I__1394 (
            .O(N__5894),
            .I(N__5885));
    Odrv12 I__1393 (
            .O(N__5891),
            .I(\U111_CYCLE_SM.TA_ENZ0 ));
    Odrv4 I__1392 (
            .O(N__5888),
            .I(\U111_CYCLE_SM.TA_ENZ0 ));
    LocalMux I__1391 (
            .O(N__5885),
            .I(\U111_CYCLE_SM.TA_ENZ0 ));
    InMux I__1390 (
            .O(N__5878),
            .I(N__5875));
    LocalMux I__1389 (
            .O(N__5875),
            .I(N__5872));
    Span4Mux_v I__1388 (
            .O(N__5872),
            .I(N__5868));
    CascadeMux I__1387 (
            .O(N__5871),
            .I(N__5863));
    Span4Mux_v I__1386 (
            .O(N__5868),
            .I(N__5860));
    InMux I__1385 (
            .O(N__5867),
            .I(N__5857));
    InMux I__1384 (
            .O(N__5866),
            .I(N__5854));
    InMux I__1383 (
            .O(N__5863),
            .I(N__5851));
    Span4Mux_v I__1382 (
            .O(N__5860),
            .I(N__5846));
    LocalMux I__1381 (
            .O(N__5857),
            .I(N__5843));
    LocalMux I__1380 (
            .O(N__5854),
            .I(N__5838));
    LocalMux I__1379 (
            .O(N__5851),
            .I(N__5838));
    InMux I__1378 (
            .O(N__5850),
            .I(N__5835));
    CascadeMux I__1377 (
            .O(N__5849),
            .I(N__5832));
    Span4Mux_v I__1376 (
            .O(N__5846),
            .I(N__5828));
    Span4Mux_v I__1375 (
            .O(N__5843),
            .I(N__5825));
    Span4Mux_h I__1374 (
            .O(N__5838),
            .I(N__5822));
    LocalMux I__1373 (
            .O(N__5835),
            .I(N__5819));
    InMux I__1372 (
            .O(N__5832),
            .I(N__5814));
    InMux I__1371 (
            .O(N__5831),
            .I(N__5814));
    Sp12to4 I__1370 (
            .O(N__5828),
            .I(N__5811));
    Sp12to4 I__1369 (
            .O(N__5825),
            .I(N__5806));
    Sp12to4 I__1368 (
            .O(N__5822),
            .I(N__5806));
    Span4Mux_h I__1367 (
            .O(N__5819),
            .I(N__5801));
    LocalMux I__1366 (
            .O(N__5814),
            .I(N__5801));
    Span12Mux_h I__1365 (
            .O(N__5811),
            .I(N__5796));
    Span12Mux_v I__1364 (
            .O(N__5806),
            .I(N__5796));
    Span4Mux_v I__1363 (
            .O(N__5801),
            .I(N__5793));
    Odrv12 I__1362 (
            .O(N__5796),
            .I(LBENn_c));
    Odrv4 I__1361 (
            .O(N__5793),
            .I(LBENn_c));
    IoInMux I__1360 (
            .O(N__5788),
            .I(N__5785));
    LocalMux I__1359 (
            .O(N__5785),
            .I(N__5782));
    Span4Mux_s2_v I__1358 (
            .O(N__5782),
            .I(N__5779));
    Span4Mux_v I__1357 (
            .O(N__5779),
            .I(N__5776));
    Span4Mux_v I__1356 (
            .O(N__5776),
            .I(N__5773));
    Odrv4 I__1355 (
            .O(N__5773),
            .I(TAn_1_i));
    InMux I__1354 (
            .O(N__5770),
            .I(N__5767));
    LocalMux I__1353 (
            .O(N__5767),
            .I(N__5763));
    InMux I__1352 (
            .O(N__5766),
            .I(N__5760));
    Span4Mux_h I__1351 (
            .O(N__5763),
            .I(N__5757));
    LocalMux I__1350 (
            .O(N__5760),
            .I(N__5754));
    Sp12to4 I__1349 (
            .O(N__5757),
            .I(N__5750));
    Span4Mux_v I__1348 (
            .O(N__5754),
            .I(N__5747));
    InMux I__1347 (
            .O(N__5753),
            .I(N__5744));
    Span12Mux_v I__1346 (
            .O(N__5750),
            .I(N__5741));
    Sp12to4 I__1345 (
            .O(N__5747),
            .I(N__5736));
    LocalMux I__1344 (
            .O(N__5744),
            .I(N__5736));
    Span12Mux_h I__1343 (
            .O(N__5741),
            .I(N__5733));
    Span12Mux_h I__1342 (
            .O(N__5736),
            .I(N__5730));
    Odrv12 I__1341 (
            .O(N__5733),
            .I(D_UM_AMIGA_in_1));
    Odrv12 I__1340 (
            .O(N__5730),
            .I(D_UM_AMIGA_in_1));
    InMux I__1339 (
            .O(N__5725),
            .I(N__5722));
    LocalMux I__1338 (
            .O(N__5722),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ));
    IoInMux I__1337 (
            .O(N__5719),
            .I(N__5716));
    LocalMux I__1336 (
            .O(N__5716),
            .I(N__5713));
    Span4Mux_s3_h I__1335 (
            .O(N__5713),
            .I(N__5710));
    Sp12to4 I__1334 (
            .O(N__5710),
            .I(N__5707));
    Span12Mux_s10_v I__1333 (
            .O(N__5707),
            .I(N__5704));
    Odrv12 I__1332 (
            .O(N__5704),
            .I(un1_D_UM_AMIGA_1));
    InMux I__1331 (
            .O(N__5701),
            .I(N__5698));
    LocalMux I__1330 (
            .O(N__5698),
            .I(N__5695));
    Sp12to4 I__1329 (
            .O(N__5695),
            .I(N__5692));
    Odrv12 I__1328 (
            .O(N__5692),
            .I(TS_CPUn_c));
    InMux I__1327 (
            .O(N__5689),
            .I(N__5683));
    InMux I__1326 (
            .O(N__5688),
            .I(N__5680));
    InMux I__1325 (
            .O(N__5687),
            .I(N__5677));
    InMux I__1324 (
            .O(N__5686),
            .I(N__5674));
    LocalMux I__1323 (
            .O(N__5683),
            .I(N__5670));
    LocalMux I__1322 (
            .O(N__5680),
            .I(N__5667));
    LocalMux I__1321 (
            .O(N__5677),
            .I(N__5664));
    LocalMux I__1320 (
            .O(N__5674),
            .I(N__5661));
    ClkMux I__1319 (
            .O(N__5673),
            .I(N__5650));
    Glb2LocalMux I__1318 (
            .O(N__5670),
            .I(N__5650));
    Glb2LocalMux I__1317 (
            .O(N__5667),
            .I(N__5650));
    Glb2LocalMux I__1316 (
            .O(N__5664),
            .I(N__5650));
    Glb2LocalMux I__1315 (
            .O(N__5661),
            .I(N__5650));
    GlobalMux I__1314 (
            .O(N__5650),
            .I(CLK40));
    InMux I__1313 (
            .O(N__5647),
            .I(N__5644));
    LocalMux I__1312 (
            .O(N__5644),
            .I(N__5641));
    Span4Mux_v I__1311 (
            .O(N__5641),
            .I(N__5638));
    Odrv4 I__1310 (
            .O(N__5638),
            .I(\U111_CYCLE_SM.TS_EN_2_0 ));
    InMux I__1309 (
            .O(N__5635),
            .I(N__5632));
    LocalMux I__1308 (
            .O(N__5632),
            .I(N__5629));
    Odrv12 I__1307 (
            .O(N__5629),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ));
    InMux I__1306 (
            .O(N__5626),
            .I(N__5622));
    InMux I__1305 (
            .O(N__5625),
            .I(N__5618));
    LocalMux I__1304 (
            .O(N__5622),
            .I(N__5615));
    InMux I__1303 (
            .O(N__5621),
            .I(N__5612));
    LocalMux I__1302 (
            .O(N__5618),
            .I(N__5609));
    Span4Mux_v I__1301 (
            .O(N__5615),
            .I(N__5606));
    LocalMux I__1300 (
            .O(N__5612),
            .I(N__5603));
    Span4Mux_v I__1299 (
            .O(N__5609),
            .I(N__5600));
    Span4Mux_h I__1298 (
            .O(N__5606),
            .I(N__5597));
    Span12Mux_h I__1297 (
            .O(N__5603),
            .I(N__5594));
    Sp12to4 I__1296 (
            .O(N__5600),
            .I(N__5589));
    Sp12to4 I__1295 (
            .O(N__5597),
            .I(N__5589));
    Span12Mux_h I__1294 (
            .O(N__5594),
            .I(N__5586));
    Span12Mux_h I__1293 (
            .O(N__5589),
            .I(N__5583));
    Odrv12 I__1292 (
            .O(N__5586),
            .I(D_UU_AMIGA_in_7));
    Odrv12 I__1291 (
            .O(N__5583),
            .I(D_UU_AMIGA_in_7));
    IoInMux I__1290 (
            .O(N__5578),
            .I(N__5575));
    LocalMux I__1289 (
            .O(N__5575),
            .I(N__5572));
    Span4Mux_s0_v I__1288 (
            .O(N__5572),
            .I(N__5569));
    Span4Mux_v I__1287 (
            .O(N__5569),
            .I(N__5566));
    Span4Mux_v I__1286 (
            .O(N__5566),
            .I(N__5563));
    Sp12to4 I__1285 (
            .O(N__5563),
            .I(N__5560));
    Odrv12 I__1284 (
            .O(N__5560),
            .I(un1_D_UU_AMIGA_7));
    InMux I__1283 (
            .O(N__5557),
            .I(N__5554));
    LocalMux I__1282 (
            .O(N__5554),
            .I(N__5551));
    Odrv12 I__1281 (
            .O(N__5551),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ));
    InMux I__1280 (
            .O(N__5548),
            .I(N__5544));
    InMux I__1279 (
            .O(N__5547),
            .I(N__5540));
    LocalMux I__1278 (
            .O(N__5544),
            .I(N__5537));
    InMux I__1277 (
            .O(N__5543),
            .I(N__5534));
    LocalMux I__1276 (
            .O(N__5540),
            .I(N__5531));
    Span4Mux_v I__1275 (
            .O(N__5537),
            .I(N__5528));
    LocalMux I__1274 (
            .O(N__5534),
            .I(N__5525));
    Sp12to4 I__1273 (
            .O(N__5531),
            .I(N__5518));
    Sp12to4 I__1272 (
            .O(N__5528),
            .I(N__5518));
    Span12Mux_s11_v I__1271 (
            .O(N__5525),
            .I(N__5518));
    Span12Mux_h I__1270 (
            .O(N__5518),
            .I(N__5515));
    Odrv12 I__1269 (
            .O(N__5515),
            .I(D_UU_AMIGA_in_2));
    IoInMux I__1268 (
            .O(N__5512),
            .I(N__5509));
    LocalMux I__1267 (
            .O(N__5509),
            .I(N__5506));
    Span12Mux_s8_v I__1266 (
            .O(N__5506),
            .I(N__5503));
    Odrv12 I__1265 (
            .O(N__5503),
            .I(un1_D_UU_AMIGA_2));
    IoInMux I__1264 (
            .O(N__5500),
            .I(N__5497));
    LocalMux I__1263 (
            .O(N__5497),
            .I(N__5494));
    IoSpan4Mux I__1262 (
            .O(N__5494),
            .I(N__5491));
    Span4Mux_s3_h I__1261 (
            .O(N__5491),
            .I(N__5488));
    Span4Mux_h I__1260 (
            .O(N__5488),
            .I(N__5485));
    Span4Mux_h I__1259 (
            .O(N__5485),
            .I(N__5482));
    Odrv4 I__1258 (
            .O(N__5482),
            .I(un1_D_UM_AMIGA_0));
    InMux I__1257 (
            .O(N__5479),
            .I(N__5473));
    InMux I__1256 (
            .O(N__5478),
            .I(N__5473));
    LocalMux I__1255 (
            .O(N__5473),
            .I(N__5470));
    Span12Mux_v I__1254 (
            .O(N__5470),
            .I(N__5467));
    Span12Mux_h I__1253 (
            .O(N__5467),
            .I(N__5464));
    Odrv12 I__1252 (
            .O(N__5464),
            .I(BGn_c));
    IoInMux I__1251 (
            .O(N__5461),
            .I(N__5458));
    LocalMux I__1250 (
            .O(N__5458),
            .I(N__5453));
    IoInMux I__1249 (
            .O(N__5457),
            .I(N__5449));
    IoInMux I__1248 (
            .O(N__5456),
            .I(N__5446));
    Span4Mux_s2_h I__1247 (
            .O(N__5453),
            .I(N__5443));
    IoInMux I__1246 (
            .O(N__5452),
            .I(N__5440));
    LocalMux I__1245 (
            .O(N__5449),
            .I(N__5430));
    LocalMux I__1244 (
            .O(N__5446),
            .I(N__5430));
    IoSpan4Mux I__1243 (
            .O(N__5443),
            .I(N__5430));
    LocalMux I__1242 (
            .O(N__5440),
            .I(N__5430));
    IoInMux I__1241 (
            .O(N__5439),
            .I(N__5427));
    IoSpan4Mux I__1240 (
            .O(N__5430),
            .I(N__5411));
    LocalMux I__1239 (
            .O(N__5427),
            .I(N__5411));
    IoInMux I__1238 (
            .O(N__5426),
            .I(N__5408));
    IoInMux I__1237 (
            .O(N__5425),
            .I(N__5405));
    IoInMux I__1236 (
            .O(N__5424),
            .I(N__5402));
    IoInMux I__1235 (
            .O(N__5423),
            .I(N__5399));
    IoInMux I__1234 (
            .O(N__5422),
            .I(N__5396));
    IoInMux I__1233 (
            .O(N__5421),
            .I(N__5393));
    IoInMux I__1232 (
            .O(N__5420),
            .I(N__5389));
    IoInMux I__1231 (
            .O(N__5419),
            .I(N__5386));
    IoInMux I__1230 (
            .O(N__5418),
            .I(N__5378));
    IoInMux I__1229 (
            .O(N__5417),
            .I(N__5375));
    IoInMux I__1228 (
            .O(N__5416),
            .I(N__5372));
    IoSpan4Mux I__1227 (
            .O(N__5411),
            .I(N__5357));
    LocalMux I__1226 (
            .O(N__5408),
            .I(N__5357));
    LocalMux I__1225 (
            .O(N__5405),
            .I(N__5357));
    LocalMux I__1224 (
            .O(N__5402),
            .I(N__5357));
    LocalMux I__1223 (
            .O(N__5399),
            .I(N__5357));
    LocalMux I__1222 (
            .O(N__5396),
            .I(N__5357));
    LocalMux I__1221 (
            .O(N__5393),
            .I(N__5357));
    IoInMux I__1220 (
            .O(N__5392),
            .I(N__5354));
    LocalMux I__1219 (
            .O(N__5389),
            .I(N__5347));
    LocalMux I__1218 (
            .O(N__5386),
            .I(N__5347));
    IoInMux I__1217 (
            .O(N__5385),
            .I(N__5344));
    IoInMux I__1216 (
            .O(N__5384),
            .I(N__5341));
    IoInMux I__1215 (
            .O(N__5383),
            .I(N__5338));
    IoInMux I__1214 (
            .O(N__5382),
            .I(N__5335));
    IoInMux I__1213 (
            .O(N__5381),
            .I(N__5332));
    LocalMux I__1212 (
            .O(N__5378),
            .I(N__5323));
    LocalMux I__1211 (
            .O(N__5375),
            .I(N__5323));
    LocalMux I__1210 (
            .O(N__5372),
            .I(N__5323));
    IoSpan4Mux I__1209 (
            .O(N__5357),
            .I(N__5317));
    LocalMux I__1208 (
            .O(N__5354),
            .I(N__5317));
    IoInMux I__1207 (
            .O(N__5353),
            .I(N__5314));
    IoInMux I__1206 (
            .O(N__5352),
            .I(N__5310));
    IoSpan4Mux I__1205 (
            .O(N__5347),
            .I(N__5299));
    LocalMux I__1204 (
            .O(N__5344),
            .I(N__5299));
    LocalMux I__1203 (
            .O(N__5341),
            .I(N__5299));
    LocalMux I__1202 (
            .O(N__5338),
            .I(N__5299));
    LocalMux I__1201 (
            .O(N__5335),
            .I(N__5299));
    LocalMux I__1200 (
            .O(N__5332),
            .I(N__5296));
    IoInMux I__1199 (
            .O(N__5331),
            .I(N__5293));
    IoInMux I__1198 (
            .O(N__5330),
            .I(N__5290));
    IoSpan4Mux I__1197 (
            .O(N__5323),
            .I(N__5287));
    IoInMux I__1196 (
            .O(N__5322),
            .I(N__5284));
    IoSpan4Mux I__1195 (
            .O(N__5317),
            .I(N__5279));
    LocalMux I__1194 (
            .O(N__5314),
            .I(N__5279));
    IoInMux I__1193 (
            .O(N__5313),
            .I(N__5276));
    LocalMux I__1192 (
            .O(N__5310),
            .I(N__5271));
    IoSpan4Mux I__1191 (
            .O(N__5299),
            .I(N__5268));
    Span4Mux_s3_v I__1190 (
            .O(N__5296),
            .I(N__5265));
    LocalMux I__1189 (
            .O(N__5293),
            .I(N__5259));
    LocalMux I__1188 (
            .O(N__5290),
            .I(N__5259));
    IoSpan4Mux I__1187 (
            .O(N__5287),
            .I(N__5254));
    LocalMux I__1186 (
            .O(N__5284),
            .I(N__5254));
    IoSpan4Mux I__1185 (
            .O(N__5279),
            .I(N__5249));
    LocalMux I__1184 (
            .O(N__5276),
            .I(N__5249));
    IoInMux I__1183 (
            .O(N__5275),
            .I(N__5246));
    IoInMux I__1182 (
            .O(N__5274),
            .I(N__5243));
    Span4Mux_s2_h I__1181 (
            .O(N__5271),
            .I(N__5236));
    Span4Mux_s3_v I__1180 (
            .O(N__5268),
            .I(N__5236));
    Span4Mux_h I__1179 (
            .O(N__5265),
            .I(N__5236));
    IoInMux I__1178 (
            .O(N__5264),
            .I(N__5233));
    Span4Mux_s3_h I__1177 (
            .O(N__5259),
            .I(N__5230));
    IoSpan4Mux I__1176 (
            .O(N__5254),
            .I(N__5225));
    IoSpan4Mux I__1175 (
            .O(N__5249),
            .I(N__5225));
    LocalMux I__1174 (
            .O(N__5246),
            .I(N__5217));
    LocalMux I__1173 (
            .O(N__5243),
            .I(N__5217));
    Sp12to4 I__1172 (
            .O(N__5236),
            .I(N__5217));
    LocalMux I__1171 (
            .O(N__5233),
            .I(N__5214));
    Span4Mux_v I__1170 (
            .O(N__5230),
            .I(N__5209));
    Span4Mux_s3_h I__1169 (
            .O(N__5225),
            .I(N__5209));
    IoInMux I__1168 (
            .O(N__5224),
            .I(N__5206));
    Span12Mux_s11_v I__1167 (
            .O(N__5217),
            .I(N__5201));
    Span12Mux_s2_h I__1166 (
            .O(N__5214),
            .I(N__5201));
    Sp12to4 I__1165 (
            .O(N__5209),
            .I(N__5196));
    LocalMux I__1164 (
            .O(N__5206),
            .I(N__5196));
    Span12Mux_h I__1163 (
            .O(N__5201),
            .I(N__5193));
    Span12Mux_s8_h I__1162 (
            .O(N__5196),
            .I(N__5190));
    Odrv12 I__1161 (
            .O(N__5193),
            .I(CPU_READ_EN_i));
    Odrv12 I__1160 (
            .O(N__5190),
            .I(CPU_READ_EN_i));
    CascadeMux I__1159 (
            .O(N__5185),
            .I(\U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0_cascade_ ));
    CascadeMux I__1158 (
            .O(N__5182),
            .I(N__5177));
    InMux I__1157 (
            .O(N__5181),
            .I(N__5172));
    InMux I__1156 (
            .O(N__5180),
            .I(N__5167));
    InMux I__1155 (
            .O(N__5177),
            .I(N__5167));
    InMux I__1154 (
            .O(N__5176),
            .I(N__5162));
    InMux I__1153 (
            .O(N__5175),
            .I(N__5162));
    LocalMux I__1152 (
            .O(N__5172),
            .I(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ));
    LocalMux I__1151 (
            .O(N__5167),
            .I(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ));
    LocalMux I__1150 (
            .O(N__5162),
            .I(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ));
    CascadeMux I__1149 (
            .O(N__5155),
            .I(\U111_CYCLE_SM.N_97_cascade_ ));
    InMux I__1148 (
            .O(N__5152),
            .I(N__5149));
    LocalMux I__1147 (
            .O(N__5149),
            .I(\U111_CYCLE_SM.LW_CYCLE_0 ));
    InMux I__1146 (
            .O(N__5146),
            .I(N__5143));
    LocalMux I__1145 (
            .O(N__5143),
            .I(N__5140));
    Span12Mux_h I__1144 (
            .O(N__5140),
            .I(N__5135));
    InMux I__1143 (
            .O(N__5139),
            .I(N__5130));
    InMux I__1142 (
            .O(N__5138),
            .I(N__5130));
    Span12Mux_v I__1141 (
            .O(N__5135),
            .I(N__5127));
    LocalMux I__1140 (
            .O(N__5130),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    Odrv12 I__1139 (
            .O(N__5127),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    InMux I__1138 (
            .O(N__5122),
            .I(N__5119));
    LocalMux I__1137 (
            .O(N__5119),
            .I(\U111_CYCLE_SM.un3_LW_CYCLE_START ));
    SRMux I__1136 (
            .O(N__5116),
            .I(N__5113));
    LocalMux I__1135 (
            .O(N__5113),
            .I(N__5110));
    Span4Mux_h I__1134 (
            .O(N__5110),
            .I(N__5107));
    Odrv4 I__1133 (
            .O(N__5107),
            .I(\U111_CYCLE_SM.RESETn_c_i ));
    InMux I__1132 (
            .O(N__5104),
            .I(N__5101));
    LocalMux I__1131 (
            .O(N__5101),
            .I(N__5098));
    Span4Mux_v I__1130 (
            .O(N__5098),
            .I(N__5095));
    Sp12to4 I__1129 (
            .O(N__5095),
            .I(N__5092));
    Span12Mux_h I__1128 (
            .O(N__5092),
            .I(N__5089));
    Odrv12 I__1127 (
            .O(N__5089),
            .I(SIZ_c_1));
    InMux I__1126 (
            .O(N__5086),
            .I(N__5083));
    LocalMux I__1125 (
            .O(N__5083),
            .I(N__5080));
    Span4Mux_v I__1124 (
            .O(N__5080),
            .I(N__5077));
    Sp12to4 I__1123 (
            .O(N__5077),
            .I(N__5074));
    Span12Mux_h I__1122 (
            .O(N__5074),
            .I(N__5071));
    Odrv12 I__1121 (
            .O(N__5071),
            .I(SIZ_c_0));
    InMux I__1120 (
            .O(N__5068),
            .I(N__5065));
    LocalMux I__1119 (
            .O(N__5065),
            .I(N__5061));
    InMux I__1118 (
            .O(N__5064),
            .I(N__5058));
    Span4Mux_v I__1117 (
            .O(N__5061),
            .I(N__5053));
    LocalMux I__1116 (
            .O(N__5058),
            .I(N__5053));
    Span4Mux_v I__1115 (
            .O(N__5053),
            .I(N__5050));
    Sp12to4 I__1114 (
            .O(N__5050),
            .I(N__5047));
    Span12Mux_h I__1113 (
            .O(N__5047),
            .I(N__5044));
    Span12Mux_v I__1112 (
            .O(N__5044),
            .I(N__5041));
    Odrv12 I__1111 (
            .O(N__5041),
            .I(PORTSIZE_c));
    InMux I__1110 (
            .O(N__5038),
            .I(N__5034));
    InMux I__1109 (
            .O(N__5037),
            .I(N__5031));
    LocalMux I__1108 (
            .O(N__5034),
            .I(N__5028));
    LocalMux I__1107 (
            .O(N__5031),
            .I(N__5025));
    Odrv12 I__1106 (
            .O(N__5028),
            .I(\U111_CYCLE_SM.LW_TRANS_0 ));
    Odrv12 I__1105 (
            .O(N__5025),
            .I(\U111_CYCLE_SM.LW_TRANS_0 ));
    InMux I__1104 (
            .O(N__5020),
            .I(N__5017));
    LocalMux I__1103 (
            .O(N__5017),
            .I(N__5014));
    Span4Mux_v I__1102 (
            .O(N__5014),
            .I(N__5011));
    Sp12to4 I__1101 (
            .O(N__5011),
            .I(N__5008));
    Span12Mux_h I__1100 (
            .O(N__5008),
            .I(N__5005));
    Odrv12 I__1099 (
            .O(N__5005),
            .I(D_LM_AMIGA_in_7));
    IoInMux I__1098 (
            .O(N__5002),
            .I(N__4999));
    LocalMux I__1097 (
            .O(N__4999),
            .I(N__4996));
    IoSpan4Mux I__1096 (
            .O(N__4996),
            .I(N__4993));
    Span4Mux_s2_h I__1095 (
            .O(N__4993),
            .I(N__4990));
    Sp12to4 I__1094 (
            .O(N__4990),
            .I(N__4987));
    Odrv12 I__1093 (
            .O(N__4987),
            .I(un1_D_LM_AMIGA_7));
    IoInMux I__1092 (
            .O(N__4984),
            .I(N__4981));
    LocalMux I__1091 (
            .O(N__4981),
            .I(N__4977));
    InMux I__1090 (
            .O(N__4980),
            .I(N__4974));
    IoSpan4Mux I__1089 (
            .O(N__4977),
            .I(N__4971));
    LocalMux I__1088 (
            .O(N__4974),
            .I(N__4968));
    Span4Mux_s3_h I__1087 (
            .O(N__4971),
            .I(N__4965));
    Span4Mux_h I__1086 (
            .O(N__4968),
            .I(N__4962));
    Sp12to4 I__1085 (
            .O(N__4965),
            .I(N__4959));
    Sp12to4 I__1084 (
            .O(N__4962),
            .I(N__4956));
    Span12Mux_v I__1083 (
            .O(N__4959),
            .I(N__4953));
    Span12Mux_v I__1082 (
            .O(N__4956),
            .I(N__4950));
    Span12Mux_h I__1081 (
            .O(N__4953),
            .I(N__4947));
    Span12Mux_v I__1080 (
            .O(N__4950),
            .I(N__4944));
    Span12Mux_h I__1079 (
            .O(N__4947),
            .I(N__4941));
    Span12Mux_h I__1078 (
            .O(N__4944),
            .I(N__4938));
    Odrv12 I__1077 (
            .O(N__4941),
            .I(D_LL_040_in_5));
    Odrv12 I__1076 (
            .O(N__4938),
            .I(D_LL_040_in_5));
    InMux I__1075 (
            .O(N__4933),
            .I(N__4930));
    LocalMux I__1074 (
            .O(N__4930),
            .I(N__4927));
    Span4Mux_v I__1073 (
            .O(N__4927),
            .I(N__4924));
    Sp12to4 I__1072 (
            .O(N__4924),
            .I(N__4921));
    Span12Mux_h I__1071 (
            .O(N__4921),
            .I(N__4918));
    Odrv12 I__1070 (
            .O(N__4918),
            .I(D_UM_040_in_5));
    IoInMux I__1069 (
            .O(N__4915),
            .I(N__4912));
    LocalMux I__1068 (
            .O(N__4912),
            .I(N__4909));
    Span12Mux_s10_v I__1067 (
            .O(N__4909),
            .I(N__4906));
    Span12Mux_h I__1066 (
            .O(N__4906),
            .I(N__4903));
    Odrv12 I__1065 (
            .O(N__4903),
            .I(un1_D_UM_040_5));
    InMux I__1064 (
            .O(N__4900),
            .I(N__4897));
    LocalMux I__1063 (
            .O(N__4897),
            .I(N__4894));
    Span4Mux_v I__1062 (
            .O(N__4894),
            .I(N__4891));
    Sp12to4 I__1061 (
            .O(N__4891),
            .I(N__4888));
    Span12Mux_h I__1060 (
            .O(N__4888),
            .I(N__4885));
    Odrv12 I__1059 (
            .O(N__4885),
            .I(D_UU_040_in_3));
    InMux I__1058 (
            .O(N__4882),
            .I(N__4875));
    InMux I__1057 (
            .O(N__4881),
            .I(N__4872));
    InMux I__1056 (
            .O(N__4880),
            .I(N__4864));
    InMux I__1055 (
            .O(N__4879),
            .I(N__4864));
    InMux I__1054 (
            .O(N__4878),
            .I(N__4861));
    LocalMux I__1053 (
            .O(N__4875),
            .I(N__4850));
    LocalMux I__1052 (
            .O(N__4872),
            .I(N__4850));
    InMux I__1051 (
            .O(N__4871),
            .I(N__4847));
    InMux I__1050 (
            .O(N__4870),
            .I(N__4844));
    InMux I__1049 (
            .O(N__4869),
            .I(N__4841));
    LocalMux I__1048 (
            .O(N__4864),
            .I(N__4836));
    LocalMux I__1047 (
            .O(N__4861),
            .I(N__4836));
    InMux I__1046 (
            .O(N__4860),
            .I(N__4831));
    InMux I__1045 (
            .O(N__4859),
            .I(N__4831));
    InMux I__1044 (
            .O(N__4858),
            .I(N__4824));
    InMux I__1043 (
            .O(N__4857),
            .I(N__4824));
    InMux I__1042 (
            .O(N__4856),
            .I(N__4821));
    InMux I__1041 (
            .O(N__4855),
            .I(N__4809));
    Span4Mux_v I__1040 (
            .O(N__4850),
            .I(N__4800));
    LocalMux I__1039 (
            .O(N__4847),
            .I(N__4800));
    LocalMux I__1038 (
            .O(N__4844),
            .I(N__4800));
    LocalMux I__1037 (
            .O(N__4841),
            .I(N__4797));
    Span4Mux_v I__1036 (
            .O(N__4836),
            .I(N__4792));
    LocalMux I__1035 (
            .O(N__4831),
            .I(N__4792));
    InMux I__1034 (
            .O(N__4830),
            .I(N__4789));
    InMux I__1033 (
            .O(N__4829),
            .I(N__4786));
    LocalMux I__1032 (
            .O(N__4824),
            .I(N__4781));
    LocalMux I__1031 (
            .O(N__4821),
            .I(N__4781));
    InMux I__1030 (
            .O(N__4820),
            .I(N__4778));
    InMux I__1029 (
            .O(N__4819),
            .I(N__4775));
    InMux I__1028 (
            .O(N__4818),
            .I(N__4770));
    InMux I__1027 (
            .O(N__4817),
            .I(N__4770));
    InMux I__1026 (
            .O(N__4816),
            .I(N__4765));
    InMux I__1025 (
            .O(N__4815),
            .I(N__4765));
    InMux I__1024 (
            .O(N__4814),
            .I(N__4762));
    InMux I__1023 (
            .O(N__4813),
            .I(N__4754));
    InMux I__1022 (
            .O(N__4812),
            .I(N__4754));
    LocalMux I__1021 (
            .O(N__4809),
            .I(N__4751));
    InMux I__1020 (
            .O(N__4808),
            .I(N__4746));
    InMux I__1019 (
            .O(N__4807),
            .I(N__4746));
    Span4Mux_v I__1018 (
            .O(N__4800),
            .I(N__4743));
    Span4Mux_v I__1017 (
            .O(N__4797),
            .I(N__4734));
    Span4Mux_v I__1016 (
            .O(N__4792),
            .I(N__4734));
    LocalMux I__1015 (
            .O(N__4789),
            .I(N__4734));
    LocalMux I__1014 (
            .O(N__4786),
            .I(N__4734));
    Span4Mux_v I__1013 (
            .O(N__4781),
            .I(N__4729));
    LocalMux I__1012 (
            .O(N__4778),
            .I(N__4729));
    LocalMux I__1011 (
            .O(N__4775),
            .I(N__4726));
    LocalMux I__1010 (
            .O(N__4770),
            .I(N__4723));
    LocalMux I__1009 (
            .O(N__4765),
            .I(N__4720));
    LocalMux I__1008 (
            .O(N__4762),
            .I(N__4717));
    InMux I__1007 (
            .O(N__4761),
            .I(N__4712));
    InMux I__1006 (
            .O(N__4760),
            .I(N__4712));
    InMux I__1005 (
            .O(N__4759),
            .I(N__4709));
    LocalMux I__1004 (
            .O(N__4754),
            .I(N__4705));
    Span12Mux_h I__1003 (
            .O(N__4751),
            .I(N__4700));
    LocalMux I__1002 (
            .O(N__4746),
            .I(N__4700));
    Span4Mux_v I__1001 (
            .O(N__4743),
            .I(N__4697));
    Span4Mux_v I__1000 (
            .O(N__4734),
            .I(N__4694));
    Span4Mux_v I__999 (
            .O(N__4729),
            .I(N__4687));
    Span4Mux_v I__998 (
            .O(N__4726),
            .I(N__4687));
    Span4Mux_h I__997 (
            .O(N__4723),
            .I(N__4687));
    Span4Mux_v I__996 (
            .O(N__4720),
            .I(N__4680));
    Span4Mux_h I__995 (
            .O(N__4717),
            .I(N__4680));
    LocalMux I__994 (
            .O(N__4712),
            .I(N__4680));
    LocalMux I__993 (
            .O(N__4709),
            .I(N__4677));
    InMux I__992 (
            .O(N__4708),
            .I(N__4674));
    Odrv12 I__991 (
            .O(N__4705),
            .I(\U111_CYCLE_SM.FLIP ));
    Odrv12 I__990 (
            .O(N__4700),
            .I(\U111_CYCLE_SM.FLIP ));
    Odrv4 I__989 (
            .O(N__4697),
            .I(\U111_CYCLE_SM.FLIP ));
    Odrv4 I__988 (
            .O(N__4694),
            .I(\U111_CYCLE_SM.FLIP ));
    Odrv4 I__987 (
            .O(N__4687),
            .I(\U111_CYCLE_SM.FLIP ));
    Odrv4 I__986 (
            .O(N__4680),
            .I(\U111_CYCLE_SM.FLIP ));
    Odrv12 I__985 (
            .O(N__4677),
            .I(\U111_CYCLE_SM.FLIP ));
    LocalMux I__984 (
            .O(N__4674),
            .I(\U111_CYCLE_SM.FLIP ));
    IoInMux I__983 (
            .O(N__4657),
            .I(N__4654));
    LocalMux I__982 (
            .O(N__4654),
            .I(N__4651));
    IoSpan4Mux I__981 (
            .O(N__4651),
            .I(N__4647));
    InMux I__980 (
            .O(N__4650),
            .I(N__4644));
    IoSpan4Mux I__979 (
            .O(N__4647),
            .I(N__4641));
    LocalMux I__978 (
            .O(N__4644),
            .I(N__4638));
    Span4Mux_s2_h I__977 (
            .O(N__4641),
            .I(N__4635));
    Span4Mux_v I__976 (
            .O(N__4638),
            .I(N__4632));
    Sp12to4 I__975 (
            .O(N__4635),
            .I(N__4629));
    Sp12to4 I__974 (
            .O(N__4632),
            .I(N__4626));
    Span12Mux_h I__973 (
            .O(N__4629),
            .I(N__4623));
    Span12Mux_v I__972 (
            .O(N__4626),
            .I(N__4620));
    Span12Mux_h I__971 (
            .O(N__4623),
            .I(N__4617));
    Span12Mux_h I__970 (
            .O(N__4620),
            .I(N__4614));
    Odrv12 I__969 (
            .O(N__4617),
            .I(D_LM_040_in_3));
    Odrv12 I__968 (
            .O(N__4614),
            .I(D_LM_040_in_3));
    IoInMux I__967 (
            .O(N__4609),
            .I(N__4606));
    LocalMux I__966 (
            .O(N__4606),
            .I(N__4603));
    IoSpan4Mux I__965 (
            .O(N__4603),
            .I(N__4600));
    IoSpan4Mux I__964 (
            .O(N__4600),
            .I(N__4597));
    Span4Mux_s2_v I__963 (
            .O(N__4597),
            .I(N__4594));
    Span4Mux_h I__962 (
            .O(N__4594),
            .I(N__4591));
    Span4Mux_v I__961 (
            .O(N__4591),
            .I(N__4588));
    Odrv4 I__960 (
            .O(N__4588),
            .I(un1_D_UU_040_3));
    IoInMux I__959 (
            .O(N__4585),
            .I(N__4582));
    LocalMux I__958 (
            .O(N__4582),
            .I(N__4579));
    Span4Mux_s2_v I__957 (
            .O(N__4579),
            .I(N__4576));
    Span4Mux_v I__956 (
            .O(N__4576),
            .I(N__4573));
    Span4Mux_h I__955 (
            .O(N__4573),
            .I(N__4570));
    Span4Mux_h I__954 (
            .O(N__4570),
            .I(N__4567));
    Odrv4 I__953 (
            .O(N__4567),
            .I(U111_CYCLE_SM_TBI_CPUn_0_i));
    InMux I__952 (
            .O(N__4564),
            .I(N__4561));
    LocalMux I__951 (
            .O(N__4561),
            .I(\U111_CYCLE_SM.TS_EN_5 ));
    InMux I__950 (
            .O(N__4558),
            .I(N__4555));
    LocalMux I__949 (
            .O(N__4555),
            .I(N__4552));
    Span12Mux_h I__948 (
            .O(N__4552),
            .I(N__4549));
    Odrv12 I__947 (
            .O(N__4549),
            .I(D_LM_AMIGA_in_1));
    CascadeMux I__946 (
            .O(N__4546),
            .I(\U111_CYCLE_SM.FLIP_cascade_ ));
    IoInMux I__945 (
            .O(N__4543),
            .I(N__4540));
    LocalMux I__944 (
            .O(N__4540),
            .I(N__4537));
    Span4Mux_s3_h I__943 (
            .O(N__4537),
            .I(N__4534));
    Sp12to4 I__942 (
            .O(N__4534),
            .I(N__4531));
    Span12Mux_v I__941 (
            .O(N__4531),
            .I(N__4528));
    Odrv12 I__940 (
            .O(N__4528),
            .I(un1_D_LM_AMIGA_1));
    IoInMux I__939 (
            .O(N__4525),
            .I(N__4522));
    LocalMux I__938 (
            .O(N__4522),
            .I(N__4516));
    IoInMux I__937 (
            .O(N__4521),
            .I(N__4513));
    IoInMux I__936 (
            .O(N__4520),
            .I(N__4510));
    IoInMux I__935 (
            .O(N__4519),
            .I(N__4507));
    IoSpan4Mux I__934 (
            .O(N__4516),
            .I(N__4504));
    LocalMux I__933 (
            .O(N__4513),
            .I(N__4501));
    LocalMux I__932 (
            .O(N__4510),
            .I(N__4498));
    LocalMux I__931 (
            .O(N__4507),
            .I(N__4495));
    IoSpan4Mux I__930 (
            .O(N__4504),
            .I(N__4490));
    IoSpan4Mux I__929 (
            .O(N__4501),
            .I(N__4490));
    IoSpan4Mux I__928 (
            .O(N__4498),
            .I(N__4487));
    IoSpan4Mux I__927 (
            .O(N__4495),
            .I(N__4484));
    Span4Mux_s2_v I__926 (
            .O(N__4490),
            .I(N__4481));
    Sp12to4 I__925 (
            .O(N__4487),
            .I(N__4478));
    Sp12to4 I__924 (
            .O(N__4484),
            .I(N__4475));
    Sp12to4 I__923 (
            .O(N__4481),
            .I(N__4472));
    Span12Mux_h I__922 (
            .O(N__4478),
            .I(N__4467));
    Span12Mux_s7_h I__921 (
            .O(N__4475),
            .I(N__4467));
    Odrv12 I__920 (
            .O(N__4472),
            .I(GB_BUFFER_CLK40_THRU_CO));
    Odrv12 I__919 (
            .O(N__4467),
            .I(GB_BUFFER_CLK40_THRU_CO));
    InMux I__918 (
            .O(N__4462),
            .I(N__4459));
    LocalMux I__917 (
            .O(N__4459),
            .I(N__4455));
    ClkMux I__916 (
            .O(N__4458),
            .I(N__4429));
    Glb2LocalMux I__915 (
            .O(N__4455),
            .I(N__4429));
    ClkMux I__914 (
            .O(N__4454),
            .I(N__4429));
    ClkMux I__913 (
            .O(N__4453),
            .I(N__4429));
    ClkMux I__912 (
            .O(N__4452),
            .I(N__4429));
    ClkMux I__911 (
            .O(N__4451),
            .I(N__4429));
    ClkMux I__910 (
            .O(N__4450),
            .I(N__4429));
    ClkMux I__909 (
            .O(N__4449),
            .I(N__4429));
    ClkMux I__908 (
            .O(N__4448),
            .I(N__4429));
    GlobalMux I__907 (
            .O(N__4429),
            .I(CLK80));
    IoInMux I__906 (
            .O(N__4426),
            .I(N__4423));
    LocalMux I__905 (
            .O(N__4423),
            .I(N__4419));
    IoInMux I__904 (
            .O(N__4422),
            .I(N__4416));
    Span12Mux_s2_v I__903 (
            .O(N__4419),
            .I(N__4413));
    LocalMux I__902 (
            .O(N__4416),
            .I(N__4410));
    Span12Mux_v I__901 (
            .O(N__4413),
            .I(N__4407));
    Span12Mux_s9_h I__900 (
            .O(N__4410),
            .I(N__4404));
    Odrv12 I__899 (
            .O(N__4407),
            .I(GB_BUFFER_CLK80_THRU_CO));
    Odrv12 I__898 (
            .O(N__4404),
            .I(GB_BUFFER_CLK80_THRU_CO));
    CascadeMux I__897 (
            .O(N__4399),
            .I(\U111_CYCLE_SM.A_OUT_0_cascade_ ));
    InMux I__896 (
            .O(N__4396),
            .I(N__4393));
    LocalMux I__895 (
            .O(N__4393),
            .I(N__4390));
    Span12Mux_s10_h I__894 (
            .O(N__4390),
            .I(N__4387));
    Span12Mux_v I__893 (
            .O(N__4387),
            .I(N__4383));
    InMux I__892 (
            .O(N__4386),
            .I(N__4380));
    Odrv12 I__891 (
            .O(N__4383),
            .I(\U111_CYCLE_SM.A_OUTZ0 ));
    LocalMux I__890 (
            .O(N__4380),
            .I(\U111_CYCLE_SM.A_OUTZ0 ));
    CascadeMux I__889 (
            .O(N__4375),
            .I(\U111_CYCLE_SM.N_75_0_cascade_ ));
    IoInMux I__888 (
            .O(N__4372),
            .I(N__4369));
    LocalMux I__887 (
            .O(N__4369),
            .I(N__4366));
    Span4Mux_s3_h I__886 (
            .O(N__4366),
            .I(N__4363));
    Span4Mux_v I__885 (
            .O(N__4363),
            .I(N__4360));
    Sp12to4 I__884 (
            .O(N__4360),
            .I(N__4357));
    Span12Mux_h I__883 (
            .O(N__4357),
            .I(N__4354));
    Odrv12 I__882 (
            .O(N__4354),
            .I(un1_D_LM_AMIGA_0));
    InMux I__881 (
            .O(N__4351),
            .I(N__4348));
    LocalMux I__880 (
            .O(N__4348),
            .I(N__4345));
    Span12Mux_v I__879 (
            .O(N__4345),
            .I(N__4342));
    Span12Mux_h I__878 (
            .O(N__4342),
            .I(N__4339));
    Odrv12 I__877 (
            .O(N__4339),
            .I(D_LL_AMIGA_in_7));
    IoInMux I__876 (
            .O(N__4336),
            .I(N__4333));
    LocalMux I__875 (
            .O(N__4333),
            .I(N__4330));
    Span4Mux_s3_h I__874 (
            .O(N__4330),
            .I(N__4327));
    Span4Mux_v I__873 (
            .O(N__4327),
            .I(N__4324));
    Span4Mux_v I__872 (
            .O(N__4324),
            .I(N__4321));
    Sp12to4 I__871 (
            .O(N__4321),
            .I(N__4318));
    Odrv12 I__870 (
            .O(N__4318),
            .I(un1_D_LL_AMIGA_7));
    IoInMux I__869 (
            .O(N__4315),
            .I(N__4312));
    LocalMux I__868 (
            .O(N__4312),
            .I(N__4308));
    InMux I__867 (
            .O(N__4311),
            .I(N__4305));
    IoSpan4Mux I__866 (
            .O(N__4308),
            .I(N__4302));
    LocalMux I__865 (
            .O(N__4305),
            .I(N__4299));
    Span4Mux_s2_h I__864 (
            .O(N__4302),
            .I(N__4296));
    Span4Mux_v I__863 (
            .O(N__4299),
            .I(N__4293));
    Sp12to4 I__862 (
            .O(N__4296),
            .I(N__4290));
    Sp12to4 I__861 (
            .O(N__4293),
            .I(N__4287));
    Span12Mux_h I__860 (
            .O(N__4290),
            .I(N__4284));
    Span12Mux_h I__859 (
            .O(N__4287),
            .I(N__4281));
    Span12Mux_h I__858 (
            .O(N__4284),
            .I(N__4278));
    Span12Mux_v I__857 (
            .O(N__4281),
            .I(N__4275));
    Odrv12 I__856 (
            .O(N__4278),
            .I(D_LL_040_in_0));
    Odrv12 I__855 (
            .O(N__4275),
            .I(D_LL_040_in_0));
    InMux I__854 (
            .O(N__4270),
            .I(N__4267));
    LocalMux I__853 (
            .O(N__4267),
            .I(N__4264));
    Span12Mux_h I__852 (
            .O(N__4264),
            .I(N__4261));
    Odrv12 I__851 (
            .O(N__4261),
            .I(D_UM_040_in_0));
    IoInMux I__850 (
            .O(N__4258),
            .I(N__4255));
    LocalMux I__849 (
            .O(N__4255),
            .I(N__4252));
    IoSpan4Mux I__848 (
            .O(N__4252),
            .I(N__4249));
    Span4Mux_s0_h I__847 (
            .O(N__4249),
            .I(N__4246));
    Sp12to4 I__846 (
            .O(N__4246),
            .I(N__4243));
    Span12Mux_s11_h I__845 (
            .O(N__4243),
            .I(N__4240));
    Odrv12 I__844 (
            .O(N__4240),
            .I(un1_D_UM_040_0));
    InMux I__843 (
            .O(N__4237),
            .I(N__4234));
    LocalMux I__842 (
            .O(N__4234),
            .I(N__4231));
    Span4Mux_h I__841 (
            .O(N__4231),
            .I(N__4228));
    Sp12to4 I__840 (
            .O(N__4228),
            .I(N__4225));
    Span12Mux_v I__839 (
            .O(N__4225),
            .I(N__4222));
    Span12Mux_h I__838 (
            .O(N__4222),
            .I(N__4219));
    Odrv12 I__837 (
            .O(N__4219),
            .I(D_UM_040_in_4));
    InMux I__836 (
            .O(N__4216),
            .I(N__4212));
    IoInMux I__835 (
            .O(N__4215),
            .I(N__4209));
    LocalMux I__834 (
            .O(N__4212),
            .I(N__4206));
    LocalMux I__833 (
            .O(N__4209),
            .I(N__4203));
    Span4Mux_v I__832 (
            .O(N__4206),
            .I(N__4200));
    Span4Mux_s2_h I__831 (
            .O(N__4203),
            .I(N__4197));
    Sp12to4 I__830 (
            .O(N__4200),
            .I(N__4194));
    Span4Mux_v I__829 (
            .O(N__4197),
            .I(N__4191));
    Span12Mux_h I__828 (
            .O(N__4194),
            .I(N__4188));
    Sp12to4 I__827 (
            .O(N__4191),
            .I(N__4185));
    Span12Mux_v I__826 (
            .O(N__4188),
            .I(N__4182));
    Span12Mux_h I__825 (
            .O(N__4185),
            .I(N__4179));
    Span12Mux_v I__824 (
            .O(N__4182),
            .I(N__4176));
    Span12Mux_h I__823 (
            .O(N__4179),
            .I(N__4173));
    Odrv12 I__822 (
            .O(N__4176),
            .I(D_LL_040_in_4));
    Odrv12 I__821 (
            .O(N__4173),
            .I(D_LL_040_in_4));
    IoInMux I__820 (
            .O(N__4168),
            .I(N__4165));
    LocalMux I__819 (
            .O(N__4165),
            .I(N__4162));
    Span12Mux_s3_h I__818 (
            .O(N__4162),
            .I(N__4159));
    Span12Mux_h I__817 (
            .O(N__4159),
            .I(N__4156));
    Odrv12 I__816 (
            .O(N__4156),
            .I(un1_D_UM_040_4));
    IoInMux I__815 (
            .O(N__4153),
            .I(N__4150));
    LocalMux I__814 (
            .O(N__4150),
            .I(N__4147));
    IoSpan4Mux I__813 (
            .O(N__4147),
            .I(N__4143));
    InMux I__812 (
            .O(N__4146),
            .I(N__4140));
    Span4Mux_s0_h I__811 (
            .O(N__4143),
            .I(N__4137));
    LocalMux I__810 (
            .O(N__4140),
            .I(N__4134));
    Span4Mux_v I__809 (
            .O(N__4137),
            .I(N__4131));
    Span4Mux_v I__808 (
            .O(N__4134),
            .I(N__4128));
    Sp12to4 I__807 (
            .O(N__4131),
            .I(N__4125));
    Sp12to4 I__806 (
            .O(N__4128),
            .I(N__4122));
    Span12Mux_h I__805 (
            .O(N__4125),
            .I(N__4119));
    Span12Mux_h I__804 (
            .O(N__4122),
            .I(N__4116));
    Span12Mux_h I__803 (
            .O(N__4119),
            .I(N__4113));
    Span12Mux_v I__802 (
            .O(N__4116),
            .I(N__4110));
    Odrv12 I__801 (
            .O(N__4113),
            .I(D_LM_040_in_5));
    Odrv12 I__800 (
            .O(N__4110),
            .I(D_LM_040_in_5));
    InMux I__799 (
            .O(N__4105),
            .I(N__4102));
    LocalMux I__798 (
            .O(N__4102),
            .I(N__4099));
    Span4Mux_v I__797 (
            .O(N__4099),
            .I(N__4096));
    Span4Mux_v I__796 (
            .O(N__4096),
            .I(N__4093));
    Sp12to4 I__795 (
            .O(N__4093),
            .I(N__4090));
    Span12Mux_h I__794 (
            .O(N__4090),
            .I(N__4087));
    Odrv12 I__793 (
            .O(N__4087),
            .I(D_UU_040_in_5));
    IoInMux I__792 (
            .O(N__4084),
            .I(N__4081));
    LocalMux I__791 (
            .O(N__4081),
            .I(N__4078));
    Span4Mux_s3_h I__790 (
            .O(N__4078),
            .I(N__4075));
    Sp12to4 I__789 (
            .O(N__4075),
            .I(N__4072));
    Span12Mux_s10_v I__788 (
            .O(N__4072),
            .I(N__4069));
    Span12Mux_h I__787 (
            .O(N__4069),
            .I(N__4066));
    Odrv12 I__786 (
            .O(N__4066),
            .I(un1_D_UU_040_5));
    IoInMux I__785 (
            .O(N__4063),
            .I(N__4060));
    LocalMux I__784 (
            .O(N__4060),
            .I(N__4057));
    IoSpan4Mux I__783 (
            .O(N__4057),
            .I(N__4053));
    InMux I__782 (
            .O(N__4056),
            .I(N__4050));
    Span4Mux_s2_h I__781 (
            .O(N__4053),
            .I(N__4047));
    LocalMux I__780 (
            .O(N__4050),
            .I(N__4044));
    Sp12to4 I__779 (
            .O(N__4047),
            .I(N__4041));
    Span4Mux_v I__778 (
            .O(N__4044),
            .I(N__4038));
    Span12Mux_h I__777 (
            .O(N__4041),
            .I(N__4035));
    Span4Mux_h I__776 (
            .O(N__4038),
            .I(N__4032));
    Span12Mux_h I__775 (
            .O(N__4035),
            .I(N__4029));
    Sp12to4 I__774 (
            .O(N__4032),
            .I(N__4026));
    Odrv12 I__773 (
            .O(N__4029),
            .I(D_LM_040_in_7));
    Odrv12 I__772 (
            .O(N__4026),
            .I(D_LM_040_in_7));
    InMux I__771 (
            .O(N__4021),
            .I(N__4018));
    LocalMux I__770 (
            .O(N__4018),
            .I(N__4015));
    Span4Mux_v I__769 (
            .O(N__4015),
            .I(N__4012));
    Sp12to4 I__768 (
            .O(N__4012),
            .I(N__4009));
    Span12Mux_h I__767 (
            .O(N__4009),
            .I(N__4006));
    Odrv12 I__766 (
            .O(N__4006),
            .I(D_UU_040_in_7));
    IoInMux I__765 (
            .O(N__4003),
            .I(N__4000));
    LocalMux I__764 (
            .O(N__4000),
            .I(N__3997));
    Span12Mux_s9_v I__763 (
            .O(N__3997),
            .I(N__3994));
    Span12Mux_h I__762 (
            .O(N__3994),
            .I(N__3991));
    Odrv12 I__761 (
            .O(N__3991),
            .I(un1_D_UU_040_7));
    InMux I__760 (
            .O(N__3988),
            .I(N__3985));
    LocalMux I__759 (
            .O(N__3985),
            .I(N__3982));
    Span4Mux_v I__758 (
            .O(N__3982),
            .I(N__3979));
    Sp12to4 I__757 (
            .O(N__3979),
            .I(N__3976));
    Span12Mux_h I__756 (
            .O(N__3976),
            .I(N__3973));
    Odrv12 I__755 (
            .O(N__3973),
            .I(D_LL_AMIGA_in_3));
    IoInMux I__754 (
            .O(N__3970),
            .I(N__3967));
    LocalMux I__753 (
            .O(N__3967),
            .I(N__3964));
    IoSpan4Mux I__752 (
            .O(N__3964),
            .I(N__3961));
    Sp12to4 I__751 (
            .O(N__3961),
            .I(N__3958));
    Span12Mux_s7_v I__750 (
            .O(N__3958),
            .I(N__3955));
    Odrv12 I__749 (
            .O(N__3955),
            .I(un1_D_LL_AMIGA_3));
    InMux I__748 (
            .O(N__3952),
            .I(N__3949));
    LocalMux I__747 (
            .O(N__3949),
            .I(N__3946));
    Span4Mux_v I__746 (
            .O(N__3946),
            .I(N__3943));
    Sp12to4 I__745 (
            .O(N__3943),
            .I(N__3940));
    Span12Mux_h I__744 (
            .O(N__3940),
            .I(N__3937));
    Odrv12 I__743 (
            .O(N__3937),
            .I(D_LL_AMIGA_in_1));
    IoInMux I__742 (
            .O(N__3934),
            .I(N__3931));
    LocalMux I__741 (
            .O(N__3931),
            .I(N__3928));
    Span12Mux_s3_h I__740 (
            .O(N__3928),
            .I(N__3925));
    Span12Mux_h I__739 (
            .O(N__3925),
            .I(N__3922));
    Odrv12 I__738 (
            .O(N__3922),
            .I(un1_D_LL_AMIGA_1));
    InMux I__737 (
            .O(N__3919),
            .I(N__3916));
    LocalMux I__736 (
            .O(N__3916),
            .I(N__3912));
    IoInMux I__735 (
            .O(N__3915),
            .I(N__3909));
    Span12Mux_h I__734 (
            .O(N__3912),
            .I(N__3906));
    LocalMux I__733 (
            .O(N__3909),
            .I(N__3903));
    Odrv12 I__732 (
            .O(N__3906),
            .I(A_AMIGA_c_1));
    Odrv12 I__731 (
            .O(N__3903),
            .I(A_AMIGA_c_1));
    IoInMux I__730 (
            .O(N__3898),
            .I(N__3894));
    InMux I__729 (
            .O(N__3897),
            .I(N__3891));
    LocalMux I__728 (
            .O(N__3894),
            .I(N__3888));
    LocalMux I__727 (
            .O(N__3891),
            .I(N__3885));
    Span4Mux_s3_h I__726 (
            .O(N__3888),
            .I(N__3882));
    Sp12to4 I__725 (
            .O(N__3885),
            .I(N__3879));
    Sp12to4 I__724 (
            .O(N__3882),
            .I(N__3876));
    Span12Mux_v I__723 (
            .O(N__3879),
            .I(N__3873));
    Span12Mux_v I__722 (
            .O(N__3876),
            .I(N__3870));
    Span12Mux_v I__721 (
            .O(N__3873),
            .I(N__3865));
    Span12Mux_h I__720 (
            .O(N__3870),
            .I(N__3865));
    Span12Mux_h I__719 (
            .O(N__3865),
            .I(N__3862));
    Odrv12 I__718 (
            .O(N__3862),
            .I(D_LL_040_in_1));
    InMux I__717 (
            .O(N__3859),
            .I(N__3856));
    LocalMux I__716 (
            .O(N__3856),
            .I(N__3853));
    Span4Mux_h I__715 (
            .O(N__3853),
            .I(N__3850));
    Span4Mux_h I__714 (
            .O(N__3850),
            .I(N__3847));
    Sp12to4 I__713 (
            .O(N__3847),
            .I(N__3844));
    Span12Mux_v I__712 (
            .O(N__3844),
            .I(N__3841));
    Odrv12 I__711 (
            .O(N__3841),
            .I(D_UM_040_in_1));
    IoInMux I__710 (
            .O(N__3838),
            .I(N__3835));
    LocalMux I__709 (
            .O(N__3835),
            .I(N__3832));
    IoSpan4Mux I__708 (
            .O(N__3832),
            .I(N__3829));
    Sp12to4 I__707 (
            .O(N__3829),
            .I(N__3826));
    Span12Mux_s6_h I__706 (
            .O(N__3826),
            .I(N__3823));
    Odrv12 I__705 (
            .O(N__3823),
            .I(un1_D_UM_040_1));
    IoInMux I__704 (
            .O(N__3820),
            .I(N__3817));
    LocalMux I__703 (
            .O(N__3817),
            .I(N__3814));
    IoSpan4Mux I__702 (
            .O(N__3814),
            .I(N__3811));
    IoSpan4Mux I__701 (
            .O(N__3811),
            .I(N__3808));
    Span4Mux_s2_v I__700 (
            .O(N__3808),
            .I(N__3805));
    Span4Mux_v I__699 (
            .O(N__3805),
            .I(N__3802));
    Odrv4 I__698 (
            .O(N__3802),
            .I(LBENn_c_i));
    IoInMux I__697 (
            .O(N__3799),
            .I(N__3796));
    LocalMux I__696 (
            .O(N__3796),
            .I(N__3793));
    Span4Mux_s3_h I__695 (
            .O(N__3793),
            .I(N__3789));
    InMux I__694 (
            .O(N__3792),
            .I(N__3786));
    Sp12to4 I__693 (
            .O(N__3789),
            .I(N__3783));
    LocalMux I__692 (
            .O(N__3786),
            .I(N__3780));
    Span12Mux_v I__691 (
            .O(N__3783),
            .I(N__3777));
    Sp12to4 I__690 (
            .O(N__3780),
            .I(N__3774));
    Span12Mux_h I__689 (
            .O(N__3777),
            .I(N__3769));
    Span12Mux_v I__688 (
            .O(N__3774),
            .I(N__3769));
    Span12Mux_h I__687 (
            .O(N__3769),
            .I(N__3766));
    Span12Mux_v I__686 (
            .O(N__3766),
            .I(N__3763));
    Odrv12 I__685 (
            .O(N__3763),
            .I(D_LM_040_in_1));
    InMux I__684 (
            .O(N__3760),
            .I(N__3757));
    LocalMux I__683 (
            .O(N__3757),
            .I(N__3754));
    Sp12to4 I__682 (
            .O(N__3754),
            .I(N__3751));
    Span12Mux_v I__681 (
            .O(N__3751),
            .I(N__3748));
    Span12Mux_h I__680 (
            .O(N__3748),
            .I(N__3745));
    Odrv12 I__679 (
            .O(N__3745),
            .I(D_UU_040_in_1));
    IoInMux I__678 (
            .O(N__3742),
            .I(N__3739));
    LocalMux I__677 (
            .O(N__3739),
            .I(N__3736));
    Span12Mux_s2_h I__676 (
            .O(N__3736),
            .I(N__3733));
    Span12Mux_h I__675 (
            .O(N__3733),
            .I(N__3730));
    Odrv12 I__674 (
            .O(N__3730),
            .I(un1_D_UU_040_1));
    IoInMux I__673 (
            .O(N__3727),
            .I(N__3724));
    LocalMux I__672 (
            .O(N__3724),
            .I(N__3721));
    Span4Mux_s1_h I__671 (
            .O(N__3721),
            .I(N__3718));
    Sp12to4 I__670 (
            .O(N__3718),
            .I(N__3714));
    InMux I__669 (
            .O(N__3717),
            .I(N__3711));
    Span12Mux_v I__668 (
            .O(N__3714),
            .I(N__3708));
    LocalMux I__667 (
            .O(N__3711),
            .I(N__3705));
    Span12Mux_h I__666 (
            .O(N__3708),
            .I(N__3702));
    Span12Mux_h I__665 (
            .O(N__3705),
            .I(N__3699));
    Span12Mux_h I__664 (
            .O(N__3702),
            .I(N__3694));
    Span12Mux_v I__663 (
            .O(N__3699),
            .I(N__3694));
    Odrv12 I__662 (
            .O(N__3694),
            .I(D_LM_040_in_4));
    InMux I__661 (
            .O(N__3691),
            .I(N__3688));
    LocalMux I__660 (
            .O(N__3688),
            .I(N__3685));
    Span4Mux_v I__659 (
            .O(N__3685),
            .I(N__3682));
    Sp12to4 I__658 (
            .O(N__3682),
            .I(N__3679));
    Span12Mux_h I__657 (
            .O(N__3679),
            .I(N__3676));
    Odrv12 I__656 (
            .O(N__3676),
            .I(D_UU_040_in_4));
    IoInMux I__655 (
            .O(N__3673),
            .I(N__3670));
    LocalMux I__654 (
            .O(N__3670),
            .I(N__3667));
    IoSpan4Mux I__653 (
            .O(N__3667),
            .I(N__3664));
    IoSpan4Mux I__652 (
            .O(N__3664),
            .I(N__3661));
    Span4Mux_s3_v I__651 (
            .O(N__3661),
            .I(N__3658));
    Odrv4 I__650 (
            .O(N__3658),
            .I(un1_D_UU_040_4));
    InMux I__649 (
            .O(N__3655),
            .I(N__3652));
    LocalMux I__648 (
            .O(N__3652),
            .I(N__3649));
    Span12Mux_v I__647 (
            .O(N__3649),
            .I(N__3646));
    Span12Mux_h I__646 (
            .O(N__3646),
            .I(N__3643));
    Odrv12 I__645 (
            .O(N__3643),
            .I(D_UU_040_in_2));
    InMux I__644 (
            .O(N__3640),
            .I(N__3637));
    LocalMux I__643 (
            .O(N__3637),
            .I(N__3633));
    IoInMux I__642 (
            .O(N__3636),
            .I(N__3630));
    Span4Mux_h I__641 (
            .O(N__3633),
            .I(N__3627));
    LocalMux I__640 (
            .O(N__3630),
            .I(N__3624));
    Span4Mux_h I__639 (
            .O(N__3627),
            .I(N__3621));
    Span12Mux_s9_h I__638 (
            .O(N__3624),
            .I(N__3618));
    Sp12to4 I__637 (
            .O(N__3621),
            .I(N__3615));
    Span12Mux_h I__636 (
            .O(N__3618),
            .I(N__3610));
    Span12Mux_v I__635 (
            .O(N__3615),
            .I(N__3610));
    Span12Mux_v I__634 (
            .O(N__3610),
            .I(N__3607));
    Odrv12 I__633 (
            .O(N__3607),
            .I(D_LM_040_in_2));
    IoInMux I__632 (
            .O(N__3604),
            .I(N__3601));
    LocalMux I__631 (
            .O(N__3601),
            .I(N__3598));
    Span4Mux_s2_v I__630 (
            .O(N__3598),
            .I(N__3595));
    Span4Mux_v I__629 (
            .O(N__3595),
            .I(N__3592));
    Sp12to4 I__628 (
            .O(N__3592),
            .I(N__3589));
    Odrv12 I__627 (
            .O(N__3589),
            .I(un1_D_UU_040_2));
    InMux I__626 (
            .O(N__3586),
            .I(N__3583));
    LocalMux I__625 (
            .O(N__3583),
            .I(N__3580));
    Span4Mux_v I__624 (
            .O(N__3580),
            .I(N__3577));
    Sp12to4 I__623 (
            .O(N__3577),
            .I(N__3574));
    Span12Mux_h I__622 (
            .O(N__3574),
            .I(N__3571));
    Odrv12 I__621 (
            .O(N__3571),
            .I(D_LL_AMIGA_in_2));
    IoInMux I__620 (
            .O(N__3568),
            .I(N__3565));
    LocalMux I__619 (
            .O(N__3565),
            .I(N__3562));
    Span12Mux_s4_h I__618 (
            .O(N__3562),
            .I(N__3559));
    Span12Mux_h I__617 (
            .O(N__3559),
            .I(N__3556));
    Odrv12 I__616 (
            .O(N__3556),
            .I(un1_D_LL_AMIGA_2));
    InMux I__615 (
            .O(N__3553),
            .I(N__3550));
    LocalMux I__614 (
            .O(N__3550),
            .I(N__3547));
    Span12Mux_v I__613 (
            .O(N__3547),
            .I(N__3544));
    Span12Mux_h I__612 (
            .O(N__3544),
            .I(N__3541));
    Odrv12 I__611 (
            .O(N__3541),
            .I(D_LL_AMIGA_in_4));
    IoInMux I__610 (
            .O(N__3538),
            .I(N__3535));
    LocalMux I__609 (
            .O(N__3535),
            .I(N__3532));
    IoSpan4Mux I__608 (
            .O(N__3532),
            .I(N__3529));
    Span4Mux_s2_h I__607 (
            .O(N__3529),
            .I(N__3526));
    Sp12to4 I__606 (
            .O(N__3526),
            .I(N__3523));
    Span12Mux_h I__605 (
            .O(N__3523),
            .I(N__3520));
    Odrv12 I__604 (
            .O(N__3520),
            .I(un1_D_LL_AMIGA_4));
    InMux I__603 (
            .O(N__3517),
            .I(N__3514));
    LocalMux I__602 (
            .O(N__3514),
            .I(N__3511));
    Span12Mux_v I__601 (
            .O(N__3511),
            .I(N__3508));
    Span12Mux_h I__600 (
            .O(N__3508),
            .I(N__3505));
    Odrv12 I__599 (
            .O(N__3505),
            .I(D_LL_AMIGA_in_6));
    IoInMux I__598 (
            .O(N__3502),
            .I(N__3499));
    LocalMux I__597 (
            .O(N__3499),
            .I(N__3496));
    Span4Mux_s0_h I__596 (
            .O(N__3496),
            .I(N__3493));
    Span4Mux_h I__595 (
            .O(N__3493),
            .I(N__3490));
    Sp12to4 I__594 (
            .O(N__3490),
            .I(N__3487));
    Span12Mux_s9_v I__593 (
            .O(N__3487),
            .I(N__3484));
    Span12Mux_h I__592 (
            .O(N__3484),
            .I(N__3481));
    Odrv12 I__591 (
            .O(N__3481),
            .I(un1_D_LL_AMIGA_6));
    InMux I__590 (
            .O(N__3478),
            .I(N__3475));
    LocalMux I__589 (
            .O(N__3475),
            .I(N__3472));
    Span4Mux_v I__588 (
            .O(N__3472),
            .I(N__3469));
    Sp12to4 I__587 (
            .O(N__3469),
            .I(N__3466));
    Span12Mux_h I__586 (
            .O(N__3466),
            .I(N__3463));
    Odrv12 I__585 (
            .O(N__3463),
            .I(D_LM_AMIGA_in_0));
    InMux I__584 (
            .O(N__3460),
            .I(N__3457));
    LocalMux I__583 (
            .O(N__3457),
            .I(N__3454));
    Span4Mux_h I__582 (
            .O(N__3454),
            .I(N__3451));
    Sp12to4 I__581 (
            .O(N__3451),
            .I(N__3448));
    Odrv12 I__580 (
            .O(N__3448),
            .I(D_LM_AMIGA_in_2));
    IoInMux I__579 (
            .O(N__3445),
            .I(N__3442));
    LocalMux I__578 (
            .O(N__3442),
            .I(N__3439));
    Span12Mux_s6_h I__577 (
            .O(N__3439),
            .I(N__3436));
    Span12Mux_v I__576 (
            .O(N__3436),
            .I(N__3433));
    Odrv12 I__575 (
            .O(N__3433),
            .I(un1_D_LM_AMIGA_2));
    IoInMux I__574 (
            .O(N__3430),
            .I(N__3427));
    LocalMux I__573 (
            .O(N__3427),
            .I(N__3423));
    InMux I__572 (
            .O(N__3426),
            .I(N__3420));
    IoSpan4Mux I__571 (
            .O(N__3423),
            .I(N__3417));
    LocalMux I__570 (
            .O(N__3420),
            .I(N__3414));
    Span4Mux_s3_h I__569 (
            .O(N__3417),
            .I(N__3411));
    Span4Mux_h I__568 (
            .O(N__3414),
            .I(N__3408));
    Sp12to4 I__567 (
            .O(N__3411),
            .I(N__3405));
    Sp12to4 I__566 (
            .O(N__3408),
            .I(N__3402));
    Span12Mux_v I__565 (
            .O(N__3405),
            .I(N__3399));
    Span12Mux_v I__564 (
            .O(N__3402),
            .I(N__3396));
    Span12Mux_h I__563 (
            .O(N__3399),
            .I(N__3391));
    Span12Mux_v I__562 (
            .O(N__3396),
            .I(N__3391));
    Span12Mux_h I__561 (
            .O(N__3391),
            .I(N__3388));
    Odrv12 I__560 (
            .O(N__3388),
            .I(D_LL_040_in_7));
    InMux I__559 (
            .O(N__3385),
            .I(N__3382));
    LocalMux I__558 (
            .O(N__3382),
            .I(N__3379));
    Span4Mux_v I__557 (
            .O(N__3379),
            .I(N__3376));
    Span4Mux_v I__556 (
            .O(N__3376),
            .I(N__3373));
    Sp12to4 I__555 (
            .O(N__3373),
            .I(N__3370));
    Span12Mux_h I__554 (
            .O(N__3370),
            .I(N__3367));
    Odrv12 I__553 (
            .O(N__3367),
            .I(D_UM_040_in_7));
    IoInMux I__552 (
            .O(N__3364),
            .I(N__3361));
    LocalMux I__551 (
            .O(N__3361),
            .I(N__3358));
    IoSpan4Mux I__550 (
            .O(N__3358),
            .I(N__3355));
    Span4Mux_s3_h I__549 (
            .O(N__3355),
            .I(N__3352));
    Span4Mux_h I__548 (
            .O(N__3352),
            .I(N__3349));
    Span4Mux_h I__547 (
            .O(N__3349),
            .I(N__3346));
    Odrv4 I__546 (
            .O(N__3346),
            .I(un1_D_UM_040_7));
    InMux I__545 (
            .O(N__3343),
            .I(N__3340));
    LocalMux I__544 (
            .O(N__3340),
            .I(N__3337));
    Span4Mux_v I__543 (
            .O(N__3337),
            .I(N__3334));
    Sp12to4 I__542 (
            .O(N__3334),
            .I(N__3331));
    Span12Mux_h I__541 (
            .O(N__3331),
            .I(N__3328));
    Odrv12 I__540 (
            .O(N__3328),
            .I(D_LL_AMIGA_in_0));
    IoInMux I__539 (
            .O(N__3325),
            .I(N__3322));
    LocalMux I__538 (
            .O(N__3322),
            .I(N__3319));
    IoSpan4Mux I__537 (
            .O(N__3319),
            .I(N__3316));
    IoSpan4Mux I__536 (
            .O(N__3316),
            .I(N__3313));
    Span4Mux_s2_h I__535 (
            .O(N__3313),
            .I(N__3310));
    Sp12to4 I__534 (
            .O(N__3310),
            .I(N__3307));
    Span12Mux_s9_h I__533 (
            .O(N__3307),
            .I(N__3304));
    Odrv12 I__532 (
            .O(N__3304),
            .I(un1_D_LL_AMIGA_0));
    IoInMux I__531 (
            .O(N__3301),
            .I(N__3298));
    LocalMux I__530 (
            .O(N__3298),
            .I(N__3295));
    Odrv12 I__529 (
            .O(N__3295),
            .I(LBENn_c_i_0));
    IoInMux I__528 (
            .O(N__3292),
            .I(N__3289));
    LocalMux I__527 (
            .O(N__3289),
            .I(N__3286));
    Span12Mux_s6_v I__526 (
            .O(N__3286),
            .I(N__3283));
    Odrv12 I__525 (
            .O(N__3283),
            .I(TSn_c));
    InMux I__524 (
            .O(N__3280),
            .I(N__3277));
    LocalMux I__523 (
            .O(N__3277),
            .I(N__3274));
    Span4Mux_v I__522 (
            .O(N__3274),
            .I(N__3271));
    Sp12to4 I__521 (
            .O(N__3271),
            .I(N__3268));
    Span12Mux_h I__520 (
            .O(N__3268),
            .I(N__3265));
    Odrv12 I__519 (
            .O(N__3265),
            .I(D_LL_AMIGA_in_5));
    IoInMux I__518 (
            .O(N__3262),
            .I(N__3259));
    LocalMux I__517 (
            .O(N__3259),
            .I(N__3256));
    Span4Mux_s3_h I__516 (
            .O(N__3256),
            .I(N__3253));
    Sp12to4 I__515 (
            .O(N__3253),
            .I(N__3250));
    Span12Mux_s11_v I__514 (
            .O(N__3250),
            .I(N__3247));
    Span12Mux_h I__513 (
            .O(N__3247),
            .I(N__3244));
    Odrv12 I__512 (
            .O(N__3244),
            .I(un1_D_LL_AMIGA_5));
    InMux I__511 (
            .O(N__3241),
            .I(N__3238));
    LocalMux I__510 (
            .O(N__3238),
            .I(N__3235));
    Span4Mux_v I__509 (
            .O(N__3235),
            .I(N__3232));
    Sp12to4 I__508 (
            .O(N__3232),
            .I(N__3229));
    Span12Mux_h I__507 (
            .O(N__3229),
            .I(N__3226));
    Odrv12 I__506 (
            .O(N__3226),
            .I(D_LM_AMIGA_in_4));
    IoInMux I__505 (
            .O(N__3223),
            .I(N__3220));
    LocalMux I__504 (
            .O(N__3220),
            .I(N__3217));
    IoSpan4Mux I__503 (
            .O(N__3217),
            .I(N__3214));
    IoSpan4Mux I__502 (
            .O(N__3214),
            .I(N__3211));
    Span4Mux_s2_h I__501 (
            .O(N__3211),
            .I(N__3208));
    Sp12to4 I__500 (
            .O(N__3208),
            .I(N__3205));
    Span12Mux_s11_h I__499 (
            .O(N__3205),
            .I(N__3202));
    Odrv12 I__498 (
            .O(N__3202),
            .I(un1_D_LM_AMIGA_4));
    InMux I__497 (
            .O(N__3199),
            .I(N__3196));
    LocalMux I__496 (
            .O(N__3196),
            .I(N__3193));
    Span12Mux_h I__495 (
            .O(N__3193),
            .I(N__3190));
    Odrv12 I__494 (
            .O(N__3190),
            .I(D_UM_040_in_6));
    IoInMux I__493 (
            .O(N__3187),
            .I(N__3184));
    LocalMux I__492 (
            .O(N__3184),
            .I(N__3181));
    IoSpan4Mux I__491 (
            .O(N__3181),
            .I(N__3177));
    InMux I__490 (
            .O(N__3180),
            .I(N__3174));
    IoSpan4Mux I__489 (
            .O(N__3177),
            .I(N__3171));
    LocalMux I__488 (
            .O(N__3174),
            .I(N__3168));
    Span4Mux_s2_h I__487 (
            .O(N__3171),
            .I(N__3165));
    Span4Mux_v I__486 (
            .O(N__3168),
            .I(N__3162));
    Sp12to4 I__485 (
            .O(N__3165),
            .I(N__3159));
    Sp12to4 I__484 (
            .O(N__3162),
            .I(N__3156));
    Span12Mux_h I__483 (
            .O(N__3159),
            .I(N__3153));
    Span12Mux_h I__482 (
            .O(N__3156),
            .I(N__3150));
    Span12Mux_h I__481 (
            .O(N__3153),
            .I(N__3145));
    Span12Mux_v I__480 (
            .O(N__3150),
            .I(N__3145));
    Odrv12 I__479 (
            .O(N__3145),
            .I(D_LL_040_in_6));
    IoInMux I__478 (
            .O(N__3142),
            .I(N__3139));
    LocalMux I__477 (
            .O(N__3139),
            .I(N__3136));
    IoSpan4Mux I__476 (
            .O(N__3136),
            .I(N__3133));
    Sp12to4 I__475 (
            .O(N__3133),
            .I(N__3130));
    Span12Mux_s6_h I__474 (
            .O(N__3130),
            .I(N__3127));
    Span12Mux_v I__473 (
            .O(N__3127),
            .I(N__3124));
    Odrv12 I__472 (
            .O(N__3124),
            .I(un1_D_UM_040_6));
    IoInMux I__471 (
            .O(N__3121),
            .I(N__3118));
    LocalMux I__470 (
            .O(N__3118),
            .I(N__3114));
    InMux I__469 (
            .O(N__3117),
            .I(N__3111));
    IoSpan4Mux I__468 (
            .O(N__3114),
            .I(N__3108));
    LocalMux I__467 (
            .O(N__3111),
            .I(N__3105));
    Span4Mux_s2_h I__466 (
            .O(N__3108),
            .I(N__3102));
    Span4Mux_v I__465 (
            .O(N__3105),
            .I(N__3099));
    Sp12to4 I__464 (
            .O(N__3102),
            .I(N__3096));
    Sp12to4 I__463 (
            .O(N__3099),
            .I(N__3093));
    Span12Mux_h I__462 (
            .O(N__3096),
            .I(N__3088));
    Span12Mux_v I__461 (
            .O(N__3093),
            .I(N__3088));
    Span12Mux_h I__460 (
            .O(N__3088),
            .I(N__3085));
    Odrv12 I__459 (
            .O(N__3085),
            .I(D_LL_040_in_2));
    InMux I__458 (
            .O(N__3082),
            .I(N__3079));
    LocalMux I__457 (
            .O(N__3079),
            .I(N__3076));
    Span12Mux_h I__456 (
            .O(N__3076),
            .I(N__3073));
    Odrv12 I__455 (
            .O(N__3073),
            .I(D_UM_040_in_2));
    IoInMux I__454 (
            .O(N__3070),
            .I(N__3067));
    LocalMux I__453 (
            .O(N__3067),
            .I(N__3064));
    Span4Mux_s3_h I__452 (
            .O(N__3064),
            .I(N__3061));
    Span4Mux_v I__451 (
            .O(N__3061),
            .I(N__3058));
    Sp12to4 I__450 (
            .O(N__3058),
            .I(N__3055));
    Odrv12 I__449 (
            .O(N__3055),
            .I(un1_D_UM_040_2));
    InMux I__448 (
            .O(N__3052),
            .I(N__3049));
    LocalMux I__447 (
            .O(N__3049),
            .I(N__3046));
    Span4Mux_v I__446 (
            .O(N__3046),
            .I(N__3043));
    Sp12to4 I__445 (
            .O(N__3043),
            .I(N__3040));
    Odrv12 I__444 (
            .O(N__3040),
            .I(D_LM_AMIGA_in_5));
    IoInMux I__443 (
            .O(N__3037),
            .I(N__3034));
    LocalMux I__442 (
            .O(N__3034),
            .I(N__3031));
    IoSpan4Mux I__441 (
            .O(N__3031),
            .I(N__3028));
    Span4Mux_s2_h I__440 (
            .O(N__3028),
            .I(N__3025));
    Span4Mux_v I__439 (
            .O(N__3025),
            .I(N__3022));
    Sp12to4 I__438 (
            .O(N__3022),
            .I(N__3019));
    Span12Mux_s11_h I__437 (
            .O(N__3019),
            .I(N__3016));
    Odrv12 I__436 (
            .O(N__3016),
            .I(un1_D_LM_AMIGA_5));
    InMux I__435 (
            .O(N__3013),
            .I(N__3010));
    LocalMux I__434 (
            .O(N__3010),
            .I(N__3007));
    Span4Mux_h I__433 (
            .O(N__3007),
            .I(N__3004));
    Span4Mux_v I__432 (
            .O(N__3004),
            .I(N__3001));
    Sp12to4 I__431 (
            .O(N__3001),
            .I(N__2998));
    Odrv12 I__430 (
            .O(N__2998),
            .I(D_LM_AMIGA_in_6));
    IoInMux I__429 (
            .O(N__2995),
            .I(N__2992));
    LocalMux I__428 (
            .O(N__2992),
            .I(N__2989));
    Span12Mux_s2_h I__427 (
            .O(N__2989),
            .I(N__2986));
    Span12Mux_h I__426 (
            .O(N__2986),
            .I(N__2983));
    Odrv12 I__425 (
            .O(N__2983),
            .I(un1_D_LM_AMIGA_6));
    InMux I__424 (
            .O(N__2980),
            .I(N__2976));
    IoInMux I__423 (
            .O(N__2979),
            .I(N__2973));
    LocalMux I__422 (
            .O(N__2976),
            .I(N__2970));
    LocalMux I__421 (
            .O(N__2973),
            .I(N__2967));
    Span4Mux_v I__420 (
            .O(N__2970),
            .I(N__2964));
    Span4Mux_s2_h I__419 (
            .O(N__2967),
            .I(N__2961));
    Sp12to4 I__418 (
            .O(N__2964),
            .I(N__2958));
    Span4Mux_v I__417 (
            .O(N__2961),
            .I(N__2955));
    Span12Mux_h I__416 (
            .O(N__2958),
            .I(N__2952));
    Sp12to4 I__415 (
            .O(N__2955),
            .I(N__2949));
    Span12Mux_v I__414 (
            .O(N__2952),
            .I(N__2946));
    Span12Mux_s11_h I__413 (
            .O(N__2949),
            .I(N__2943));
    Span12Mux_v I__412 (
            .O(N__2946),
            .I(N__2938));
    Span12Mux_h I__411 (
            .O(N__2943),
            .I(N__2938));
    Odrv12 I__410 (
            .O(N__2938),
            .I(D_LL_040_in_3));
    InMux I__409 (
            .O(N__2935),
            .I(N__2932));
    LocalMux I__408 (
            .O(N__2932),
            .I(N__2929));
    Sp12to4 I__407 (
            .O(N__2929),
            .I(N__2926));
    Span12Mux_v I__406 (
            .O(N__2926),
            .I(N__2923));
    Span12Mux_h I__405 (
            .O(N__2923),
            .I(N__2920));
    Odrv12 I__404 (
            .O(N__2920),
            .I(D_UM_040_in_3));
    IoInMux I__403 (
            .O(N__2917),
            .I(N__2914));
    LocalMux I__402 (
            .O(N__2914),
            .I(N__2911));
    IoSpan4Mux I__401 (
            .O(N__2911),
            .I(N__2908));
    Span4Mux_s3_h I__400 (
            .O(N__2908),
            .I(N__2905));
    Span4Mux_h I__399 (
            .O(N__2905),
            .I(N__2902));
    Span4Mux_h I__398 (
            .O(N__2902),
            .I(N__2899));
    Odrv4 I__397 (
            .O(N__2899),
            .I(un1_D_UM_040_3));
    IoInMux I__396 (
            .O(N__2896),
            .I(N__2893));
    LocalMux I__395 (
            .O(N__2893),
            .I(N__2888));
    IoInMux I__394 (
            .O(N__2892),
            .I(N__2883));
    IoInMux I__393 (
            .O(N__2891),
            .I(N__2883));
    Span4Mux_s0_v I__392 (
            .O(N__2888),
            .I(N__2879));
    LocalMux I__391 (
            .O(N__2883),
            .I(N__2876));
    IoInMux I__390 (
            .O(N__2882),
            .I(N__2873));
    Span4Mux_h I__389 (
            .O(N__2879),
            .I(N__2870));
    Span4Mux_s0_v I__388 (
            .O(N__2876),
            .I(N__2867));
    LocalMux I__387 (
            .O(N__2873),
            .I(N__2864));
    Span4Mux_h I__386 (
            .O(N__2870),
            .I(N__2859));
    Span4Mux_h I__385 (
            .O(N__2867),
            .I(N__2859));
    Span12Mux_s7_h I__384 (
            .O(N__2864),
            .I(N__2856));
    Span4Mux_v I__383 (
            .O(N__2859),
            .I(N__2853));
    Span12Mux_h I__382 (
            .O(N__2856),
            .I(N__2850));
    Span4Mux_v I__381 (
            .O(N__2853),
            .I(N__2847));
    Odrv12 I__380 (
            .O(N__2850),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__379 (
            .O(N__2847),
            .I(CONSTANT_ONE_NET));
    InMux I__378 (
            .O(N__2842),
            .I(N__2839));
    LocalMux I__377 (
            .O(N__2839),
            .I(N__2836));
    Span4Mux_v I__376 (
            .O(N__2836),
            .I(N__2833));
    Span4Mux_h I__375 (
            .O(N__2833),
            .I(N__2830));
    Sp12to4 I__374 (
            .O(N__2830),
            .I(N__2827));
    Span12Mux_h I__373 (
            .O(N__2827),
            .I(N__2824));
    Odrv12 I__372 (
            .O(N__2824),
            .I(D_UU_040_in_6));
    IoInMux I__371 (
            .O(N__2821),
            .I(N__2818));
    LocalMux I__370 (
            .O(N__2818),
            .I(N__2815));
    Span4Mux_s2_h I__369 (
            .O(N__2815),
            .I(N__2811));
    InMux I__368 (
            .O(N__2814),
            .I(N__2808));
    Span4Mux_v I__367 (
            .O(N__2811),
            .I(N__2805));
    LocalMux I__366 (
            .O(N__2808),
            .I(N__2802));
    Sp12to4 I__365 (
            .O(N__2805),
            .I(N__2799));
    Sp12to4 I__364 (
            .O(N__2802),
            .I(N__2796));
    Span12Mux_h I__363 (
            .O(N__2799),
            .I(N__2791));
    Span12Mux_s11_v I__362 (
            .O(N__2796),
            .I(N__2791));
    Span12Mux_h I__361 (
            .O(N__2791),
            .I(N__2788));
    Odrv12 I__360 (
            .O(N__2788),
            .I(D_LM_040_in_6));
    IoInMux I__359 (
            .O(N__2785),
            .I(N__2782));
    LocalMux I__358 (
            .O(N__2782),
            .I(N__2779));
    IoSpan4Mux I__357 (
            .O(N__2779),
            .I(N__2776));
    Sp12to4 I__356 (
            .O(N__2776),
            .I(N__2773));
    Span12Mux_s6_v I__355 (
            .O(N__2773),
            .I(N__2770));
    Odrv12 I__354 (
            .O(N__2770),
            .I(un1_D_UU_040_6));
    InMux I__353 (
            .O(N__2767),
            .I(N__2764));
    LocalMux I__352 (
            .O(N__2764),
            .I(N__2761));
    Span4Mux_v I__351 (
            .O(N__2761),
            .I(N__2758));
    Span4Mux_h I__350 (
            .O(N__2758),
            .I(N__2755));
    Sp12to4 I__349 (
            .O(N__2755),
            .I(N__2752));
    Span12Mux_h I__348 (
            .O(N__2752),
            .I(N__2749));
    Odrv12 I__347 (
            .O(N__2749),
            .I(D_UU_040_in_0));
    IoInMux I__346 (
            .O(N__2746),
            .I(N__2742));
    InMux I__345 (
            .O(N__2745),
            .I(N__2739));
    LocalMux I__344 (
            .O(N__2742),
            .I(N__2736));
    LocalMux I__343 (
            .O(N__2739),
            .I(N__2733));
    IoSpan4Mux I__342 (
            .O(N__2736),
            .I(N__2730));
    Span4Mux_v I__341 (
            .O(N__2733),
            .I(N__2727));
    IoSpan4Mux I__340 (
            .O(N__2730),
            .I(N__2724));
    Sp12to4 I__339 (
            .O(N__2727),
            .I(N__2721));
    Span4Mux_s2_h I__338 (
            .O(N__2724),
            .I(N__2718));
    Span12Mux_h I__337 (
            .O(N__2721),
            .I(N__2715));
    Sp12to4 I__336 (
            .O(N__2718),
            .I(N__2712));
    Span12Mux_v I__335 (
            .O(N__2715),
            .I(N__2709));
    Span12Mux_h I__334 (
            .O(N__2712),
            .I(N__2706));
    Span12Mux_v I__333 (
            .O(N__2709),
            .I(N__2701));
    Span12Mux_h I__332 (
            .O(N__2706),
            .I(N__2701));
    Odrv12 I__331 (
            .O(N__2701),
            .I(D_LM_040_in_0));
    IoInMux I__330 (
            .O(N__2698),
            .I(N__2695));
    LocalMux I__329 (
            .O(N__2695),
            .I(N__2692));
    IoSpan4Mux I__328 (
            .O(N__2692),
            .I(N__2689));
    IoSpan4Mux I__327 (
            .O(N__2689),
            .I(N__2686));
    Span4Mux_s3_v I__326 (
            .O(N__2686),
            .I(N__2683));
    Odrv4 I__325 (
            .O(N__2683),
            .I(un1_D_UU_040_0));
    InMux I__324 (
            .O(N__2680),
            .I(N__2677));
    LocalMux I__323 (
            .O(N__2677),
            .I(N__2674));
    Span12Mux_v I__322 (
            .O(N__2674),
            .I(N__2671));
    Span12Mux_h I__321 (
            .O(N__2671),
            .I(N__2668));
    Odrv12 I__320 (
            .O(N__2668),
            .I(D_LM_AMIGA_in_3));
    IoInMux I__319 (
            .O(N__2665),
            .I(N__2662));
    LocalMux I__318 (
            .O(N__2662),
            .I(N__2659));
    Span4Mux_s0_h I__317 (
            .O(N__2659),
            .I(N__2656));
    Sp12to4 I__316 (
            .O(N__2656),
            .I(N__2653));
    Span12Mux_v I__315 (
            .O(N__2653),
            .I(N__2650));
    Span12Mux_h I__314 (
            .O(N__2650),
            .I(N__2647));
    Odrv12 I__313 (
            .O(N__2647),
            .I(un1_D_LM_AMIGA_3));
    IoInMux I__312 (
            .O(N__2644),
            .I(N__2641));
    LocalMux I__311 (
            .O(N__2641),
            .I(N__2638));
    Span4Mux_s0_v I__310 (
            .O(N__2638),
            .I(N__2635));
    Sp12to4 I__309 (
            .O(N__2635),
            .I(N__2632));
    Span12Mux_h I__308 (
            .O(N__2632),
            .I(N__2629));
    Span12Mux_v I__307 (
            .O(N__2629),
            .I(N__2626));
    Span12Mux_v I__306 (
            .O(N__2626),
            .I(N__2623));
    Odrv12 I__305 (
            .O(N__2623),
            .I(TAn_in));
    InMux I__304 (
            .O(N__2620),
            .I(N__2617));
    LocalMux I__303 (
            .O(N__2617),
            .I(N__2614));
    Span12Mux_h I__302 (
            .O(N__2614),
            .I(N__2611));
    Odrv12 I__301 (
            .O(N__2611),
            .I(A_040_c_1));
    InMux I__300 (
            .O(N__2608),
            .I(N__2605));
    LocalMux I__299 (
            .O(N__2605),
            .I(N__2602));
    Span4Mux_h I__298 (
            .O(N__2602),
            .I(N__2599));
    Span4Mux_v I__297 (
            .O(N__2599),
            .I(N__2596));
    Odrv4 I__296 (
            .O(N__2596),
            .I(A_040_c_0));
    IoInMux I__295 (
            .O(N__2593),
            .I(N__2590));
    LocalMux I__294 (
            .O(N__2590),
            .I(N__2587));
    Span4Mux_s2_v I__293 (
            .O(N__2587),
            .I(N__2584));
    Span4Mux_v I__292 (
            .O(N__2584),
            .I(N__2581));
    Odrv4 I__291 (
            .O(N__2581),
            .I(A_AMIGA_c_0));
    IoInMux I__290 (
            .O(N__2578),
            .I(N__2575));
    LocalMux I__289 (
            .O(N__2575),
            .I(N__2569));
    IoInMux I__288 (
            .O(N__2574),
            .I(N__2566));
    IoInMux I__287 (
            .O(N__2573),
            .I(N__2563));
    IoInMux I__286 (
            .O(N__2572),
            .I(N__2560));
    IoSpan4Mux I__285 (
            .O(N__2569),
            .I(N__2549));
    LocalMux I__284 (
            .O(N__2566),
            .I(N__2549));
    LocalMux I__283 (
            .O(N__2563),
            .I(N__2549));
    LocalMux I__282 (
            .O(N__2560),
            .I(N__2549));
    IoInMux I__281 (
            .O(N__2559),
            .I(N__2546));
    IoInMux I__280 (
            .O(N__2558),
            .I(N__2543));
    IoSpan4Mux I__279 (
            .O(N__2549),
            .I(N__2535));
    LocalMux I__278 (
            .O(N__2546),
            .I(N__2535));
    LocalMux I__277 (
            .O(N__2543),
            .I(N__2535));
    IoInMux I__276 (
            .O(N__2542),
            .I(N__2532));
    IoSpan4Mux I__275 (
            .O(N__2535),
            .I(N__2526));
    LocalMux I__274 (
            .O(N__2532),
            .I(N__2523));
    IoInMux I__273 (
            .O(N__2531),
            .I(N__2520));
    IoInMux I__272 (
            .O(N__2530),
            .I(N__2517));
    IoInMux I__271 (
            .O(N__2529),
            .I(N__2514));
    IoSpan4Mux I__270 (
            .O(N__2526),
            .I(N__2496));
    IoSpan4Mux I__269 (
            .O(N__2523),
            .I(N__2496));
    LocalMux I__268 (
            .O(N__2520),
            .I(N__2496));
    LocalMux I__267 (
            .O(N__2517),
            .I(N__2496));
    LocalMux I__266 (
            .O(N__2514),
            .I(N__2496));
    IoInMux I__265 (
            .O(N__2513),
            .I(N__2493));
    IoInMux I__264 (
            .O(N__2512),
            .I(N__2490));
    IoInMux I__263 (
            .O(N__2511),
            .I(N__2485));
    IoInMux I__262 (
            .O(N__2510),
            .I(N__2482));
    IoInMux I__261 (
            .O(N__2509),
            .I(N__2479));
    IoInMux I__260 (
            .O(N__2508),
            .I(N__2476));
    IoInMux I__259 (
            .O(N__2507),
            .I(N__2469));
    IoSpan4Mux I__258 (
            .O(N__2496),
            .I(N__2460));
    LocalMux I__257 (
            .O(N__2493),
            .I(N__2460));
    LocalMux I__256 (
            .O(N__2490),
            .I(N__2460));
    IoInMux I__255 (
            .O(N__2489),
            .I(N__2457));
    IoInMux I__254 (
            .O(N__2488),
            .I(N__2454));
    LocalMux I__253 (
            .O(N__2485),
            .I(N__2440));
    LocalMux I__252 (
            .O(N__2482),
            .I(N__2440));
    LocalMux I__251 (
            .O(N__2479),
            .I(N__2440));
    LocalMux I__250 (
            .O(N__2476),
            .I(N__2440));
    IoInMux I__249 (
            .O(N__2475),
            .I(N__2437));
    IoInMux I__248 (
            .O(N__2474),
            .I(N__2434));
    IoInMux I__247 (
            .O(N__2473),
            .I(N__2431));
    IoInMux I__246 (
            .O(N__2472),
            .I(N__2428));
    LocalMux I__245 (
            .O(N__2469),
            .I(N__2425));
    IoInMux I__244 (
            .O(N__2468),
            .I(N__2422));
    IoInMux I__243 (
            .O(N__2467),
            .I(N__2419));
    IoSpan4Mux I__242 (
            .O(N__2460),
            .I(N__2412));
    LocalMux I__241 (
            .O(N__2457),
            .I(N__2412));
    LocalMux I__240 (
            .O(N__2454),
            .I(N__2412));
    IoInMux I__239 (
            .O(N__2453),
            .I(N__2409));
    IoInMux I__238 (
            .O(N__2452),
            .I(N__2406));
    IoInMux I__237 (
            .O(N__2451),
            .I(N__2403));
    IoInMux I__236 (
            .O(N__2450),
            .I(N__2400));
    IoInMux I__235 (
            .O(N__2449),
            .I(N__2397));
    IoSpan4Mux I__234 (
            .O(N__2440),
            .I(N__2386));
    LocalMux I__233 (
            .O(N__2437),
            .I(N__2386));
    LocalMux I__232 (
            .O(N__2434),
            .I(N__2386));
    LocalMux I__231 (
            .O(N__2431),
            .I(N__2386));
    LocalMux I__230 (
            .O(N__2428),
            .I(N__2371));
    IoSpan4Mux I__229 (
            .O(N__2425),
            .I(N__2371));
    LocalMux I__228 (
            .O(N__2422),
            .I(N__2371));
    LocalMux I__227 (
            .O(N__2419),
            .I(N__2371));
    IoSpan4Mux I__226 (
            .O(N__2412),
            .I(N__2371));
    LocalMux I__225 (
            .O(N__2409),
            .I(N__2371));
    LocalMux I__224 (
            .O(N__2406),
            .I(N__2371));
    LocalMux I__223 (
            .O(N__2403),
            .I(N__2366));
    LocalMux I__222 (
            .O(N__2400),
            .I(N__2366));
    LocalMux I__221 (
            .O(N__2397),
            .I(N__2363));
    IoInMux I__220 (
            .O(N__2396),
            .I(N__2360));
    IoInMux I__219 (
            .O(N__2395),
            .I(N__2357));
    IoSpan4Mux I__218 (
            .O(N__2386),
            .I(N__2354));
    IoSpan4Mux I__217 (
            .O(N__2371),
            .I(N__2351));
    Span12Mux_s7_h I__216 (
            .O(N__2366),
            .I(N__2348));
    Span12Mux_s9_h I__215 (
            .O(N__2363),
            .I(N__2345));
    LocalMux I__214 (
            .O(N__2360),
            .I(N__2340));
    LocalMux I__213 (
            .O(N__2357),
            .I(N__2340));
    Span4Mux_s1_v I__212 (
            .O(N__2354),
            .I(N__2337));
    Span4Mux_s3_h I__211 (
            .O(N__2351),
            .I(N__2334));
    Span12Mux_v I__210 (
            .O(N__2348),
            .I(N__2331));
    Span12Mux_v I__209 (
            .O(N__2345),
            .I(N__2326));
    Span12Mux_s9_h I__208 (
            .O(N__2340),
            .I(N__2326));
    Span4Mux_v I__207 (
            .O(N__2337),
            .I(N__2323));
    Span4Mux_h I__206 (
            .O(N__2334),
            .I(N__2320));
    Odrv12 I__205 (
            .O(N__2331),
            .I(RnW_c_i));
    Odrv12 I__204 (
            .O(N__2326),
            .I(RnW_c_i));
    Odrv4 I__203 (
            .O(N__2323),
            .I(RnW_c_i));
    Odrv4 I__202 (
            .O(N__2320),
            .I(RnW_c_i));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net ),
            .I(N__4454));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .I(N__4452));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net ),
            .I(N__4458));
    INV \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C  (
            .O(\INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net ),
            .I(N__4449));
    INV \INVU111_CYCLE_SM.LW_CYCLEC  (
            .O(\INVU111_CYCLE_SM.LW_CYCLEC_net ),
            .I(N__4451));
    INV \INVU111_CYCLE_SM.CYCLE_STATE_1C  (
            .O(\INVU111_CYCLE_SM.CYCLE_STATE_1C_net ),
            .I(N__4453));
    INV \INVU111_CYCLE_SM.TA_ENC  (
            .O(\INVU111_CYCLE_SM.TA_ENC_net ),
            .I(N__4448));
    INV \INVU111_CYCLE_SM.LW_CYCLE_STARTC  (
            .O(\INVU111_CYCLE_SM.LW_CYCLE_STARTC_net ),
            .I(N__4450));
    INV \INVU111_CYCLE_SM.TSnC  (
            .O(\INVU111_CYCLE_SM.TSnC_net ),
            .I(N__5673));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_1  (
            .in0(N__4396),
            .in1(N__2620),
            .in2(_gnd_net_),
            .in3(N__7272),
            .lcout(A_AMIGA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_7  (
            .in0(N__2608),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7273),
            .lcout(A_AMIGA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RnW_c_sbtinv_LC_6_18_6.C_ON=1'b0;
    defparam RnW_c_sbtinv_LC_6_18_6.SEQ_MODE=4'b0000;
    defparam RnW_c_sbtinv_LC_6_18_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 RnW_c_sbtinv_LC_6_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6041),
            .lcout(RnW_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_9_10_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_9_10_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_9_10_7  (
            .in0(N__3117),
            .in1(N__4759),
            .in2(_gnd_net_),
            .in3(N__3082),
            .lcout(un1_D_UM_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_9_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_9_15_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_9_15_0  (
            .in0(N__3052),
            .in1(N__4859),
            .in2(_gnd_net_),
            .in3(N__6825),
            .lcout(un1_D_LM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_9_15_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_9_15_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_9_15_3  (
            .in0(N__4860),
            .in1(N__6554),
            .in2(_gnd_net_),
            .in3(N__3013),
            .lcout(un1_D_LM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_9_18_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_9_18_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_9_18_1  (
            .in0(N__2980),
            .in1(N__4869),
            .in2(_gnd_net_),
            .in3(N__2935),
            .lcout(un1_D_UM_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_9_18_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_9_18_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_9_18_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_9_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_9_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_9_20_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_9_20_3  (
            .in0(N__4879),
            .in1(N__2842),
            .in2(_gnd_net_),
            .in3(N__2814),
            .lcout(un1_D_UU_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_9_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_9_20_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_9_20_4  (
            .in0(N__2767),
            .in1(N__4880),
            .in2(_gnd_net_),
            .in3(N__2745),
            .lcout(un1_D_UU_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_10_12_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_10_12_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_10_12_2  (
            .in0(N__6680),
            .in1(N__4830),
            .in2(_gnd_net_),
            .in3(N__2680),
            .lcout(un1_D_LM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_10_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_10_12_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_10_12_4  (
            .in0(N__4829),
            .in1(N__5548),
            .in2(_gnd_net_),
            .in3(N__3460),
            .lcout(un1_D_LM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_10_19_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_10_19_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_10_19_1  (
            .in0(N__3426),
            .in1(N__4878),
            .in2(_gnd_net_),
            .in3(N__3385),
            .lcout(un1_D_UM_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_11_1_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_11_1_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_11_1_0  (
            .in0(N__3343),
            .in1(N__4855),
            .in2(_gnd_net_),
            .in3(N__6466),
            .lcout(un1_D_LL_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LBENn_c_sbtinv_LC_11_1_1.C_ON=1'b0;
    defparam LBENn_c_sbtinv_LC_11_1_1.SEQ_MODE=4'b0000;
    defparam LBENn_c_sbtinv_LC_11_1_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 LBENn_c_sbtinv_LC_11_1_1 (
            .in0(N__5831),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(LBENn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TSn_LC_11_1_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TSn_LC_11_1_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TSn_LC_11_1_7 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \U111_CYCLE_SM.TSn_LC_11_1_7  (
            .in0(N__6094),
            .in1(_gnd_net_),
            .in2(N__5849),
            .in3(N__5146),
            .lcout(TSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TSnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_6  (
            .in0(N__6772),
            .in1(N__4814),
            .in2(_gnd_net_),
            .in3(N__3280),
            .lcout(un1_D_LL_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_11_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_11_13_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_11_13_2  (
            .in0(N__4818),
            .in1(N__6634),
            .in2(_gnd_net_),
            .in3(N__3241),
            .lcout(un1_D_LM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_11_13_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_11_13_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_11_13_4  (
            .in0(N__4817),
            .in1(N__3199),
            .in2(_gnd_net_),
            .in3(N__3180),
            .lcout(un1_D_UM_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_11_15_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_11_15_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_11_15_4  (
            .in0(N__3897),
            .in1(N__4870),
            .in2(_gnd_net_),
            .in3(N__3859),
            .lcout(un1_D_UM_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BUFENn_obuf_RNO_LC_11_18_1.C_ON=1'b0;
    defparam BUFENn_obuf_RNO_LC_11_18_1.SEQ_MODE=4'b0000;
    defparam BUFENn_obuf_RNO_LC_11_18_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 BUFENn_obuf_RNO_LC_11_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5867),
            .lcout(LBENn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_11_18_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_11_18_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_11_18_3  (
            .in0(N__3792),
            .in1(N__4871),
            .in2(_gnd_net_),
            .in3(N__3760),
            .lcout(un1_D_UU_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_11_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_11_20_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_11_20_2  (
            .in0(N__3717),
            .in1(N__4882),
            .in2(_gnd_net_),
            .in3(N__3691),
            .lcout(un1_D_UU_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_11_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_11_20_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_11_20_7  (
            .in0(N__3655),
            .in1(N__4881),
            .in2(_gnd_net_),
            .in3(N__3640),
            .lcout(un1_D_UU_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_12_3_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_12_3_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_12_3_6  (
            .in0(N__6367),
            .in1(N__4815),
            .in2(_gnd_net_),
            .in3(N__3586),
            .lcout(un1_D_LL_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_12_3_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_12_3_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_12_3_7  (
            .in0(N__4816),
            .in1(N__7324),
            .in2(_gnd_net_),
            .in3(N__3553),
            .lcout(un1_D_LL_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_12_6_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_12_6_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_12_6_2  (
            .in0(N__6415),
            .in1(N__4819),
            .in2(_gnd_net_),
            .in3(N__3517),
            .lcout(un1_D_LL_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_12_7_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_12_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_12_7_0  (
            .in0(N__4760),
            .in1(N__6910),
            .in2(_gnd_net_),
            .in3(N__3478),
            .lcout(un1_D_LM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_12_7_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_12_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_12_7_5  (
            .in0(N__6974),
            .in1(N__4761),
            .in2(_gnd_net_),
            .in3(N__4351),
            .lcout(un1_D_LL_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_12_9_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_12_9_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_12_9_0  (
            .in0(N__4708),
            .in1(N__4311),
            .in2(_gnd_net_),
            .in3(N__4270),
            .lcout(un1_D_UM_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_12_19_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_12_19_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_12_19_3  (
            .in0(N__4856),
            .in1(N__4237),
            .in2(_gnd_net_),
            .in3(N__4216),
            .lcout(un1_D_UM_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_12_20_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_12_20_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_12_20_0  (
            .in0(N__4146),
            .in1(N__4857),
            .in2(_gnd_net_),
            .in3(N__4105),
            .lcout(un1_D_UU_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_12_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_12_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_12_20_1  (
            .in0(N__4858),
            .in1(N__4056),
            .in2(_gnd_net_),
            .in3(N__4021),
            .lcout(un1_D_UU_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_13_2_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_13_2_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_13_2_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_13_2_4  (
            .in0(N__3988),
            .in1(N__4808),
            .in2(_gnd_net_),
            .in3(N__7123),
            .lcout(un1_D_LL_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_13_2_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_13_2_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_13_2_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_13_2_6  (
            .in0(N__5770),
            .in1(N__4807),
            .in2(_gnd_net_),
            .in3(N__3952),
            .lcout(un1_D_LL_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIM3VM1_LC_13_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIM3VM1_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIM3VM1_LC_13_10_3 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIM3VM1_LC_13_10_3  (
            .in0(N__7263),
            .in1(N__5038),
            .in2(_gnd_net_),
            .in3(N__3919),
            .lcout(\U111_CYCLE_SM.FLIP ),
            .ltout(\U111_CYCLE_SM.FLIP_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_13_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_13_10_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_13_10_4  (
            .in0(N__4558),
            .in1(_gnd_net_),
            .in2(N__4546),
            .in3(N__5977),
            .lcout(un1_D_LM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_13_11_0.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_13_11_0.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_13_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_THRU_LUT4_0_LC_13_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5689),
            .lcout(GB_BUFFER_CLK40_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_11_2.C_ON=1'b0;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_11_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_11_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_11_2 (
            .in0(N__4462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_CLK80_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_START_LC_13_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_LC_13_13_0 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_START_LC_13_13_0  (
            .in0(N__7189),
            .in1(N__5122),
            .in2(N__6148),
            .in3(N__5180),
            .lcout(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.LW_CYCLE_STARTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A_OUT_RNO_0_LC_13_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A_OUT_RNO_0_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A_OUT_RNO_0_LC_13_13_1 .LUT_INIT=16'b1100110010101110;
    LogicCell40 \U111_CYCLE_SM.A_OUT_RNO_0_LC_13_13_1  (
            .in0(N__6198),
            .in1(N__4386),
            .in2(N__5182),
            .in3(N__6247),
            .lcout(),
            .ltout(\U111_CYCLE_SM.A_OUT_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A_OUT_LC_13_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A_OUT_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.A_OUT_LC_13_13_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U111_CYCLE_SM.A_OUT_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4399),
            .in3(N__6129),
            .lcout(\U111_CYCLE_SM.A_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.LW_CYCLE_STARTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_13_13_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_13_13_3 .LUT_INIT=16'b1011101110011001;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_0_LC_13_13_3  (
            .in0(N__6197),
            .in1(N__6246),
            .in2(_gnd_net_),
            .in3(N__5687),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_75_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_LC_13_13_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_LC_13_13_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TS_EN_LC_13_13_4 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \U111_CYCLE_SM.TS_EN_LC_13_13_4  (
            .in0(N__5139),
            .in1(N__6130),
            .in2(N__4375),
            .in3(N__4564),
            .lcout(\U111_CYCLE_SM.TS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.LW_CYCLE_STARTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_EN_RNO_0_LC_13_13_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_EN_RNO_0_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_EN_RNO_0_LC_13_13_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \U111_CYCLE_SM.TA_EN_RNO_0_LC_13_13_6  (
            .in0(N__6137),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.RESETn_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_13_13_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_13_13_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_13_13_7  (
            .in0(N__5064),
            .in1(N__5037),
            .in2(N__5871),
            .in3(N__5138),
            .lcout(\U111_CYCLE_SM.un3_LW_CYCLE_START ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_EN_LC_13_14_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_EN_LC_13_14_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.TA_EN_LC_13_14_6 .LUT_INIT=16'b1111000011011100;
    LogicCell40 \U111_CYCLE_SM.TA_EN_LC_13_14_6  (
            .in0(N__5181),
            .in1(N__6201),
            .in2(N__5903),
            .in3(N__6248),
            .lcout(\U111_CYCLE_SM.TA_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TA_ENC_net ),
            .ce(),
            .sr(N__5116));
    defparam \U111_CYCLE_SM.LW_TRANS_LC_13_16_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_13_16_0 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \U111_CYCLE_SM.LW_TRANS_LC_13_16_0  (
            .in0(N__5104),
            .in1(N__5086),
            .in2(_gnd_net_),
            .in3(N__5068),
            .lcout(\U111_CYCLE_SM.LW_TRANS_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_13_16_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_13_16_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_13_16_4  (
            .in0(N__5625),
            .in1(N__4820),
            .in2(_gnd_net_),
            .in3(N__5020),
            .lcout(un1_D_LM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_13_20_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_13_20_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_13_20_0  (
            .in0(N__4980),
            .in1(N__4813),
            .in2(_gnd_net_),
            .in3(N__4933),
            .lcout(un1_D_UM_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_13_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_13_20_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_13_20_2  (
            .in0(N__4900),
            .in1(N__4812),
            .in2(_gnd_net_),
            .in3(N__4650),
            .lcout(un1_D_UU_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_EN_RNI4SHG_LC_14_1_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_EN_RNI4SHG_LC_14_1_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_EN_RNI4SHG_LC_14_1_2 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U111_CYCLE_SM.TA_EN_RNI4SHG_LC_14_1_2  (
            .in0(N__5911),
            .in1(N__6275),
            .in2(_gnd_net_),
            .in3(N__5850),
            .lcout(U111_CYCLE_SM_TBI_CPUn_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_14_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_14_13_1 .LUT_INIT=16'b0001101100001010;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_1_LC_14_13_1  (
            .in0(N__6192),
            .in1(N__5479),
            .in2(N__6250),
            .in3(N__5647),
            .lcout(\U111_CYCLE_SM.TS_EN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CPU_READ_EN_i_LC_14_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CPU_READ_EN_i_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CPU_READ_EN_i_LC_14_13_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U111_CYCLE_SM.CPU_READ_EN_i_LC_14_13_2  (
            .in0(N__5478),
            .in1(N__6045),
            .in2(_gnd_net_),
            .in3(N__5866),
            .lcout(CPU_READ_EN_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_14_13_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_14_13_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_14_13_5 .LUT_INIT=16'b1001000010100000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_1_LC_14_13_5  (
            .in0(N__6193),
            .in1(N__6282),
            .in2(N__6154),
            .in3(N__6249),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.CYCLE_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_14_14_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_14_14_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__5175),
            .in2(_gnd_net_),
            .in3(N__6241),
            .lcout(),
            .ltout(\U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_LC_14_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_CYCLE_LC_14_14_1 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_LC_14_14_1  (
            .in0(N__6152),
            .in1(N__5152),
            .in2(N__5185),
            .in3(N__6200),
            .lcout(\U111_CYCLE_SM.LW_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.LW_CYCLEC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_14_14_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_14_14_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_14_14_4  (
            .in0(N__6199),
            .in1(N__5176),
            .in2(_gnd_net_),
            .in3(N__5688),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_97_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_14_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_14_14_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_14_14_5 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_0_LC_14_14_5  (
            .in0(N__6242),
            .in1(N__6301),
            .in2(N__5155),
            .in3(N__6147),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.LW_CYCLEC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_14_14_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_14_14_7 .LUT_INIT=16'b1100110001001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_14_14_7  (
            .in0(N__6240),
            .in1(N__7188),
            .in2(N__6202),
            .in3(N__6302),
            .lcout(\U111_CYCLE_SM.LW_CYCLE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_14_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_14_15_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_14_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5547),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net ),
            .ce(N__7045),
            .sr(N__7005));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_14_15_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_14_15_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_14_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5621),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net ),
            .ce(N__7045),
            .sr(N__7005));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_14_15_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_14_15_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_14_15_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_14_15_3  (
            .in0(N__5973),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net ),
            .ce(N__7045),
            .sr(N__7005));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_14_15_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_14_15_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_14_15_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_14_15_7  (
            .in0(N__5766),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net ),
            .ce(N__7045),
            .sr(N__7005));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_14_16_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_14_16_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_14_16_0  (
            .in0(N__7228),
            .in1(N__5983),
            .in2(_gnd_net_),
            .in3(N__5972),
            .lcout(un1_D_UU_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_EN_RNIVCEG_LC_14_16_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_EN_RNIVCEG_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_EN_RNIVCEG_LC_14_16_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.TA_EN_RNIVCEG_LC_14_16_4  (
            .in0(N__5904),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5878),
            .lcout(TAn_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_14_16_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_14_16_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_14_16_5  (
            .in0(N__5753),
            .in1(N__5725),
            .in2(_gnd_net_),
            .in3(N__7227),
            .lcout(un1_D_UM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_2_LC_14_18_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_2_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_2_LC_14_18_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_2_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__5701),
            .in2(_gnd_net_),
            .in3(N__5686),
            .lcout(\U111_CYCLE_SM.TS_EN_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_14_18_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_14_18_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_14_18_6  (
            .in0(N__7230),
            .in1(N__5635),
            .in2(_gnd_net_),
            .in3(N__5626),
            .lcout(un1_D_UU_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_14_18_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_14_18_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_14_18_7  (
            .in0(N__5557),
            .in1(N__5543),
            .in2(_gnd_net_),
            .in3(N__7229),
            .lcout(un1_D_UU_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_15_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_15_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_15_11_0  (
            .in0(N__6424),
            .in1(N__6459),
            .in2(_gnd_net_),
            .in3(N__7249),
            .lcout(un1_D_UM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_15_11_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_15_11_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_15_11_5  (
            .in0(N__7250),
            .in1(N__6325),
            .in2(_gnd_net_),
            .in3(N__6360),
            .lcout(un1_D_UM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_15_12_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_15_12_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_15_12_1  (
            .in0(N__6373),
            .in1(N__6401),
            .in2(_gnd_net_),
            .in3(N__7248),
            .lcout(un1_D_UM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_15_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_15_13_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_15_13_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_15_13_1  (
            .in0(N__6458),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net ),
            .ce(N__7036),
            .sr(N__7003));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_15_13_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_15_13_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_15_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6411),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net ),
            .ce(N__7036),
            .sr(N__7003));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_15_13_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_15_13_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_15_13_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_15_13_6  (
            .in0(N__6359),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net ),
            .ce(N__7036),
            .sr(N__7003));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIULFD_0_LC_15_14_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIULFD_0_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIULFD_0_LC_15_14_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIULFD_0_LC_15_14_4  (
            .in0(N__6303),
            .in1(N__6239),
            .in2(_gnd_net_),
            .in3(N__6191),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa ),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1_0_LC_15_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1_0_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1_0_LC_15_14_5 .LUT_INIT=16'b0011001111110011;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1_0_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(N__6153),
            .in2(N__6055),
            .in3(N__6037),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0 ),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIE3PP1_0_LC_15_14_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIE3PP1_0_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIE3PP1_0_LC_15_14_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIE3PP1_0_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5992),
            .in3(N__5989),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_15_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_15_15_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_15_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7119),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__7044),
            .sr(N__7004));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_15_15_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_15_15_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_15_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6764),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__7044),
            .sr(N__7004));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_15_15_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_15_15_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_15_15_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_15_15_4  (
            .in0(N__6694),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__7044),
            .sr(N__7004));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_15_15_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_15_15_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_15_15_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_15_15_6  (
            .in0(N__6630),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__7044),
            .sr(N__7004));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_15_15_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_15_15_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_15_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6562),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__7044),
            .sr(N__7004));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_15_16_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_15_16_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_15_16_0  (
            .in0(N__7231),
            .in1(N__6778),
            .in2(_gnd_net_),
            .in3(N__6771),
            .lcout(un1_D_UM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_15_16_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_15_16_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_15_16_2  (
            .in0(N__7232),
            .in1(N__6700),
            .in2(_gnd_net_),
            .in3(N__6693),
            .lcout(un1_D_UU_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_15_16_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_15_16_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_15_16_6  (
            .in0(N__7233),
            .in1(N__6640),
            .in2(_gnd_net_),
            .in3(N__6629),
            .lcout(un1_D_UU_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_15_18_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_15_18_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_15_18_2  (
            .in0(N__7262),
            .in1(N__6571),
            .in2(_gnd_net_),
            .in3(N__6561),
            .lcout(un1_D_UU_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_15_18_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_15_18_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_15_18_7  (
            .in0(N__7112),
            .in1(N__7075),
            .in2(_gnd_net_),
            .in3(N__7261),
            .lcout(un1_D_UM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_16_15_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_16_15_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_16_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7320),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net ),
            .ce(N__7043),
            .sr(N__7006));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_16_15_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_16_15_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_16_15_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_16_15_2  (
            .in0(N__6841),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net ),
            .ce(N__7043),
            .sr(N__7006));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_16_15_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_16_15_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_16_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6906),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net ),
            .ce(N__7043),
            .sr(N__7006));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_16_15_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_16_15_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_16_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6976),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net ),
            .ce(N__7043),
            .sr(N__7006));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_16_16_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_16_16_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_16_16_0  (
            .in0(N__7258),
            .in1(N__6982),
            .in2(_gnd_net_),
            .in3(N__6975),
            .lcout(un1_D_UM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_16_16_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_16_16_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_16_16_2  (
            .in0(N__7260),
            .in1(N__6916),
            .in2(_gnd_net_),
            .in3(N__6905),
            .lcout(un1_D_UU_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_16_16_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_16_16_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_16_16_3  (
            .in0(N__6847),
            .in1(N__6837),
            .in2(_gnd_net_),
            .in3(N__7259),
            .lcout(un1_D_UU_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_16_16_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_16_16_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_16_16_7  (
            .in0(N__7330),
            .in1(N__7319),
            .in2(_gnd_net_),
            .in3(N__7257),
            .lcout(un1_D_UM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U111_TOP

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 25 2025 21:58:51

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    TT,
    A,
    TICK50,
    nROMEN,
    nCIACS1,
    TICK60,
    CLKCIA,
    CLK6,
    CLK40_IN,
    CLK28_IN,
    TSn,
    nBUFEN,
    nREGSPACE,
    nRAMSPACE,
    RESETn,
    OVL,
    TACKn,
    nCIACS0,
    PORTSIZE);

    input [1:0] TT;
    input [31:1] A;
    output TICK50;
    output nROMEN;
    output nCIACS1;
    output TICK60;
    output CLKCIA;
    input CLK6;
    input CLK40_IN;
    input CLK28_IN;
    input TSn;
    output nBUFEN;
    output nREGSPACE;
    output nRAMSPACE;
    input RESETn;
    input OVL;
    inout TACKn;
    output nCIACS0;
    output PORTSIZE;

    wire N__6546;
    wire N__6545;
    wire N__6544;
    wire N__6536;
    wire N__6535;
    wire N__6534;
    wire N__6525;
    wire N__6524;
    wire N__6523;
    wire N__6516;
    wire N__6515;
    wire N__6514;
    wire N__6507;
    wire N__6506;
    wire N__6505;
    wire N__6498;
    wire N__6497;
    wire N__6496;
    wire N__6489;
    wire N__6488;
    wire N__6487;
    wire N__6480;
    wire N__6479;
    wire N__6478;
    wire N__6471;
    wire N__6470;
    wire N__6469;
    wire N__6462;
    wire N__6461;
    wire N__6460;
    wire N__6453;
    wire N__6452;
    wire N__6451;
    wire N__6444;
    wire N__6443;
    wire N__6442;
    wire N__6435;
    wire N__6434;
    wire N__6433;
    wire N__6426;
    wire N__6425;
    wire N__6424;
    wire N__6417;
    wire N__6416;
    wire N__6415;
    wire N__6408;
    wire N__6407;
    wire N__6406;
    wire N__6399;
    wire N__6398;
    wire N__6397;
    wire N__6390;
    wire N__6389;
    wire N__6388;
    wire N__6381;
    wire N__6380;
    wire N__6379;
    wire N__6372;
    wire N__6371;
    wire N__6370;
    wire N__6363;
    wire N__6362;
    wire N__6361;
    wire N__6354;
    wire N__6353;
    wire N__6352;
    wire N__6345;
    wire N__6344;
    wire N__6343;
    wire N__6336;
    wire N__6335;
    wire N__6334;
    wire N__6327;
    wire N__6326;
    wire N__6325;
    wire N__6318;
    wire N__6317;
    wire N__6316;
    wire N__6309;
    wire N__6308;
    wire N__6307;
    wire N__6300;
    wire N__6299;
    wire N__6298;
    wire N__6291;
    wire N__6290;
    wire N__6289;
    wire N__6282;
    wire N__6281;
    wire N__6280;
    wire N__6273;
    wire N__6272;
    wire N__6271;
    wire N__6264;
    wire N__6263;
    wire N__6262;
    wire N__6255;
    wire N__6254;
    wire N__6253;
    wire N__6246;
    wire N__6245;
    wire N__6244;
    wire N__6237;
    wire N__6236;
    wire N__6235;
    wire N__6228;
    wire N__6227;
    wire N__6226;
    wire N__6219;
    wire N__6218;
    wire N__6217;
    wire N__6200;
    wire N__6199;
    wire N__6198;
    wire N__6195;
    wire N__6188;
    wire N__6185;
    wire N__6184;
    wire N__6183;
    wire N__6176;
    wire N__6173;
    wire N__6172;
    wire N__6169;
    wire N__6166;
    wire N__6161;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6151;
    wire N__6148;
    wire N__6147;
    wire N__6144;
    wire N__6141;
    wire N__6138;
    wire N__6135;
    wire N__6132;
    wire N__6127;
    wire N__6126;
    wire N__6125;
    wire N__6120;
    wire N__6117;
    wire N__6116;
    wire N__6113;
    wire N__6112;
    wire N__6111;
    wire N__6110;
    wire N__6109;
    wire N__6108;
    wire N__6107;
    wire N__6106;
    wire N__6103;
    wire N__6098;
    wire N__6093;
    wire N__6090;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6080;
    wire N__6075;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6050;
    wire N__6041;
    wire N__6038;
    wire N__6035;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6001;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5984;
    wire N__5983;
    wire N__5980;
    wire N__5977;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5957;
    wire N__5954;
    wire N__5951;
    wire N__5948;
    wire N__5947;
    wire N__5944;
    wire N__5943;
    wire N__5940;
    wire N__5937;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5903;
    wire N__5900;
    wire N__5897;
    wire N__5894;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5866;
    wire N__5865;
    wire N__5864;
    wire N__5863;
    wire N__5862;
    wire N__5861;
    wire N__5856;
    wire N__5849;
    wire N__5844;
    wire N__5837;
    wire N__5834;
    wire N__5831;
    wire N__5830;
    wire N__5829;
    wire N__5826;
    wire N__5823;
    wire N__5822;
    wire N__5819;
    wire N__5814;
    wire N__5811;
    wire N__5804;
    wire N__5803;
    wire N__5802;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5790;
    wire N__5783;
    wire N__5782;
    wire N__5781;
    wire N__5780;
    wire N__5775;
    wire N__5772;
    wire N__5769;
    wire N__5762;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5750;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5742;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5723;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5710;
    wire N__5707;
    wire N__5704;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5692;
    wire N__5687;
    wire N__5684;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5676;
    wire N__5675;
    wire N__5674;
    wire N__5673;
    wire N__5668;
    wire N__5665;
    wire N__5662;
    wire N__5659;
    wire N__5658;
    wire N__5655;
    wire N__5648;
    wire N__5645;
    wire N__5644;
    wire N__5641;
    wire N__5638;
    wire N__5633;
    wire N__5630;
    wire N__5627;
    wire N__5624;
    wire N__5621;
    wire N__5616;
    wire N__5613;
    wire N__5610;
    wire N__5607;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5593;
    wire N__5590;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5577;
    wire N__5574;
    wire N__5571;
    wire N__5568;
    wire N__5563;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5528;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5482;
    wire N__5481;
    wire N__5480;
    wire N__5479;
    wire N__5478;
    wire N__5477;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5463;
    wire N__5454;
    wire N__5447;
    wire N__5444;
    wire N__5443;
    wire N__5442;
    wire N__5441;
    wire N__5440;
    wire N__5439;
    wire N__5436;
    wire N__5429;
    wire N__5424;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5403;
    wire N__5400;
    wire N__5397;
    wire N__5394;
    wire N__5387;
    wire N__5386;
    wire N__5385;
    wire N__5384;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5347;
    wire N__5346;
    wire N__5345;
    wire N__5344;
    wire N__5337;
    wire N__5332;
    wire N__5327;
    wire N__5326;
    wire N__5325;
    wire N__5324;
    wire N__5323;
    wire N__5316;
    wire N__5311;
    wire N__5306;
    wire N__5305;
    wire N__5304;
    wire N__5301;
    wire N__5300;
    wire N__5297;
    wire N__5296;
    wire N__5289;
    wire N__5284;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5269;
    wire N__5268;
    wire N__5267;
    wire N__5266;
    wire N__5265;
    wire N__5264;
    wire N__5261;
    wire N__5256;
    wire N__5253;
    wire N__5246;
    wire N__5237;
    wire N__5236;
    wire N__5235;
    wire N__5234;
    wire N__5233;
    wire N__5232;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5218;
    wire N__5213;
    wire N__5204;
    wire N__5203;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5195;
    wire N__5194;
    wire N__5193;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5180;
    wire N__5175;
    wire N__5170;
    wire N__5167;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5146;
    wire N__5143;
    wire N__5140;
    wire N__5137;
    wire N__5134;
    wire N__5129;
    wire N__5128;
    wire N__5127;
    wire N__5126;
    wire N__5125;
    wire N__5124;
    wire N__5123;
    wire N__5122;
    wire N__5121;
    wire N__5120;
    wire N__5119;
    wire N__5118;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5071;
    wire N__5070;
    wire N__5067;
    wire N__5062;
    wire N__5057;
    wire N__5054;
    wire N__5053;
    wire N__5050;
    wire N__5049;
    wire N__5048;
    wire N__5045;
    wire N__5040;
    wire N__5037;
    wire N__5030;
    wire N__5029;
    wire N__5026;
    wire N__5025;
    wire N__5020;
    wire N__5017;
    wire N__5014;
    wire N__5011;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4990;
    wire N__4989;
    wire N__4986;
    wire N__4981;
    wire N__4976;
    wire N__4975;
    wire N__4974;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4960;
    wire N__4955;
    wire N__4954;
    wire N__4953;
    wire N__4952;
    wire N__4951;
    wire N__4948;
    wire N__4939;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4924;
    wire N__4923;
    wire N__4922;
    wire N__4919;
    wire N__4912;
    wire N__4907;
    wire N__4904;
    wire N__4903;
    wire N__4902;
    wire N__4895;
    wire N__4892;
    wire N__4891;
    wire N__4890;
    wire N__4887;
    wire N__4882;
    wire N__4877;
    wire N__4876;
    wire N__4871;
    wire N__4868;
    wire N__4867;
    wire N__4864;
    wire N__4861;
    wire N__4858;
    wire N__4853;
    wire N__4852;
    wire N__4849;
    wire N__4846;
    wire N__4841;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4829;
    wire N__4828;
    wire N__4825;
    wire N__4822;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4810;
    wire N__4807;
    wire N__4804;
    wire N__4799;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4774;
    wire N__4771;
    wire N__4768;
    wire N__4763;
    wire N__4762;
    wire N__4759;
    wire N__4756;
    wire N__4751;
    wire N__4750;
    wire N__4747;
    wire N__4744;
    wire N__4739;
    wire N__4738;
    wire N__4737;
    wire N__4736;
    wire N__4733;
    wire N__4730;
    wire N__4725;
    wire N__4722;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4697;
    wire N__4694;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4672;
    wire N__4669;
    wire N__4666;
    wire N__4661;
    wire N__4660;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4571;
    wire N__4570;
    wire N__4567;
    wire N__4564;
    wire N__4559;
    wire N__4558;
    wire N__4555;
    wire N__4552;
    wire N__4547;
    wire N__4546;
    wire N__4543;
    wire N__4542;
    wire N__4537;
    wire N__4534;
    wire N__4529;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4480;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4468;
    wire N__4465;
    wire N__4464;
    wire N__4461;
    wire N__4460;
    wire N__4459;
    wire N__4458;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4445;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4420;
    wire N__4417;
    wire N__4412;
    wire N__4405;
    wire N__4402;
    wire N__4399;
    wire N__4394;
    wire N__4393;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4385;
    wire N__4384;
    wire N__4381;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4371;
    wire N__4368;
    wire N__4367;
    wire N__4366;
    wire N__4365;
    wire N__4362;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4321;
    wire N__4316;
    wire N__4309;
    wire N__4304;
    wire N__4301;
    wire N__4300;
    wire N__4297;
    wire N__4296;
    wire N__4293;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4282;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4261;
    wire N__4258;
    wire N__4255;
    wire N__4248;
    wire N__4245;
    wire N__4240;
    wire N__4235;
    wire N__4232;
    wire N__4229;
    wire N__4228;
    wire N__4225;
    wire N__4222;
    wire N__4217;
    wire N__4214;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4150;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4114;
    wire N__4111;
    wire N__4110;
    wire N__4107;
    wire N__4106;
    wire N__4105;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4093;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4075;
    wire N__4072;
    wire N__4065;
    wire N__4062;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4037;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4025;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire N__3983;
    wire N__3982;
    wire N__3979;
    wire N__3976;
    wire N__3973;
    wire N__3972;
    wire N__3971;
    wire N__3970;
    wire N__3969;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3951;
    wire N__3944;
    wire N__3943;
    wire N__3942;
    wire N__3941;
    wire N__3940;
    wire N__3937;
    wire N__3934;
    wire N__3927;
    wire N__3920;
    wire N__3919;
    wire N__3918;
    wire N__3917;
    wire N__3914;
    wire N__3911;
    wire N__3906;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3892;
    wire N__3891;
    wire N__3888;
    wire N__3883;
    wire N__3878;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3847;
    wire N__3844;
    wire N__3843;
    wire N__3840;
    wire N__3837;
    wire N__3834;
    wire N__3827;
    wire N__3826;
    wire N__3825;
    wire N__3824;
    wire N__3821;
    wire N__3818;
    wire N__3815;
    wire N__3812;
    wire N__3803;
    wire N__3802;
    wire N__3801;
    wire N__3798;
    wire N__3797;
    wire N__3792;
    wire N__3787;
    wire N__3782;
    wire N__3781;
    wire N__3780;
    wire N__3777;
    wire N__3776;
    wire N__3773;
    wire N__3770;
    wire N__3767;
    wire N__3764;
    wire N__3761;
    wire N__3756;
    wire N__3749;
    wire N__3748;
    wire N__3747;
    wire N__3746;
    wire N__3745;
    wire N__3742;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3728;
    wire N__3723;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3709;
    wire N__3704;
    wire N__3701;
    wire N__3698;
    wire N__3697;
    wire N__3694;
    wire N__3693;
    wire N__3692;
    wire N__3689;
    wire N__3688;
    wire N__3683;
    wire N__3676;
    wire N__3671;
    wire N__3668;
    wire N__3665;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3637;
    wire N__3636;
    wire N__3633;
    wire N__3630;
    wire N__3627;
    wire N__3624;
    wire N__3621;
    wire N__3618;
    wire N__3611;
    wire N__3608;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire N__3596;
    wire N__3593;
    wire N__3590;
    wire N__3587;
    wire N__3584;
    wire N__3581;
    wire N__3578;
    wire N__3575;
    wire N__3572;
    wire N__3569;
    wire N__3566;
    wire N__3563;
    wire N__3560;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3548;
    wire N__3547;
    wire N__3546;
    wire N__3545;
    wire N__3544;
    wire N__3543;
    wire N__3542;
    wire N__3533;
    wire N__3530;
    wire N__3529;
    wire N__3526;
    wire N__3523;
    wire N__3520;
    wire N__3515;
    wire N__3506;
    wire N__3503;
    wire N__3502;
    wire N__3501;
    wire N__3500;
    wire N__3499;
    wire N__3498;
    wire N__3497;
    wire N__3496;
    wire N__3493;
    wire N__3486;
    wire N__3483;
    wire N__3476;
    wire N__3467;
    wire N__3466;
    wire N__3465;
    wire N__3464;
    wire N__3461;
    wire N__3460;
    wire N__3457;
    wire N__3454;
    wire N__3451;
    wire N__3450;
    wire N__3449;
    wire N__3448;
    wire N__3445;
    wire N__3442;
    wire N__3435;
    wire N__3432;
    wire N__3427;
    wire N__3416;
    wire N__3413;
    wire N__3410;
    wire N__3407;
    wire N__3406;
    wire N__3403;
    wire N__3400;
    wire N__3397;
    wire N__3392;
    wire N__3391;
    wire N__3386;
    wire N__3383;
    wire N__3380;
    wire N__3377;
    wire N__3374;
    wire N__3373;
    wire N__3368;
    wire N__3365;
    wire N__3362;
    wire N__3359;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3347;
    wire N__3344;
    wire N__3341;
    wire N__3340;
    wire N__3337;
    wire N__3334;
    wire N__3329;
    wire N__3326;
    wire N__3323;
    wire N__3320;
    wire N__3319;
    wire N__3316;
    wire N__3313;
    wire N__3312;
    wire N__3307;
    wire N__3304;
    wire N__3299;
    wire N__3298;
    wire N__3297;
    wire N__3296;
    wire N__3293;
    wire N__3286;
    wire N__3283;
    wire N__3278;
    wire N__3275;
    wire N__3272;
    wire N__3269;
    wire N__3268;
    wire N__3265;
    wire N__3262;
    wire N__3257;
    wire N__3254;
    wire N__3251;
    wire N__3250;
    wire N__3247;
    wire N__3244;
    wire N__3239;
    wire N__3236;
    wire N__3233;
    wire N__3230;
    wire N__3229;
    wire N__3226;
    wire N__3223;
    wire N__3218;
    wire N__3215;
    wire N__3212;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3200;
    wire N__3197;
    wire N__3194;
    wire N__3193;
    wire N__3190;
    wire N__3187;
    wire N__3182;
    wire N__3179;
    wire N__3176;
    wire N__3173;
    wire N__3170;
    wire N__3167;
    wire N__3166;
    wire N__3163;
    wire N__3160;
    wire N__3155;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3143;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3131;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3119;
    wire N__3118;
    wire N__3115;
    wire N__3112;
    wire N__3107;
    wire N__3104;
    wire N__3101;
    wire N__3098;
    wire N__3097;
    wire N__3094;
    wire N__3091;
    wire N__3086;
    wire N__3085;
    wire N__3082;
    wire N__3079;
    wire N__3074;
    wire N__3071;
    wire N__3068;
    wire N__3065;
    wire N__3062;
    wire N__3059;
    wire N__3056;
    wire N__3053;
    wire N__3050;
    wire N__3047;
    wire N__3044;
    wire N__3043;
    wire N__3038;
    wire N__3037;
    wire N__3034;
    wire N__3031;
    wire N__3026;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3013;
    wire N__3010;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__3000;
    wire N__2999;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2981;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2966;
    wire N__2963;
    wire N__2960;
    wire N__2957;
    wire N__2954;
    wire N__2951;
    wire N__2948;
    wire N__2945;
    wire N__2942;
    wire N__2939;
    wire N__2936;
    wire N__2933;
    wire N__2930;
    wire N__2927;
    wire N__2924;
    wire N__2921;
    wire N__2918;
    wire N__2915;
    wire N__2912;
    wire N__2909;
    wire N__2906;
    wire N__2903;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2890;
    wire N__2889;
    wire N__2886;
    wire N__2883;
    wire N__2880;
    wire N__2877;
    wire N__2872;
    wire N__2869;
    wire N__2866;
    wire N__2863;
    wire N__2860;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2842;
    wire N__2841;
    wire N__2838;
    wire N__2833;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2819;
    wire N__2816;
    wire N__2813;
    wire N__2810;
    wire N__2809;
    wire N__2808;
    wire N__2805;
    wire N__2800;
    wire N__2795;
    wire N__2792;
    wire N__2789;
    wire N__2788;
    wire N__2785;
    wire N__2784;
    wire N__2781;
    wire N__2778;
    wire N__2773;
    wire N__2768;
    wire N__2765;
    wire N__2764;
    wire N__2763;
    wire N__2760;
    wire N__2755;
    wire N__2750;
    wire N__2747;
    wire N__2744;
    wire N__2741;
    wire N__2738;
    wire N__2735;
    wire N__2732;
    wire N__2729;
    wire N__2728;
    wire N__2727;
    wire N__2720;
    wire N__2717;
    wire N__2714;
    wire N__2711;
    wire N__2708;
    wire N__2707;
    wire N__2706;
    wire N__2699;
    wire N__2696;
    wire N__2693;
    wire N__2690;
    wire N__2687;
    wire N__2684;
    wire N__2683;
    wire N__2680;
    wire N__2677;
    wire N__2676;
    wire N__2673;
    wire N__2668;
    wire N__2663;
    wire N__2660;
    wire N__2657;
    wire N__2654;
    wire N__2653;
    wire N__2650;
    wire N__2649;
    wire N__2646;
    wire N__2639;
    wire N__2636;
    wire N__2633;
    wire N__2630;
    wire N__2627;
    wire N__2624;
    wire N__2621;
    wire N__2618;
    wire N__2615;
    wire N__2612;
    wire N__2609;
    wire N__2608;
    wire N__2605;
    wire N__2602;
    wire N__2597;
    wire N__2594;
    wire N__2591;
    wire N__2588;
    wire N__2585;
    wire N__2582;
    wire N__2579;
    wire N__2576;
    wire N__2573;
    wire N__2570;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2558;
    wire N__2555;
    wire N__2554;
    wire N__2551;
    wire N__2548;
    wire N__2545;
    wire N__2540;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2525;
    wire N__2524;
    wire N__2519;
    wire N__2516;
    wire N__2513;
    wire N__2510;
    wire N__2507;
    wire N__2504;
    wire N__2503;
    wire N__2502;
    wire N__2501;
    wire N__2500;
    wire N__2499;
    wire N__2498;
    wire N__2497;
    wire N__2496;
    wire N__2495;
    wire N__2474;
    wire CLK80_OUT;
    wire GNDG0;
    wire VCCG0;
    wire A_c_18;
    wire A_c_17;
    wire \U409_CIA.g0Z0Z_2_cascade_ ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_ ;
    wire A_c_26;
    wire A_c_27;
    wire A_c_25;
    wire A_c_24;
    wire \U409_CIA.g0Z0Z_10 ;
    wire A_c_31;
    wire A_c_28;
    wire A_c_30;
    wire A_c_29;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ;
    wire \U409_CIA.g0Z0Z_8 ;
    wire A_c_16;
    wire \U409_CIA.g0Z0Z_11 ;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8 ;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEm_3_cascade_ ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEm_6 ;
    wire A_c_20;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_0 ;
    wire TT_c_1;
    wire TT_c_0;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACE_1Z0Z_0 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEm_cascade_ ;
    wire PORTSIZE_0_i;
    wire \U409_ADDRESS_DECODE.CIA_SPACEm_3 ;
    wire A_c_19;
    wire bfn_8_5_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire bfn_8_6_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.TICK503_11 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire TICK50_c;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ;
    wire U409_ADDRESS_DECODE_un1_nREGSPACE_i;
    wire bfn_11_5_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire bfn_11_6_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.m9_am_cascade_ ;
    wire \U409_TRANSFER_ACK.i6_mux_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire \U409_TRANSFER_ACK.N_105_cascade_ ;
    wire \U409_TRANSFER_ACK.m9_bm ;
    wire \U409_TRANSFER_ACK.N_4 ;
    wire A_c_22;
    wire A_c_23;
    wire A_c_21;
    wire \U409_ADDRESS_DECODE.LOWROMZ0 ;
    wire \U409_ADDRESS_DECODE.HIROMZ0 ;
    wire ROMENm_i;
    wire AUTOVECTORm;
    wire TSn_c;
    wire CLK40_IN_c;
    wire ROMENm;
    wire CONSTANT_ONE_NET;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_nCIACS0_i;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_nCIACS1_i;
    wire U409_ADDRESS_DECODE_un1_nRAMSPACE_i;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire TICK60_c;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.TICK603_10_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire \U409_TICK.TICK603_11 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.TICK603_8_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire CIA_ENABLEm;
    wire \U409_CIA.N_9_cascade_ ;
    wire \U409_CIA.g0Z0Z_14 ;
    wire \U409_CIA.VMAZ0 ;
    wire \U409_CIA.g0Z0Z_13 ;
    wire \U409_CIA.CIA_HOLDZ0 ;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_105 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_0C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire CLK6_c_g;
    wire bfn_13_7_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a2_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_ ;
    wire \U409_CIA.N_20_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CLKCIAZ0_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire CLKCIA_c;
    wire CLK28_IN_c_g;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.CLKCIA6_0_a2_1 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CLKCIA8_0_a2_0 ;
    wire RESETn_c_i;
    wire \U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ;
    wire \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0 ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0 ;
    wire OVL_c;
    wire TACK_OUTn;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER5_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ;
    wire \INVU409_TRANSFER_ACK.TACK_EN_iC_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ;
    wire RESETn_c;
    wire nBUFEN_c;
    wire TACKn_in;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire TACK_EN_i;
    wire N_365_i;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__4118),
            .RESETB(N__4040),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6544),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__6546),
            .DIN(N__6545),
            .DOUT(N__6544),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__6546),
            .PADOUT(N__6545),
            .PADIN(N__6544),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6534),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__6536),
            .DIN(N__6535),
            .DOUT(N__6534),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__6536),
            .PADOUT(N__6535),
            .PADIN(N__6534),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__6525),
            .DIN(N__6524),
            .DOUT(N__6523),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__6525),
            .PADOUT(N__6524),
            .PADIN(N__6523),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKCIA_obuf_iopad (
            .OE(N__6516),
            .DIN(N__6515),
            .DOUT(N__6514),
            .PACKAGEPIN(CLKCIA));
    defparam CLKCIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKCIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKCIA_obuf_preio (
            .PADOEN(N__6516),
            .PADOUT(N__6515),
            .PADIN(N__6514),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5417),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_24_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_24_iopad (
            .OE(N__6507),
            .DIN(N__6506),
            .DOUT(N__6505),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__6507),
            .PADOUT(N__6506),
            .PADIN(N__6505),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nCIACS0_obuf_iopad (
            .OE(N__6498),
            .DIN(N__6497),
            .DOUT(N__6496),
            .PACKAGEPIN(nCIACS0));
    defparam nCIACS0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCIACS0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCIACS0_obuf_preio (
            .PADOEN(N__6498),
            .PADOUT(N__6497),
            .PADIN(N__6496),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4010),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nCIACS1_obuf_iopad (
            .OE(N__6489),
            .DIN(N__6488),
            .DOUT(N__6487),
            .PACKAGEPIN(nCIACS1));
    defparam nCIACS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCIACS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCIACS1_obuf_preio (
            .PADOEN(N__6489),
            .PADOUT(N__6488),
            .PADIN(N__6487),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4628),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_31_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_31_iopad (
            .OE(N__6480),
            .DIN(N__6479),
            .DOUT(N__6478),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__6480),
            .PADOUT(N__6479),
            .PADIN(N__6478),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_17_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_17_iopad (
            .OE(N__6471),
            .DIN(N__6470),
            .DOUT(N__6469),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__6471),
            .PADOUT(N__6470),
            .PADIN(N__6469),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_21_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_21_iopad (
            .OE(N__6462),
            .DIN(N__6461),
            .DOUT(N__6460),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__6462),
            .PADOUT(N__6461),
            .PADIN(N__6460),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_iobuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__6453),
            .DIN(N__6452),
            .DOUT(N__6451),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__6453),
            .PADOUT(N__6452),
            .PADIN(N__6451),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5885),
            .DIN0(TACKn_in),
            .DOUT0(N__5555),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_12_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_12_iopad (
            .OE(N__6444),
            .DIN(N__6443),
            .DOUT(N__6442),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__6444),
            .PADOUT(N__6443),
            .PADIN(N__6442),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__6435),
            .DIN(N__6434),
            .DOUT(N__6433),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__6435),
            .PADOUT(N__6434),
            .PADIN(N__6433),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__6426),
            .DIN(N__6425),
            .DOUT(N__6424),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__6426),
            .PADOUT(N__6425),
            .PADIN(N__6424),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PORTSIZE_obuf_iopad.PULLUP=1'b1;
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__6417),
            .DIN(N__6416),
            .DOUT(N__6415),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__6417),
            .PADOUT(N__6416),
            .PADIN(N__6415),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2909),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nRAMSPACE_obuf_iopad (
            .OE(N__6408),
            .DIN(N__6407),
            .DOUT(N__6406),
            .PACKAGEPIN(nRAMSPACE));
    defparam nRAMSPACE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nRAMSPACE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nRAMSPACE_obuf_preio (
            .PADOEN(N__6408),
            .PADOUT(N__6407),
            .PADIN(N__6406),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4613),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nROMEN_obuf_iopad (
            .OE(N__6399),
            .DIN(N__6398),
            .DOUT(N__6397),
            .PACKAGEPIN(nROMEN));
    defparam nROMEN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nROMEN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nROMEN_obuf_preio (
            .PADOEN(N__6399),
            .PADOUT(N__6398),
            .PADIN(N__6397),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4187),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_18_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_18_iopad (
            .OE(N__6390),
            .DIN(N__6389),
            .DOUT(N__6388),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__6390),
            .PADOUT(N__6389),
            .PADIN(N__6388),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_29_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_29_iopad (
            .OE(N__6381),
            .DIN(N__6380),
            .DOUT(N__6379),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__6381),
            .PADOUT(N__6380),
            .PADIN(N__6379),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nBUFEN_obuf_iopad (
            .OE(N__6372),
            .DIN(N__6371),
            .DOUT(N__6370),
            .PACKAGEPIN(nBUFEN));
    defparam nBUFEN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nBUFEN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nBUFEN_obuf_preio (
            .PADOEN(N__6372),
            .PADOUT(N__6371),
            .PADIN(N__6370),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5996),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_22_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_22_iopad (
            .OE(N__6363),
            .DIN(N__6362),
            .DOUT(N__6361),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__6363),
            .PADOUT(N__6362),
            .PADIN(N__6361),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_27_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_27_iopad (
            .OE(N__6354),
            .DIN(N__6353),
            .DOUT(N__6352),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__6354),
            .PADOUT(N__6353),
            .PADIN(N__6352),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__6345),
            .DIN(N__6344),
            .DOUT(N__6343),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__6345),
            .PADOUT(N__6344),
            .PADIN(N__6343),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__6336),
            .DIN(N__6335),
            .DOUT(N__6334),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__6336),
            .PADOUT(N__6335),
            .PADIN(N__6334),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_20_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_20_iopad (
            .OE(N__6327),
            .DIN(N__6326),
            .DOUT(N__6325),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__6327),
            .PADOUT(N__6326),
            .PADIN(N__6325),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_13_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_13_iopad (
            .OE(N__6318),
            .DIN(N__6317),
            .DOUT(N__6316),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__6318),
            .PADOUT(N__6317),
            .PADIN(N__6316),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_25_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_25_iopad (
            .OE(N__6309),
            .DIN(N__6308),
            .DOUT(N__6307),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__6309),
            .PADOUT(N__6308),
            .PADIN(N__6307),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nREGSPACE_obuf_iopad (
            .OE(N__6300),
            .DIN(N__6299),
            .DOUT(N__6298),
            .PACKAGEPIN(nREGSPACE));
    defparam nREGSPACE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nREGSPACE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nREGSPACE_obuf_preio (
            .PADOEN(N__6300),
            .PADOUT(N__6299),
            .PADIN(N__6298),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3611),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__6291),
            .DIN(N__6290),
            .DOUT(N__6289),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__6291),
            .PADOUT(N__6290),
            .PADIN(N__6289),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3572),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_19_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_19_iopad (
            .OE(N__6282),
            .DIN(N__6281),
            .DOUT(N__6280),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__6282),
            .PADOUT(N__6281),
            .PADIN(N__6280),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_28_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_28_iopad (
            .OE(N__6273),
            .DIN(N__6272),
            .DOUT(N__6271),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__6273),
            .PADOUT(N__6272),
            .PADIN(N__6271),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_30_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_30_iopad (
            .OE(N__6264),
            .DIN(N__6263),
            .DOUT(N__6262),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__6264),
            .PADOUT(N__6263),
            .PADIN(N__6262),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__6255),
            .DIN(N__6254),
            .DOUT(N__6253),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__6255),
            .PADOUT(N__6254),
            .PADIN(N__6253),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_16_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_16_iopad (
            .OE(N__6246),
            .DIN(N__6245),
            .DOUT(N__6244),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__6246),
            .PADOUT(N__6245),
            .PADIN(N__6244),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__6237),
            .DIN(N__6236),
            .DOUT(N__6235),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__6237),
            .PADOUT(N__6236),
            .PADIN(N__6235),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4595),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_26_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_26_iopad (
            .OE(N__6228),
            .DIN(N__6227),
            .DOUT(N__6226),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__6228),
            .PADOUT(N__6227),
            .PADIN(N__6226),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_23_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_23_iopad (
            .OE(N__6219),
            .DIN(N__6218),
            .DOUT(N__6217),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__6219),
            .PADOUT(N__6218),
            .PADIN(N__6217),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__1457 (
            .O(N__6200),
            .I(N__6195));
    InMux I__1456 (
            .O(N__6199),
            .I(N__6188));
    InMux I__1455 (
            .O(N__6198),
            .I(N__6188));
    InMux I__1454 (
            .O(N__6195),
            .I(N__6188));
    LocalMux I__1453 (
            .O(N__6188),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    InMux I__1452 (
            .O(N__6185),
            .I(N__6176));
    InMux I__1451 (
            .O(N__6184),
            .I(N__6176));
    InMux I__1450 (
            .O(N__6183),
            .I(N__6176));
    LocalMux I__1449 (
            .O(N__6176),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    InMux I__1448 (
            .O(N__6173),
            .I(N__6169));
    InMux I__1447 (
            .O(N__6172),
            .I(N__6166));
    LocalMux I__1446 (
            .O(N__6169),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ));
    LocalMux I__1445 (
            .O(N__6166),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ));
    CEMux I__1444 (
            .O(N__6161),
            .I(N__6158));
    LocalMux I__1443 (
            .O(N__6158),
            .I(N__6155));
    Odrv4 I__1442 (
            .O(N__6155),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ));
    InMux I__1441 (
            .O(N__6152),
            .I(N__6148));
    CascadeMux I__1440 (
            .O(N__6151),
            .I(N__6144));
    LocalMux I__1439 (
            .O(N__6148),
            .I(N__6141));
    InMux I__1438 (
            .O(N__6147),
            .I(N__6138));
    InMux I__1437 (
            .O(N__6144),
            .I(N__6135));
    Span4Mux_v I__1436 (
            .O(N__6141),
            .I(N__6132));
    LocalMux I__1435 (
            .O(N__6138),
            .I(N__6127));
    LocalMux I__1434 (
            .O(N__6135),
            .I(N__6127));
    Span4Mux_h I__1433 (
            .O(N__6132),
            .I(N__6120));
    Span4Mux_v I__1432 (
            .O(N__6127),
            .I(N__6120));
    CascadeMux I__1431 (
            .O(N__6126),
            .I(N__6117));
    CascadeMux I__1430 (
            .O(N__6125),
            .I(N__6113));
    Span4Mux_h I__1429 (
            .O(N__6120),
            .I(N__6103));
    InMux I__1428 (
            .O(N__6117),
            .I(N__6098));
    InMux I__1427 (
            .O(N__6116),
            .I(N__6098));
    InMux I__1426 (
            .O(N__6113),
            .I(N__6093));
    InMux I__1425 (
            .O(N__6112),
            .I(N__6093));
    InMux I__1424 (
            .O(N__6111),
            .I(N__6090));
    InMux I__1423 (
            .O(N__6110),
            .I(N__6086));
    InMux I__1422 (
            .O(N__6109),
            .I(N__6083));
    InMux I__1421 (
            .O(N__6108),
            .I(N__6080));
    InMux I__1420 (
            .O(N__6107),
            .I(N__6075));
    InMux I__1419 (
            .O(N__6106),
            .I(N__6075));
    Span4Mux_h I__1418 (
            .O(N__6103),
            .I(N__6070));
    LocalMux I__1417 (
            .O(N__6098),
            .I(N__6070));
    LocalMux I__1416 (
            .O(N__6093),
            .I(N__6067));
    LocalMux I__1415 (
            .O(N__6090),
            .I(N__6064));
    InMux I__1414 (
            .O(N__6089),
            .I(N__6061));
    LocalMux I__1413 (
            .O(N__6086),
            .I(N__6058));
    LocalMux I__1412 (
            .O(N__6083),
            .I(N__6055));
    LocalMux I__1411 (
            .O(N__6080),
            .I(N__6050));
    LocalMux I__1410 (
            .O(N__6075),
            .I(N__6050));
    Span4Mux_v I__1409 (
            .O(N__6070),
            .I(N__6041));
    Span4Mux_v I__1408 (
            .O(N__6067),
            .I(N__6041));
    Span4Mux_h I__1407 (
            .O(N__6064),
            .I(N__6041));
    LocalMux I__1406 (
            .O(N__6061),
            .I(N__6041));
    Span4Mux_v I__1405 (
            .O(N__6058),
            .I(N__6038));
    Sp12to4 I__1404 (
            .O(N__6055),
            .I(N__6035));
    Span4Mux_v I__1403 (
            .O(N__6050),
            .I(N__6032));
    Span4Mux_v I__1402 (
            .O(N__6041),
            .I(N__6029));
    Sp12to4 I__1401 (
            .O(N__6038),
            .I(N__6026));
    Span12Mux_v I__1400 (
            .O(N__6035),
            .I(N__6021));
    Sp12to4 I__1399 (
            .O(N__6032),
            .I(N__6021));
    Sp12to4 I__1398 (
            .O(N__6029),
            .I(N__6018));
    Span12Mux_h I__1397 (
            .O(N__6026),
            .I(N__6015));
    Span12Mux_v I__1396 (
            .O(N__6021),
            .I(N__6012));
    Span12Mux_h I__1395 (
            .O(N__6018),
            .I(N__6009));
    Span12Mux_v I__1394 (
            .O(N__6015),
            .I(N__6006));
    Span12Mux_h I__1393 (
            .O(N__6012),
            .I(N__6001));
    Span12Mux_v I__1392 (
            .O(N__6009),
            .I(N__6001));
    Odrv12 I__1391 (
            .O(N__6006),
            .I(RESETn_c));
    Odrv12 I__1390 (
            .O(N__6001),
            .I(RESETn_c));
    IoInMux I__1389 (
            .O(N__5996),
            .I(N__5993));
    LocalMux I__1388 (
            .O(N__5993),
            .I(N__5990));
    Span4Mux_s3_v I__1387 (
            .O(N__5990),
            .I(N__5987));
    Sp12to4 I__1386 (
            .O(N__5987),
            .I(N__5984));
    Span12Mux_h I__1385 (
            .O(N__5984),
            .I(N__5980));
    InMux I__1384 (
            .O(N__5983),
            .I(N__5977));
    Span12Mux_v I__1383 (
            .O(N__5980),
            .I(N__5972));
    LocalMux I__1382 (
            .O(N__5977),
            .I(N__5972));
    Odrv12 I__1381 (
            .O(N__5972),
            .I(nBUFEN_c));
    InMux I__1380 (
            .O(N__5969),
            .I(N__5966));
    LocalMux I__1379 (
            .O(N__5966),
            .I(N__5963));
    Span4Mux_v I__1378 (
            .O(N__5963),
            .I(N__5960));
    Sp12to4 I__1377 (
            .O(N__5960),
            .I(N__5957));
    Span12Mux_h I__1376 (
            .O(N__5957),
            .I(N__5954));
    Span12Mux_v I__1375 (
            .O(N__5954),
            .I(N__5951));
    Odrv12 I__1374 (
            .O(N__5951),
            .I(TACKn_in));
    SRMux I__1373 (
            .O(N__5948),
            .I(N__5944));
    SRMux I__1372 (
            .O(N__5947),
            .I(N__5940));
    LocalMux I__1371 (
            .O(N__5944),
            .I(N__5937));
    SRMux I__1370 (
            .O(N__5943),
            .I(N__5933));
    LocalMux I__1369 (
            .O(N__5940),
            .I(N__5930));
    Span4Mux_v I__1368 (
            .O(N__5937),
            .I(N__5927));
    SRMux I__1367 (
            .O(N__5936),
            .I(N__5924));
    LocalMux I__1366 (
            .O(N__5933),
            .I(N__5921));
    Span4Mux_v I__1365 (
            .O(N__5930),
            .I(N__5914));
    Span4Mux_v I__1364 (
            .O(N__5927),
            .I(N__5914));
    LocalMux I__1363 (
            .O(N__5924),
            .I(N__5914));
    Span4Mux_v I__1362 (
            .O(N__5921),
            .I(N__5911));
    Span4Mux_h I__1361 (
            .O(N__5914),
            .I(N__5908));
    Span4Mux_h I__1360 (
            .O(N__5911),
            .I(N__5903));
    Span4Mux_h I__1359 (
            .O(N__5908),
            .I(N__5903));
    Odrv4 I__1358 (
            .O(N__5903),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__1357 (
            .O(N__5900),
            .I(N__5897));
    LocalMux I__1356 (
            .O(N__5897),
            .I(N__5894));
    Span4Mux_v I__1355 (
            .O(N__5894),
            .I(N__5891));
    Span4Mux_h I__1354 (
            .O(N__5891),
            .I(N__5888));
    Odrv4 I__1353 (
            .O(N__5888),
            .I(TACK_EN_i));
    IoInMux I__1352 (
            .O(N__5885),
            .I(N__5882));
    LocalMux I__1351 (
            .O(N__5882),
            .I(N__5879));
    Span4Mux_s2_v I__1350 (
            .O(N__5879),
            .I(N__5876));
    Span4Mux_h I__1349 (
            .O(N__5876),
            .I(N__5873));
    Span4Mux_v I__1348 (
            .O(N__5873),
            .I(N__5870));
    Odrv4 I__1347 (
            .O(N__5870),
            .I(N_365_i));
    InMux I__1346 (
            .O(N__5867),
            .I(N__5856));
    InMux I__1345 (
            .O(N__5866),
            .I(N__5856));
    InMux I__1344 (
            .O(N__5865),
            .I(N__5849));
    InMux I__1343 (
            .O(N__5864),
            .I(N__5849));
    InMux I__1342 (
            .O(N__5863),
            .I(N__5849));
    InMux I__1341 (
            .O(N__5862),
            .I(N__5844));
    InMux I__1340 (
            .O(N__5861),
            .I(N__5844));
    LocalMux I__1339 (
            .O(N__5856),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1338 (
            .O(N__5849),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1337 (
            .O(N__5844),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    InMux I__1336 (
            .O(N__5837),
            .I(N__5834));
    LocalMux I__1335 (
            .O(N__5834),
            .I(\U409_CIA.CLKCIA6_0_a2_1 ));
    CascadeMux I__1334 (
            .O(N__5831),
            .I(N__5826));
    CascadeMux I__1333 (
            .O(N__5830),
            .I(N__5823));
    InMux I__1332 (
            .O(N__5829),
            .I(N__5819));
    InMux I__1331 (
            .O(N__5826),
            .I(N__5814));
    InMux I__1330 (
            .O(N__5823),
            .I(N__5814));
    InMux I__1329 (
            .O(N__5822),
            .I(N__5811));
    LocalMux I__1328 (
            .O(N__5819),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1327 (
            .O(N__5814),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1326 (
            .O(N__5811),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    InMux I__1325 (
            .O(N__5804),
            .I(N__5798));
    InMux I__1324 (
            .O(N__5803),
            .I(N__5795));
    InMux I__1323 (
            .O(N__5802),
            .I(N__5790));
    InMux I__1322 (
            .O(N__5801),
            .I(N__5790));
    LocalMux I__1321 (
            .O(N__5798),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1320 (
            .O(N__5795),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1319 (
            .O(N__5790),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    InMux I__1318 (
            .O(N__5783),
            .I(N__5775));
    InMux I__1317 (
            .O(N__5782),
            .I(N__5775));
    InMux I__1316 (
            .O(N__5781),
            .I(N__5772));
    InMux I__1315 (
            .O(N__5780),
            .I(N__5769));
    LocalMux I__1314 (
            .O(N__5775),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1313 (
            .O(N__5772),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1312 (
            .O(N__5769),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    InMux I__1311 (
            .O(N__5762),
            .I(N__5758));
    InMux I__1310 (
            .O(N__5761),
            .I(N__5755));
    LocalMux I__1309 (
            .O(N__5758),
            .I(\U409_CIA.CLKCIA8_0_a2_0 ));
    LocalMux I__1308 (
            .O(N__5755),
            .I(\U409_CIA.CLKCIA8_0_a2_0 ));
    SRMux I__1307 (
            .O(N__5750),
            .I(N__5746));
    SRMux I__1306 (
            .O(N__5749),
            .I(N__5743));
    LocalMux I__1305 (
            .O(N__5746),
            .I(N__5737));
    LocalMux I__1304 (
            .O(N__5743),
            .I(N__5737));
    SRMux I__1303 (
            .O(N__5742),
            .I(N__5734));
    Span4Mux_v I__1302 (
            .O(N__5737),
            .I(N__5731));
    LocalMux I__1301 (
            .O(N__5734),
            .I(N__5728));
    Odrv4 I__1300 (
            .O(N__5731),
            .I(RESETn_c_i));
    Odrv4 I__1299 (
            .O(N__5728),
            .I(RESETn_c_i));
    InMux I__1298 (
            .O(N__5723),
            .I(N__5720));
    LocalMux I__1297 (
            .O(N__5720),
            .I(N__5717));
    Span4Mux_v I__1296 (
            .O(N__5717),
            .I(N__5714));
    Odrv4 I__1295 (
            .O(N__5714),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ));
    InMux I__1294 (
            .O(N__5711),
            .I(N__5707));
    InMux I__1293 (
            .O(N__5710),
            .I(N__5704));
    LocalMux I__1292 (
            .O(N__5707),
            .I(N__5701));
    LocalMux I__1291 (
            .O(N__5704),
            .I(N__5698));
    Span4Mux_v I__1290 (
            .O(N__5701),
            .I(N__5695));
    Span4Mux_v I__1289 (
            .O(N__5698),
            .I(N__5692));
    Odrv4 I__1288 (
            .O(N__5695),
            .I(\U409_ADDRESS_DECODE.un5_nRAMSPACEZ0 ));
    Odrv4 I__1287 (
            .O(N__5692),
            .I(\U409_ADDRESS_DECODE.un5_nRAMSPACEZ0 ));
    CascadeMux I__1286 (
            .O(N__5687),
            .I(N__5684));
    InMux I__1285 (
            .O(N__5684),
            .I(N__5680));
    InMux I__1284 (
            .O(N__5683),
            .I(N__5677));
    LocalMux I__1283 (
            .O(N__5680),
            .I(N__5668));
    LocalMux I__1282 (
            .O(N__5677),
            .I(N__5668));
    InMux I__1281 (
            .O(N__5676),
            .I(N__5665));
    InMux I__1280 (
            .O(N__5675),
            .I(N__5662));
    InMux I__1279 (
            .O(N__5674),
            .I(N__5659));
    InMux I__1278 (
            .O(N__5673),
            .I(N__5655));
    Span4Mux_h I__1277 (
            .O(N__5668),
            .I(N__5648));
    LocalMux I__1276 (
            .O(N__5665),
            .I(N__5648));
    LocalMux I__1275 (
            .O(N__5662),
            .I(N__5648));
    LocalMux I__1274 (
            .O(N__5659),
            .I(N__5645));
    CascadeMux I__1273 (
            .O(N__5658),
            .I(N__5641));
    LocalMux I__1272 (
            .O(N__5655),
            .I(N__5638));
    Span4Mux_v I__1271 (
            .O(N__5648),
            .I(N__5633));
    Span4Mux_v I__1270 (
            .O(N__5645),
            .I(N__5633));
    InMux I__1269 (
            .O(N__5644),
            .I(N__5630));
    InMux I__1268 (
            .O(N__5641),
            .I(N__5627));
    Span12Mux_h I__1267 (
            .O(N__5638),
            .I(N__5624));
    Sp12to4 I__1266 (
            .O(N__5633),
            .I(N__5621));
    LocalMux I__1265 (
            .O(N__5630),
            .I(N__5616));
    LocalMux I__1264 (
            .O(N__5627),
            .I(N__5616));
    Span12Mux_v I__1263 (
            .O(N__5624),
            .I(N__5613));
    Span12Mux_h I__1262 (
            .O(N__5621),
            .I(N__5610));
    Span4Mux_v I__1261 (
            .O(N__5616),
            .I(N__5607));
    Odrv12 I__1260 (
            .O(N__5613),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ));
    Odrv12 I__1259 (
            .O(N__5610),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ));
    Odrv4 I__1258 (
            .O(N__5607),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ));
    CascadeMux I__1257 (
            .O(N__5600),
            .I(N__5597));
    InMux I__1256 (
            .O(N__5597),
            .I(N__5594));
    LocalMux I__1255 (
            .O(N__5594),
            .I(N__5590));
    InMux I__1254 (
            .O(N__5593),
            .I(N__5586));
    Span4Mux_v I__1253 (
            .O(N__5590),
            .I(N__5583));
    InMux I__1252 (
            .O(N__5589),
            .I(N__5580));
    LocalMux I__1251 (
            .O(N__5586),
            .I(N__5577));
    Span4Mux_v I__1250 (
            .O(N__5583),
            .I(N__5574));
    LocalMux I__1249 (
            .O(N__5580),
            .I(N__5571));
    Span12Mux_h I__1248 (
            .O(N__5577),
            .I(N__5568));
    Sp12to4 I__1247 (
            .O(N__5574),
            .I(N__5563));
    Span12Mux_v I__1246 (
            .O(N__5571),
            .I(N__5563));
    Span12Mux_v I__1245 (
            .O(N__5568),
            .I(N__5558));
    Span12Mux_h I__1244 (
            .O(N__5563),
            .I(N__5558));
    Odrv12 I__1243 (
            .O(N__5558),
            .I(OVL_c));
    IoInMux I__1242 (
            .O(N__5555),
            .I(N__5552));
    LocalMux I__1241 (
            .O(N__5552),
            .I(N__5549));
    Span4Mux_s3_v I__1240 (
            .O(N__5549),
            .I(N__5546));
    Span4Mux_h I__1239 (
            .O(N__5546),
            .I(N__5543));
    Sp12to4 I__1238 (
            .O(N__5543),
            .I(N__5540));
    Span12Mux_v I__1237 (
            .O(N__5540),
            .I(N__5536));
    InMux I__1236 (
            .O(N__5539),
            .I(N__5533));
    Odrv12 I__1235 (
            .O(N__5536),
            .I(TACK_OUTn));
    LocalMux I__1234 (
            .O(N__5533),
            .I(TACK_OUTn));
    InMux I__1233 (
            .O(N__5528),
            .I(N__5524));
    InMux I__1232 (
            .O(N__5527),
            .I(N__5521));
    LocalMux I__1231 (
            .O(N__5524),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__1230 (
            .O(N__5521),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__1229 (
            .O(N__5516),
            .I(N__5513));
    LocalMux I__1228 (
            .O(N__5513),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER5_0 ));
    CascadeMux I__1227 (
            .O(N__5510),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ));
    InMux I__1226 (
            .O(N__5507),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    CascadeMux I__1225 (
            .O(N__5504),
            .I(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ));
    InMux I__1224 (
            .O(N__5501),
            .I(N__5498));
    LocalMux I__1223 (
            .O(N__5498),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ));
    InMux I__1222 (
            .O(N__5495),
            .I(N__5492));
    LocalMux I__1221 (
            .O(N__5492),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ));
    CascadeMux I__1220 (
            .O(N__5489),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_ ));
    CascadeMux I__1219 (
            .O(N__5486),
            .I(\U409_CIA.N_20_cascade_ ));
    CascadeMux I__1218 (
            .O(N__5483),
            .I(N__5473));
    InMux I__1217 (
            .O(N__5482),
            .I(N__5470));
    InMux I__1216 (
            .O(N__5481),
            .I(N__5463));
    InMux I__1215 (
            .O(N__5480),
            .I(N__5463));
    InMux I__1214 (
            .O(N__5479),
            .I(N__5463));
    InMux I__1213 (
            .O(N__5478),
            .I(N__5454));
    InMux I__1212 (
            .O(N__5477),
            .I(N__5454));
    InMux I__1211 (
            .O(N__5476),
            .I(N__5454));
    InMux I__1210 (
            .O(N__5473),
            .I(N__5454));
    LocalMux I__1209 (
            .O(N__5470),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1208 (
            .O(N__5463),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1207 (
            .O(N__5454),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    CascadeMux I__1206 (
            .O(N__5447),
            .I(\U409_CIA.CLKCIAZ0_cascade_ ));
    InMux I__1205 (
            .O(N__5444),
            .I(N__5436));
    InMux I__1204 (
            .O(N__5443),
            .I(N__5429));
    InMux I__1203 (
            .O(N__5442),
            .I(N__5429));
    InMux I__1202 (
            .O(N__5441),
            .I(N__5429));
    InMux I__1201 (
            .O(N__5440),
            .I(N__5424));
    InMux I__1200 (
            .O(N__5439),
            .I(N__5424));
    LocalMux I__1199 (
            .O(N__5436),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1198 (
            .O(N__5429),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1197 (
            .O(N__5424),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    IoInMux I__1196 (
            .O(N__5417),
            .I(N__5414));
    LocalMux I__1195 (
            .O(N__5414),
            .I(N__5411));
    Span12Mux_s6_v I__1194 (
            .O(N__5411),
            .I(N__5407));
    InMux I__1193 (
            .O(N__5410),
            .I(N__5404));
    Span12Mux_v I__1192 (
            .O(N__5407),
            .I(N__5400));
    LocalMux I__1191 (
            .O(N__5404),
            .I(N__5397));
    InMux I__1190 (
            .O(N__5403),
            .I(N__5394));
    Odrv12 I__1189 (
            .O(N__5400),
            .I(CLKCIA_c));
    Odrv4 I__1188 (
            .O(N__5397),
            .I(CLKCIA_c));
    LocalMux I__1187 (
            .O(N__5394),
            .I(CLKCIA_c));
    ClkMux I__1186 (
            .O(N__5387),
            .I(N__5375));
    ClkMux I__1185 (
            .O(N__5386),
            .I(N__5375));
    ClkMux I__1184 (
            .O(N__5385),
            .I(N__5375));
    ClkMux I__1183 (
            .O(N__5384),
            .I(N__5375));
    GlobalMux I__1182 (
            .O(N__5375),
            .I(N__5372));
    gio2CtrlBuf I__1181 (
            .O(N__5372),
            .I(CLK28_IN_c_g));
    CascadeMux I__1180 (
            .O(N__5369),
            .I(N__5365));
    CascadeMux I__1179 (
            .O(N__5368),
            .I(N__5362));
    InMux I__1178 (
            .O(N__5365),
            .I(N__5357));
    InMux I__1177 (
            .O(N__5362),
            .I(N__5357));
    LocalMux I__1176 (
            .O(N__5357),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ));
    InMux I__1175 (
            .O(N__5354),
            .I(N__5351));
    LocalMux I__1174 (
            .O(N__5351),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ));
    InMux I__1173 (
            .O(N__5348),
            .I(N__5337));
    InMux I__1172 (
            .O(N__5347),
            .I(N__5337));
    InMux I__1171 (
            .O(N__5346),
            .I(N__5337));
    InMux I__1170 (
            .O(N__5345),
            .I(N__5332));
    InMux I__1169 (
            .O(N__5344),
            .I(N__5332));
    LocalMux I__1168 (
            .O(N__5337),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1167 (
            .O(N__5332),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    InMux I__1166 (
            .O(N__5327),
            .I(N__5316));
    InMux I__1165 (
            .O(N__5326),
            .I(N__5316));
    InMux I__1164 (
            .O(N__5325),
            .I(N__5316));
    InMux I__1163 (
            .O(N__5324),
            .I(N__5311));
    InMux I__1162 (
            .O(N__5323),
            .I(N__5311));
    LocalMux I__1161 (
            .O(N__5316),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1160 (
            .O(N__5311),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    CascadeMux I__1159 (
            .O(N__5306),
            .I(N__5301));
    CascadeMux I__1158 (
            .O(N__5305),
            .I(N__5297));
    InMux I__1157 (
            .O(N__5304),
            .I(N__5289));
    InMux I__1156 (
            .O(N__5301),
            .I(N__5289));
    InMux I__1155 (
            .O(N__5300),
            .I(N__5289));
    InMux I__1154 (
            .O(N__5297),
            .I(N__5284));
    InMux I__1153 (
            .O(N__5296),
            .I(N__5284));
    LocalMux I__1152 (
            .O(N__5289),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1151 (
            .O(N__5284),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__1150 (
            .O(N__5279),
            .I(N__5276));
    LocalMux I__1149 (
            .O(N__5276),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0 ));
    InMux I__1148 (
            .O(N__5273),
            .I(N__5270));
    LocalMux I__1147 (
            .O(N__5270),
            .I(N__5261));
    InMux I__1146 (
            .O(N__5269),
            .I(N__5256));
    InMux I__1145 (
            .O(N__5268),
            .I(N__5256));
    InMux I__1144 (
            .O(N__5267),
            .I(N__5253));
    InMux I__1143 (
            .O(N__5266),
            .I(N__5246));
    InMux I__1142 (
            .O(N__5265),
            .I(N__5246));
    InMux I__1141 (
            .O(N__5264),
            .I(N__5246));
    Odrv4 I__1140 (
            .O(N__5261),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__1139 (
            .O(N__5256),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__1138 (
            .O(N__5253),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__1137 (
            .O(N__5246),
            .I(\U409_TICK.TICK603_14 ));
    InMux I__1136 (
            .O(N__5237),
            .I(N__5228));
    InMux I__1135 (
            .O(N__5236),
            .I(N__5225));
    InMux I__1134 (
            .O(N__5235),
            .I(N__5218));
    InMux I__1133 (
            .O(N__5234),
            .I(N__5218));
    InMux I__1132 (
            .O(N__5233),
            .I(N__5218));
    InMux I__1131 (
            .O(N__5232),
            .I(N__5213));
    InMux I__1130 (
            .O(N__5231),
            .I(N__5213));
    LocalMux I__1129 (
            .O(N__5228),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__1128 (
            .O(N__5225),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__1127 (
            .O(N__5218),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__1126 (
            .O(N__5213),
            .I(\U409_TICK.TICK603_10 ));
    CascadeMux I__1125 (
            .O(N__5204),
            .I(N__5199));
    CascadeMux I__1124 (
            .O(N__5203),
            .I(N__5196));
    CascadeMux I__1123 (
            .O(N__5202),
            .I(N__5189));
    InMux I__1122 (
            .O(N__5199),
            .I(N__5186));
    InMux I__1121 (
            .O(N__5196),
            .I(N__5183));
    InMux I__1120 (
            .O(N__5195),
            .I(N__5180));
    InMux I__1119 (
            .O(N__5194),
            .I(N__5175));
    InMux I__1118 (
            .O(N__5193),
            .I(N__5175));
    InMux I__1117 (
            .O(N__5192),
            .I(N__5170));
    InMux I__1116 (
            .O(N__5189),
            .I(N__5170));
    LocalMux I__1115 (
            .O(N__5186),
            .I(N__5167));
    LocalMux I__1114 (
            .O(N__5183),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__1113 (
            .O(N__5180),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__1112 (
            .O(N__5175),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__1111 (
            .O(N__5170),
            .I(\U409_TICK.TICK603_9 ));
    Odrv4 I__1110 (
            .O(N__5167),
            .I(\U409_TICK.TICK603_9 ));
    InMux I__1109 (
            .O(N__5156),
            .I(N__5153));
    LocalMux I__1108 (
            .O(N__5153),
            .I(N__5150));
    Odrv4 I__1107 (
            .O(N__5150),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__1106 (
            .O(N__5147),
            .I(N__5143));
    InMux I__1105 (
            .O(N__5146),
            .I(N__5140));
    LocalMux I__1104 (
            .O(N__5143),
            .I(N__5137));
    LocalMux I__1103 (
            .O(N__5140),
            .I(N__5134));
    Odrv4 I__1102 (
            .O(N__5137),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    Odrv4 I__1101 (
            .O(N__5134),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    ClkMux I__1100 (
            .O(N__5129),
            .I(N__5093));
    ClkMux I__1099 (
            .O(N__5128),
            .I(N__5093));
    ClkMux I__1098 (
            .O(N__5127),
            .I(N__5093));
    ClkMux I__1097 (
            .O(N__5126),
            .I(N__5093));
    ClkMux I__1096 (
            .O(N__5125),
            .I(N__5093));
    ClkMux I__1095 (
            .O(N__5124),
            .I(N__5093));
    ClkMux I__1094 (
            .O(N__5123),
            .I(N__5093));
    ClkMux I__1093 (
            .O(N__5122),
            .I(N__5093));
    ClkMux I__1092 (
            .O(N__5121),
            .I(N__5093));
    ClkMux I__1091 (
            .O(N__5120),
            .I(N__5093));
    ClkMux I__1090 (
            .O(N__5119),
            .I(N__5093));
    ClkMux I__1089 (
            .O(N__5118),
            .I(N__5093));
    GlobalMux I__1088 (
            .O(N__5093),
            .I(N__5090));
    gio2CtrlBuf I__1087 (
            .O(N__5090),
            .I(CLK6_c_g));
    InMux I__1086 (
            .O(N__5087),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__1085 (
            .O(N__5084),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__1084 (
            .O(N__5081),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__1083 (
            .O(N__5078),
            .I(N__5075));
    LocalMux I__1082 (
            .O(N__5075),
            .I(N__5072));
    Span4Mux_v I__1081 (
            .O(N__5072),
            .I(N__5067));
    InMux I__1080 (
            .O(N__5071),
            .I(N__5062));
    InMux I__1079 (
            .O(N__5070),
            .I(N__5062));
    Sp12to4 I__1078 (
            .O(N__5067),
            .I(N__5057));
    LocalMux I__1077 (
            .O(N__5062),
            .I(N__5057));
    Odrv12 I__1076 (
            .O(N__5057),
            .I(\U409_CIA.g0Z0Z_14 ));
    CascadeMux I__1075 (
            .O(N__5054),
            .I(N__5050));
    InMux I__1074 (
            .O(N__5053),
            .I(N__5045));
    InMux I__1073 (
            .O(N__5050),
            .I(N__5040));
    InMux I__1072 (
            .O(N__5049),
            .I(N__5040));
    InMux I__1071 (
            .O(N__5048),
            .I(N__5037));
    LocalMux I__1070 (
            .O(N__5045),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__1069 (
            .O(N__5040),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__1068 (
            .O(N__5037),
            .I(\U409_CIA.VMAZ0 ));
    CascadeMux I__1067 (
            .O(N__5030),
            .I(N__5026));
    InMux I__1066 (
            .O(N__5029),
            .I(N__5020));
    InMux I__1065 (
            .O(N__5026),
            .I(N__5020));
    CascadeMux I__1064 (
            .O(N__5025),
            .I(N__5017));
    LocalMux I__1063 (
            .O(N__5020),
            .I(N__5014));
    InMux I__1062 (
            .O(N__5017),
            .I(N__5011));
    Span4Mux_v I__1061 (
            .O(N__5014),
            .I(N__5006));
    LocalMux I__1060 (
            .O(N__5011),
            .I(N__5006));
    Span4Mux_v I__1059 (
            .O(N__5006),
            .I(N__5003));
    Sp12to4 I__1058 (
            .O(N__5003),
            .I(N__5000));
    Span12Mux_h I__1057 (
            .O(N__5000),
            .I(N__4997));
    Odrv12 I__1056 (
            .O(N__4997),
            .I(\U409_CIA.g0Z0Z_13 ));
    InMux I__1055 (
            .O(N__4994),
            .I(N__4991));
    LocalMux I__1054 (
            .O(N__4991),
            .I(N__4986));
    InMux I__1053 (
            .O(N__4990),
            .I(N__4981));
    InMux I__1052 (
            .O(N__4989),
            .I(N__4981));
    Odrv4 I__1051 (
            .O(N__4986),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    LocalMux I__1050 (
            .O(N__4981),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    CascadeMux I__1049 (
            .O(N__4976),
            .I(N__4970));
    InMux I__1048 (
            .O(N__4975),
            .I(N__4967));
    InMux I__1047 (
            .O(N__4974),
            .I(N__4960));
    InMux I__1046 (
            .O(N__4973),
            .I(N__4960));
    InMux I__1045 (
            .O(N__4970),
            .I(N__4960));
    LocalMux I__1044 (
            .O(N__4967),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1043 (
            .O(N__4960),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    InMux I__1042 (
            .O(N__4955),
            .I(N__4948));
    InMux I__1041 (
            .O(N__4954),
            .I(N__4939));
    InMux I__1040 (
            .O(N__4953),
            .I(N__4939));
    InMux I__1039 (
            .O(N__4952),
            .I(N__4939));
    InMux I__1038 (
            .O(N__4951),
            .I(N__4939));
    LocalMux I__1037 (
            .O(N__4948),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__1036 (
            .O(N__4939),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    CascadeMux I__1035 (
            .O(N__4934),
            .I(N__4931));
    InMux I__1034 (
            .O(N__4931),
            .I(N__4928));
    LocalMux I__1033 (
            .O(N__4928),
            .I(\U409_TRANSFER_ACK.N_105 ));
    InMux I__1032 (
            .O(N__4925),
            .I(N__4919));
    InMux I__1031 (
            .O(N__4924),
            .I(N__4912));
    InMux I__1030 (
            .O(N__4923),
            .I(N__4912));
    InMux I__1029 (
            .O(N__4922),
            .I(N__4912));
    LocalMux I__1028 (
            .O(N__4919),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__1027 (
            .O(N__4912),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    CascadeMux I__1026 (
            .O(N__4907),
            .I(N__4904));
    InMux I__1025 (
            .O(N__4904),
            .I(N__4895));
    InMux I__1024 (
            .O(N__4903),
            .I(N__4895));
    InMux I__1023 (
            .O(N__4902),
            .I(N__4895));
    LocalMux I__1022 (
            .O(N__4895),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    InMux I__1021 (
            .O(N__4892),
            .I(N__4887));
    InMux I__1020 (
            .O(N__4891),
            .I(N__4882));
    InMux I__1019 (
            .O(N__4890),
            .I(N__4882));
    LocalMux I__1018 (
            .O(N__4887),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__1017 (
            .O(N__4882),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__1016 (
            .O(N__4877),
            .I(N__4871));
    InMux I__1015 (
            .O(N__4876),
            .I(N__4871));
    LocalMux I__1014 (
            .O(N__4871),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    InMux I__1013 (
            .O(N__4868),
            .I(N__4864));
    InMux I__1012 (
            .O(N__4867),
            .I(N__4861));
    LocalMux I__1011 (
            .O(N__4864),
            .I(N__4858));
    LocalMux I__1010 (
            .O(N__4861),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    Odrv4 I__1009 (
            .O(N__4858),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    InMux I__1008 (
            .O(N__4853),
            .I(N__4849));
    InMux I__1007 (
            .O(N__4852),
            .I(N__4846));
    LocalMux I__1006 (
            .O(N__4849),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__1005 (
            .O(N__4846),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    InMux I__1004 (
            .O(N__4841),
            .I(N__4837));
    InMux I__1003 (
            .O(N__4840),
            .I(N__4834));
    LocalMux I__1002 (
            .O(N__4837),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__1001 (
            .O(N__4834),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__1000 (
            .O(N__4829),
            .I(N__4825));
    InMux I__999 (
            .O(N__4828),
            .I(N__4822));
    LocalMux I__998 (
            .O(N__4825),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__997 (
            .O(N__4822),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    CascadeMux I__996 (
            .O(N__4817),
            .I(N__4814));
    InMux I__995 (
            .O(N__4814),
            .I(N__4811));
    LocalMux I__994 (
            .O(N__4811),
            .I(N__4807));
    InMux I__993 (
            .O(N__4810),
            .I(N__4804));
    Odrv4 I__992 (
            .O(N__4807),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__991 (
            .O(N__4804),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    CascadeMux I__990 (
            .O(N__4799),
            .I(N__4795));
    InMux I__989 (
            .O(N__4798),
            .I(N__4792));
    InMux I__988 (
            .O(N__4795),
            .I(N__4789));
    LocalMux I__987 (
            .O(N__4792),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__986 (
            .O(N__4789),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    CascadeMux I__985 (
            .O(N__4784),
            .I(\U409_TICK.TICK603_10_cascade_ ));
    InMux I__984 (
            .O(N__4781),
            .I(N__4778));
    LocalMux I__983 (
            .O(N__4778),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__982 (
            .O(N__4775),
            .I(N__4771));
    InMux I__981 (
            .O(N__4774),
            .I(N__4768));
    LocalMux I__980 (
            .O(N__4771),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__979 (
            .O(N__4768),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    InMux I__978 (
            .O(N__4763),
            .I(N__4759));
    InMux I__977 (
            .O(N__4762),
            .I(N__4756));
    LocalMux I__976 (
            .O(N__4759),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__975 (
            .O(N__4756),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__974 (
            .O(N__4751),
            .I(N__4747));
    InMux I__973 (
            .O(N__4750),
            .I(N__4744));
    LocalMux I__972 (
            .O(N__4747),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__971 (
            .O(N__4744),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    CascadeMux I__970 (
            .O(N__4739),
            .I(N__4733));
    InMux I__969 (
            .O(N__4738),
            .I(N__4730));
    InMux I__968 (
            .O(N__4737),
            .I(N__4725));
    InMux I__967 (
            .O(N__4736),
            .I(N__4725));
    InMux I__966 (
            .O(N__4733),
            .I(N__4722));
    LocalMux I__965 (
            .O(N__4730),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__964 (
            .O(N__4725),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__963 (
            .O(N__4722),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__962 (
            .O(N__4715),
            .I(N__4712));
    LocalMux I__961 (
            .O(N__4712),
            .I(\U409_TICK.TICK603_11 ));
    InMux I__960 (
            .O(N__4709),
            .I(N__4705));
    InMux I__959 (
            .O(N__4708),
            .I(N__4702));
    LocalMux I__958 (
            .O(N__4705),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__957 (
            .O(N__4702),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    CascadeMux I__956 (
            .O(N__4697),
            .I(\U409_TICK.TICK603_8_cascade_ ));
    InMux I__955 (
            .O(N__4694),
            .I(N__4690));
    InMux I__954 (
            .O(N__4693),
            .I(N__4687));
    LocalMux I__953 (
            .O(N__4690),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__952 (
            .O(N__4687),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    CascadeMux I__951 (
            .O(N__4682),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    InMux I__950 (
            .O(N__4679),
            .I(N__4676));
    LocalMux I__949 (
            .O(N__4676),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__948 (
            .O(N__4673),
            .I(N__4669));
    InMux I__947 (
            .O(N__4672),
            .I(N__4666));
    LocalMux I__946 (
            .O(N__4669),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__945 (
            .O(N__4666),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    InMux I__944 (
            .O(N__4661),
            .I(N__4655));
    InMux I__943 (
            .O(N__4660),
            .I(N__4655));
    LocalMux I__942 (
            .O(N__4655),
            .I(N__4652));
    Odrv4 I__941 (
            .O(N__4652),
            .I(CIA_ENABLEm));
    CascadeMux I__940 (
            .O(N__4649),
            .I(\U409_CIA.N_9_cascade_ ));
    InMux I__939 (
            .O(N__4646),
            .I(N__4643));
    LocalMux I__938 (
            .O(N__4643),
            .I(N__4640));
    Span4Mux_v I__937 (
            .O(N__4640),
            .I(N__4637));
    Sp12to4 I__936 (
            .O(N__4637),
            .I(N__4634));
    Span12Mux_h I__935 (
            .O(N__4634),
            .I(N__4631));
    Odrv12 I__934 (
            .O(N__4631),
            .I(A_c_13));
    IoInMux I__933 (
            .O(N__4628),
            .I(N__4625));
    LocalMux I__932 (
            .O(N__4625),
            .I(N__4622));
    Span12Mux_s4_h I__931 (
            .O(N__4622),
            .I(N__4619));
    Span12Mux_h I__930 (
            .O(N__4619),
            .I(N__4616));
    Odrv12 I__929 (
            .O(N__4616),
            .I(U409_ADDRESS_DECODE_un1_nCIACS1_i));
    IoInMux I__928 (
            .O(N__4613),
            .I(N__4610));
    LocalMux I__927 (
            .O(N__4610),
            .I(N__4607));
    Span12Mux_s4_v I__926 (
            .O(N__4607),
            .I(N__4604));
    Odrv12 I__925 (
            .O(N__4604),
            .I(U409_ADDRESS_DECODE_un1_nRAMSPACE_i));
    InMux I__924 (
            .O(N__4601),
            .I(N__4598));
    LocalMux I__923 (
            .O(N__4598),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    IoInMux I__922 (
            .O(N__4595),
            .I(N__4592));
    LocalMux I__921 (
            .O(N__4592),
            .I(N__4589));
    Span4Mux_s3_v I__920 (
            .O(N__4589),
            .I(N__4586));
    Sp12to4 I__919 (
            .O(N__4586),
            .I(N__4583));
    Span12Mux_h I__918 (
            .O(N__4583),
            .I(N__4579));
    InMux I__917 (
            .O(N__4582),
            .I(N__4576));
    Odrv12 I__916 (
            .O(N__4579),
            .I(TICK60_c));
    LocalMux I__915 (
            .O(N__4576),
            .I(TICK60_c));
    InMux I__914 (
            .O(N__4571),
            .I(N__4567));
    InMux I__913 (
            .O(N__4570),
            .I(N__4564));
    LocalMux I__912 (
            .O(N__4567),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__911 (
            .O(N__4564),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__910 (
            .O(N__4559),
            .I(N__4555));
    InMux I__909 (
            .O(N__4558),
            .I(N__4552));
    LocalMux I__908 (
            .O(N__4555),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__907 (
            .O(N__4552),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    CascadeMux I__906 (
            .O(N__4547),
            .I(N__4543));
    InMux I__905 (
            .O(N__4546),
            .I(N__4537));
    InMux I__904 (
            .O(N__4543),
            .I(N__4537));
    InMux I__903 (
            .O(N__4542),
            .I(N__4534));
    LocalMux I__902 (
            .O(N__4537),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__901 (
            .O(N__4534),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    InMux I__900 (
            .O(N__4529),
            .I(N__4525));
    InMux I__899 (
            .O(N__4528),
            .I(N__4522));
    LocalMux I__898 (
            .O(N__4525),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__897 (
            .O(N__4522),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    CascadeMux I__896 (
            .O(N__4517),
            .I(N__4514));
    InMux I__895 (
            .O(N__4514),
            .I(N__4511));
    LocalMux I__894 (
            .O(N__4511),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    CascadeMux I__893 (
            .O(N__4508),
            .I(N__4505));
    InMux I__892 (
            .O(N__4505),
            .I(N__4501));
    InMux I__891 (
            .O(N__4504),
            .I(N__4498));
    LocalMux I__890 (
            .O(N__4501),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__889 (
            .O(N__4498),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    CascadeMux I__888 (
            .O(N__4493),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    CascadeMux I__887 (
            .O(N__4490),
            .I(\U409_TRANSFER_ACK.N_105_cascade_ ));
    InMux I__886 (
            .O(N__4487),
            .I(N__4484));
    LocalMux I__885 (
            .O(N__4484),
            .I(\U409_TRANSFER_ACK.m9_bm ));
    InMux I__884 (
            .O(N__4481),
            .I(N__4475));
    InMux I__883 (
            .O(N__4480),
            .I(N__4475));
    LocalMux I__882 (
            .O(N__4475),
            .I(\U409_TRANSFER_ACK.N_4 ));
    InMux I__881 (
            .O(N__4472),
            .I(N__4469));
    LocalMux I__880 (
            .O(N__4469),
            .I(N__4465));
    InMux I__879 (
            .O(N__4468),
            .I(N__4461));
    Span4Mux_v I__878 (
            .O(N__4465),
            .I(N__4454));
    InMux I__877 (
            .O(N__4464),
            .I(N__4451));
    LocalMux I__876 (
            .O(N__4461),
            .I(N__4448));
    CascadeMux I__875 (
            .O(N__4460),
            .I(N__4445));
    InMux I__874 (
            .O(N__4459),
            .I(N__4442));
    InMux I__873 (
            .O(N__4458),
            .I(N__4439));
    InMux I__872 (
            .O(N__4457),
            .I(N__4436));
    Sp12to4 I__871 (
            .O(N__4454),
            .I(N__4431));
    LocalMux I__870 (
            .O(N__4451),
            .I(N__4431));
    Span4Mux_v I__869 (
            .O(N__4448),
            .I(N__4428));
    InMux I__868 (
            .O(N__4445),
            .I(N__4425));
    LocalMux I__867 (
            .O(N__4442),
            .I(N__4420));
    LocalMux I__866 (
            .O(N__4439),
            .I(N__4420));
    LocalMux I__865 (
            .O(N__4436),
            .I(N__4417));
    Span12Mux_h I__864 (
            .O(N__4431),
            .I(N__4412));
    Sp12to4 I__863 (
            .O(N__4428),
            .I(N__4412));
    LocalMux I__862 (
            .O(N__4425),
            .I(N__4405));
    Sp12to4 I__861 (
            .O(N__4420),
            .I(N__4405));
    Sp12to4 I__860 (
            .O(N__4417),
            .I(N__4405));
    Span12Mux_v I__859 (
            .O(N__4412),
            .I(N__4402));
    Span12Mux_v I__858 (
            .O(N__4405),
            .I(N__4399));
    Odrv12 I__857 (
            .O(N__4402),
            .I(A_c_22));
    Odrv12 I__856 (
            .O(N__4399),
            .I(A_c_22));
    InMux I__855 (
            .O(N__4394),
            .I(N__4389));
    InMux I__854 (
            .O(N__4393),
            .I(N__4386));
    InMux I__853 (
            .O(N__4392),
            .I(N__4381));
    LocalMux I__852 (
            .O(N__4389),
            .I(N__4378));
    LocalMux I__851 (
            .O(N__4386),
            .I(N__4375));
    InMux I__850 (
            .O(N__4385),
            .I(N__4372));
    InMux I__849 (
            .O(N__4384),
            .I(N__4368));
    LocalMux I__848 (
            .O(N__4381),
            .I(N__4362));
    Span4Mux_v I__847 (
            .O(N__4378),
            .I(N__4355));
    Span4Mux_h I__846 (
            .O(N__4375),
            .I(N__4355));
    LocalMux I__845 (
            .O(N__4372),
            .I(N__4355));
    InMux I__844 (
            .O(N__4371),
            .I(N__4352));
    LocalMux I__843 (
            .O(N__4368),
            .I(N__4349));
    InMux I__842 (
            .O(N__4367),
            .I(N__4346));
    InMux I__841 (
            .O(N__4366),
            .I(N__4343));
    InMux I__840 (
            .O(N__4365),
            .I(N__4340));
    Span4Mux_v I__839 (
            .O(N__4362),
            .I(N__4335));
    Span4Mux_v I__838 (
            .O(N__4355),
            .I(N__4335));
    LocalMux I__837 (
            .O(N__4352),
            .I(N__4332));
    Span4Mux_v I__836 (
            .O(N__4349),
            .I(N__4329));
    LocalMux I__835 (
            .O(N__4346),
            .I(N__4326));
    LocalMux I__834 (
            .O(N__4343),
            .I(N__4321));
    LocalMux I__833 (
            .O(N__4340),
            .I(N__4321));
    Span4Mux_h I__832 (
            .O(N__4335),
            .I(N__4316));
    Span4Mux_v I__831 (
            .O(N__4332),
            .I(N__4316));
    Span4Mux_v I__830 (
            .O(N__4329),
            .I(N__4309));
    Span4Mux_v I__829 (
            .O(N__4326),
            .I(N__4309));
    Span4Mux_v I__828 (
            .O(N__4321),
            .I(N__4309));
    Sp12to4 I__827 (
            .O(N__4316),
            .I(N__4304));
    Sp12to4 I__826 (
            .O(N__4309),
            .I(N__4304));
    Odrv12 I__825 (
            .O(N__4304),
            .I(A_c_23));
    InMux I__824 (
            .O(N__4301),
            .I(N__4297));
    InMux I__823 (
            .O(N__4300),
            .I(N__4293));
    LocalMux I__822 (
            .O(N__4297),
            .I(N__4289));
    InMux I__821 (
            .O(N__4296),
            .I(N__4286));
    LocalMux I__820 (
            .O(N__4293),
            .I(N__4283));
    CascadeMux I__819 (
            .O(N__4292),
            .I(N__4278));
    Span4Mux_v I__818 (
            .O(N__4289),
            .I(N__4275));
    LocalMux I__817 (
            .O(N__4286),
            .I(N__4272));
    Span4Mux_h I__816 (
            .O(N__4283),
            .I(N__4269));
    InMux I__815 (
            .O(N__4282),
            .I(N__4266));
    InMux I__814 (
            .O(N__4281),
            .I(N__4261));
    InMux I__813 (
            .O(N__4278),
            .I(N__4261));
    Span4Mux_v I__812 (
            .O(N__4275),
            .I(N__4258));
    Span4Mux_v I__811 (
            .O(N__4272),
            .I(N__4255));
    Span4Mux_h I__810 (
            .O(N__4269),
            .I(N__4248));
    LocalMux I__809 (
            .O(N__4266),
            .I(N__4248));
    LocalMux I__808 (
            .O(N__4261),
            .I(N__4248));
    Span4Mux_h I__807 (
            .O(N__4258),
            .I(N__4245));
    Span4Mux_v I__806 (
            .O(N__4255),
            .I(N__4240));
    Span4Mux_v I__805 (
            .O(N__4248),
            .I(N__4240));
    Sp12to4 I__804 (
            .O(N__4245),
            .I(N__4235));
    Sp12to4 I__803 (
            .O(N__4240),
            .I(N__4235));
    Odrv12 I__802 (
            .O(N__4235),
            .I(A_c_21));
    CascadeMux I__801 (
            .O(N__4232),
            .I(N__4229));
    InMux I__800 (
            .O(N__4229),
            .I(N__4225));
    InMux I__799 (
            .O(N__4228),
            .I(N__4222));
    LocalMux I__798 (
            .O(N__4225),
            .I(N__4217));
    LocalMux I__797 (
            .O(N__4222),
            .I(N__4217));
    Odrv12 I__796 (
            .O(N__4217),
            .I(\U409_ADDRESS_DECODE.LOWROMZ0 ));
    CascadeMux I__795 (
            .O(N__4214),
            .I(N__4210));
    InMux I__794 (
            .O(N__4213),
            .I(N__4207));
    InMux I__793 (
            .O(N__4210),
            .I(N__4204));
    LocalMux I__792 (
            .O(N__4207),
            .I(N__4201));
    LocalMux I__791 (
            .O(N__4204),
            .I(N__4198));
    Span12Mux_v I__790 (
            .O(N__4201),
            .I(N__4195));
    Span4Mux_h I__789 (
            .O(N__4198),
            .I(N__4192));
    Odrv12 I__788 (
            .O(N__4195),
            .I(\U409_ADDRESS_DECODE.HIROMZ0 ));
    Odrv4 I__787 (
            .O(N__4192),
            .I(\U409_ADDRESS_DECODE.HIROMZ0 ));
    IoInMux I__786 (
            .O(N__4187),
            .I(N__4184));
    LocalMux I__785 (
            .O(N__4184),
            .I(N__4181));
    Span4Mux_s0_v I__784 (
            .O(N__4181),
            .I(N__4178));
    Span4Mux_v I__783 (
            .O(N__4178),
            .I(N__4175));
    Sp12to4 I__782 (
            .O(N__4175),
            .I(N__4172));
    Span12Mux_h I__781 (
            .O(N__4172),
            .I(N__4169));
    Odrv12 I__780 (
            .O(N__4169),
            .I(ROMENm_i));
    InMux I__779 (
            .O(N__4166),
            .I(N__4163));
    LocalMux I__778 (
            .O(N__4163),
            .I(N__4160));
    Span4Mux_v I__777 (
            .O(N__4160),
            .I(N__4157));
    Span4Mux_h I__776 (
            .O(N__4157),
            .I(N__4154));
    Odrv4 I__775 (
            .O(N__4154),
            .I(AUTOVECTORm));
    InMux I__774 (
            .O(N__4151),
            .I(N__4145));
    InMux I__773 (
            .O(N__4150),
            .I(N__4145));
    LocalMux I__772 (
            .O(N__4145),
            .I(N__4142));
    Span4Mux_v I__771 (
            .O(N__4142),
            .I(N__4139));
    Span4Mux_v I__770 (
            .O(N__4139),
            .I(N__4135));
    InMux I__769 (
            .O(N__4138),
            .I(N__4132));
    Sp12to4 I__768 (
            .O(N__4135),
            .I(N__4127));
    LocalMux I__767 (
            .O(N__4132),
            .I(N__4127));
    Span12Mux_h I__766 (
            .O(N__4127),
            .I(N__4124));
    Span12Mux_v I__765 (
            .O(N__4124),
            .I(N__4121));
    Odrv12 I__764 (
            .O(N__4121),
            .I(TSn_c));
    IoInMux I__763 (
            .O(N__4118),
            .I(N__4115));
    LocalMux I__762 (
            .O(N__4115),
            .I(N__4111));
    CascadeMux I__761 (
            .O(N__4114),
            .I(N__4107));
    IoSpan4Mux I__760 (
            .O(N__4111),
            .I(N__4102));
    InMux I__759 (
            .O(N__4110),
            .I(N__4099));
    InMux I__758 (
            .O(N__4107),
            .I(N__4096));
    CascadeMux I__757 (
            .O(N__4106),
            .I(N__4093));
    CascadeMux I__756 (
            .O(N__4105),
            .I(N__4090));
    Span4Mux_s0_v I__755 (
            .O(N__4102),
            .I(N__4087));
    LocalMux I__754 (
            .O(N__4099),
            .I(N__4084));
    LocalMux I__753 (
            .O(N__4096),
            .I(N__4081));
    InMux I__752 (
            .O(N__4093),
            .I(N__4078));
    InMux I__751 (
            .O(N__4090),
            .I(N__4075));
    Sp12to4 I__750 (
            .O(N__4087),
            .I(N__4072));
    Span4Mux_v I__749 (
            .O(N__4084),
            .I(N__4065));
    Span4Mux_v I__748 (
            .O(N__4081),
            .I(N__4065));
    LocalMux I__747 (
            .O(N__4078),
            .I(N__4065));
    LocalMux I__746 (
            .O(N__4075),
            .I(N__4062));
    Span12Mux_v I__745 (
            .O(N__4072),
            .I(N__4055));
    Sp12to4 I__744 (
            .O(N__4065),
            .I(N__4055));
    Sp12to4 I__743 (
            .O(N__4062),
            .I(N__4055));
    Span12Mux_v I__742 (
            .O(N__4055),
            .I(N__4052));
    Odrv12 I__741 (
            .O(N__4052),
            .I(CLK40_IN_c));
    InMux I__740 (
            .O(N__4049),
            .I(N__4046));
    LocalMux I__739 (
            .O(N__4046),
            .I(N__4043));
    Odrv4 I__738 (
            .O(N__4043),
            .I(ROMENm));
    IoInMux I__737 (
            .O(N__4040),
            .I(N__4037));
    LocalMux I__736 (
            .O(N__4037),
            .I(N__4034));
    Span4Mux_s3_v I__735 (
            .O(N__4034),
            .I(N__4031));
    Span4Mux_h I__734 (
            .O(N__4031),
            .I(N__4028));
    Odrv4 I__733 (
            .O(N__4028),
            .I(CONSTANT_ONE_NET));
    InMux I__732 (
            .O(N__4025),
            .I(N__4022));
    LocalMux I__731 (
            .O(N__4022),
            .I(N__4019));
    Span12Mux_s10_v I__730 (
            .O(N__4019),
            .I(N__4016));
    Span12Mux_h I__729 (
            .O(N__4016),
            .I(N__4013));
    Odrv12 I__728 (
            .O(N__4013),
            .I(A_c_12));
    IoInMux I__727 (
            .O(N__4010),
            .I(N__4007));
    LocalMux I__726 (
            .O(N__4007),
            .I(N__4004));
    IoSpan4Mux I__725 (
            .O(N__4004),
            .I(N__4001));
    Span4Mux_s3_h I__724 (
            .O(N__4001),
            .I(N__3998));
    Span4Mux_v I__723 (
            .O(N__3998),
            .I(N__3995));
    Span4Mux_h I__722 (
            .O(N__3995),
            .I(N__3992));
    Sp12to4 I__721 (
            .O(N__3992),
            .I(N__3989));
    Odrv12 I__720 (
            .O(N__3989),
            .I(U409_ADDRESS_DECODE_un1_nCIACS0_i));
    CascadeMux I__719 (
            .O(N__3986),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    CascadeMux I__718 (
            .O(N__3983),
            .I(N__3979));
    InMux I__717 (
            .O(N__3982),
            .I(N__3976));
    InMux I__716 (
            .O(N__3979),
            .I(N__3973));
    LocalMux I__715 (
            .O(N__3976),
            .I(N__3965));
    LocalMux I__714 (
            .O(N__3973),
            .I(N__3962));
    InMux I__713 (
            .O(N__3972),
            .I(N__3951));
    InMux I__712 (
            .O(N__3971),
            .I(N__3951));
    InMux I__711 (
            .O(N__3970),
            .I(N__3951));
    InMux I__710 (
            .O(N__3969),
            .I(N__3951));
    InMux I__709 (
            .O(N__3968),
            .I(N__3951));
    Odrv4 I__708 (
            .O(N__3965),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    Odrv4 I__707 (
            .O(N__3962),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__706 (
            .O(N__3951),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    InMux I__705 (
            .O(N__3944),
            .I(N__3937));
    InMux I__704 (
            .O(N__3943),
            .I(N__3934));
    InMux I__703 (
            .O(N__3942),
            .I(N__3927));
    InMux I__702 (
            .O(N__3941),
            .I(N__3927));
    InMux I__701 (
            .O(N__3940),
            .I(N__3927));
    LocalMux I__700 (
            .O(N__3937),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__699 (
            .O(N__3934),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__698 (
            .O(N__3927),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    InMux I__697 (
            .O(N__3920),
            .I(N__3914));
    InMux I__696 (
            .O(N__3919),
            .I(N__3911));
    InMux I__695 (
            .O(N__3918),
            .I(N__3906));
    InMux I__694 (
            .O(N__3917),
            .I(N__3906));
    LocalMux I__693 (
            .O(N__3914),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__692 (
            .O(N__3911),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__691 (
            .O(N__3906),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    InMux I__690 (
            .O(N__3899),
            .I(N__3896));
    LocalMux I__689 (
            .O(N__3896),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    InMux I__688 (
            .O(N__3893),
            .I(N__3888));
    InMux I__687 (
            .O(N__3892),
            .I(N__3883));
    InMux I__686 (
            .O(N__3891),
            .I(N__3883));
    LocalMux I__685 (
            .O(N__3888),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    LocalMux I__684 (
            .O(N__3883),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    CascadeMux I__683 (
            .O(N__3878),
            .I(\U409_TRANSFER_ACK.m9_am_cascade_ ));
    CascadeMux I__682 (
            .O(N__3875),
            .I(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ));
    CascadeMux I__681 (
            .O(N__3872),
            .I(N__3869));
    InMux I__680 (
            .O(N__3869),
            .I(N__3866));
    LocalMux I__679 (
            .O(N__3866),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__678 (
            .O(N__3863),
            .I(N__3860));
    LocalMux I__677 (
            .O(N__3860),
            .I(N__3857));
    Odrv4 I__676 (
            .O(N__3857),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ));
    InMux I__675 (
            .O(N__3854),
            .I(N__3851));
    LocalMux I__674 (
            .O(N__3851),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3 ));
    InMux I__673 (
            .O(N__3848),
            .I(N__3844));
    InMux I__672 (
            .O(N__3847),
            .I(N__3840));
    LocalMux I__671 (
            .O(N__3844),
            .I(N__3837));
    InMux I__670 (
            .O(N__3843),
            .I(N__3834));
    LocalMux I__669 (
            .O(N__3840),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    Odrv4 I__668 (
            .O(N__3837),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__667 (
            .O(N__3834),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    InMux I__666 (
            .O(N__3827),
            .I(N__3821));
    InMux I__665 (
            .O(N__3826),
            .I(N__3818));
    InMux I__664 (
            .O(N__3825),
            .I(N__3815));
    InMux I__663 (
            .O(N__3824),
            .I(N__3812));
    LocalMux I__662 (
            .O(N__3821),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__661 (
            .O(N__3818),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__660 (
            .O(N__3815),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__659 (
            .O(N__3812),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__658 (
            .O(N__3803),
            .I(N__3798));
    InMux I__657 (
            .O(N__3802),
            .I(N__3792));
    InMux I__656 (
            .O(N__3801),
            .I(N__3792));
    InMux I__655 (
            .O(N__3798),
            .I(N__3787));
    InMux I__654 (
            .O(N__3797),
            .I(N__3787));
    LocalMux I__653 (
            .O(N__3792),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__652 (
            .O(N__3787),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    CascadeMux I__651 (
            .O(N__3782),
            .I(N__3777));
    InMux I__650 (
            .O(N__3781),
            .I(N__3773));
    InMux I__649 (
            .O(N__3780),
            .I(N__3770));
    InMux I__648 (
            .O(N__3777),
            .I(N__3767));
    InMux I__647 (
            .O(N__3776),
            .I(N__3764));
    LocalMux I__646 (
            .O(N__3773),
            .I(N__3761));
    LocalMux I__645 (
            .O(N__3770),
            .I(N__3756));
    LocalMux I__644 (
            .O(N__3767),
            .I(N__3756));
    LocalMux I__643 (
            .O(N__3764),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    Odrv4 I__642 (
            .O(N__3761),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    Odrv4 I__641 (
            .O(N__3756),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    InMux I__640 (
            .O(N__3749),
            .I(N__3742));
    InMux I__639 (
            .O(N__3748),
            .I(N__3737));
    InMux I__638 (
            .O(N__3747),
            .I(N__3737));
    InMux I__637 (
            .O(N__3746),
            .I(N__3734));
    InMux I__636 (
            .O(N__3745),
            .I(N__3731));
    LocalMux I__635 (
            .O(N__3742),
            .I(N__3728));
    LocalMux I__634 (
            .O(N__3737),
            .I(N__3723));
    LocalMux I__633 (
            .O(N__3734),
            .I(N__3723));
    LocalMux I__632 (
            .O(N__3731),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    Odrv4 I__631 (
            .O(N__3728),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    Odrv4 I__630 (
            .O(N__3723),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    CascadeMux I__629 (
            .O(N__3716),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ));
    CascadeMux I__628 (
            .O(N__3713),
            .I(N__3710));
    InMux I__627 (
            .O(N__3710),
            .I(N__3704));
    InMux I__626 (
            .O(N__3709),
            .I(N__3704));
    LocalMux I__625 (
            .O(N__3704),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    CascadeMux I__624 (
            .O(N__3701),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ));
    CascadeMux I__623 (
            .O(N__3698),
            .I(N__3694));
    CascadeMux I__622 (
            .O(N__3697),
            .I(N__3689));
    InMux I__621 (
            .O(N__3694),
            .I(N__3683));
    InMux I__620 (
            .O(N__3693),
            .I(N__3683));
    InMux I__619 (
            .O(N__3692),
            .I(N__3676));
    InMux I__618 (
            .O(N__3689),
            .I(N__3676));
    InMux I__617 (
            .O(N__3688),
            .I(N__3676));
    LocalMux I__616 (
            .O(N__3683),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__615 (
            .O(N__3676),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    InMux I__614 (
            .O(N__3671),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__613 (
            .O(N__3668),
            .I(bfn_11_6_0_));
    InMux I__612 (
            .O(N__3665),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__611 (
            .O(N__3662),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__610 (
            .O(N__3659),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__609 (
            .O(N__3656),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__608 (
            .O(N__3653),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__607 (
            .O(N__3650),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__606 (
            .O(N__3647),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__605 (
            .O(N__3644),
            .I(N__3641));
    LocalMux I__604 (
            .O(N__3641),
            .I(N__3638));
    Span4Mux_v I__603 (
            .O(N__3638),
            .I(N__3633));
    InMux I__602 (
            .O(N__3637),
            .I(N__3630));
    InMux I__601 (
            .O(N__3636),
            .I(N__3627));
    Span4Mux_h I__600 (
            .O(N__3633),
            .I(N__3624));
    LocalMux I__599 (
            .O(N__3630),
            .I(N__3621));
    LocalMux I__598 (
            .O(N__3627),
            .I(N__3618));
    Odrv4 I__597 (
            .O(N__3624),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ));
    Odrv12 I__596 (
            .O(N__3621),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ));
    Odrv12 I__595 (
            .O(N__3618),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ));
    IoInMux I__594 (
            .O(N__3611),
            .I(N__3608));
    LocalMux I__593 (
            .O(N__3608),
            .I(N__3605));
    IoSpan4Mux I__592 (
            .O(N__3605),
            .I(N__3602));
    Sp12to4 I__591 (
            .O(N__3602),
            .I(N__3599));
    Span12Mux_s6_v I__590 (
            .O(N__3599),
            .I(N__3596));
    Span12Mux_h I__589 (
            .O(N__3596),
            .I(N__3593));
    Odrv12 I__588 (
            .O(N__3593),
            .I(U409_ADDRESS_DECODE_un1_nREGSPACE_i));
    InMux I__587 (
            .O(N__3590),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__586 (
            .O(N__3587),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__585 (
            .O(N__3584),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__584 (
            .O(N__3581),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    InMux I__583 (
            .O(N__3578),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__582 (
            .O(N__3575),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    IoInMux I__581 (
            .O(N__3572),
            .I(N__3569));
    LocalMux I__580 (
            .O(N__3569),
            .I(N__3566));
    Span4Mux_s1_v I__579 (
            .O(N__3566),
            .I(N__3563));
    Sp12to4 I__578 (
            .O(N__3563),
            .I(N__3560));
    Span12Mux_h I__577 (
            .O(N__3560),
            .I(N__3556));
    InMux I__576 (
            .O(N__3559),
            .I(N__3553));
    Odrv12 I__575 (
            .O(N__3556),
            .I(TICK50_c));
    LocalMux I__574 (
            .O(N__3553),
            .I(TICK50_c));
    InMux I__573 (
            .O(N__3548),
            .I(N__3533));
    InMux I__572 (
            .O(N__3547),
            .I(N__3533));
    InMux I__571 (
            .O(N__3546),
            .I(N__3533));
    InMux I__570 (
            .O(N__3545),
            .I(N__3533));
    CascadeMux I__569 (
            .O(N__3544),
            .I(N__3530));
    InMux I__568 (
            .O(N__3543),
            .I(N__3526));
    InMux I__567 (
            .O(N__3542),
            .I(N__3523));
    LocalMux I__566 (
            .O(N__3533),
            .I(N__3520));
    InMux I__565 (
            .O(N__3530),
            .I(N__3515));
    InMux I__564 (
            .O(N__3529),
            .I(N__3515));
    LocalMux I__563 (
            .O(N__3526),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__562 (
            .O(N__3523),
            .I(\U409_TICK.TICK503_14 ));
    Odrv4 I__561 (
            .O(N__3520),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__560 (
            .O(N__3515),
            .I(\U409_TICK.TICK503_14 ));
    CascadeMux I__559 (
            .O(N__3506),
            .I(N__3503));
    InMux I__558 (
            .O(N__3503),
            .I(N__3493));
    InMux I__557 (
            .O(N__3502),
            .I(N__3486));
    InMux I__556 (
            .O(N__3501),
            .I(N__3486));
    InMux I__555 (
            .O(N__3500),
            .I(N__3486));
    InMux I__554 (
            .O(N__3499),
            .I(N__3483));
    InMux I__553 (
            .O(N__3498),
            .I(N__3476));
    InMux I__552 (
            .O(N__3497),
            .I(N__3476));
    InMux I__551 (
            .O(N__3496),
            .I(N__3476));
    LocalMux I__550 (
            .O(N__3493),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__549 (
            .O(N__3486),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__548 (
            .O(N__3483),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__547 (
            .O(N__3476),
            .I(\U409_TICK.TICK503_9 ));
    CascadeMux I__546 (
            .O(N__3467),
            .I(N__3461));
    CascadeMux I__545 (
            .O(N__3466),
            .I(N__3457));
    CascadeMux I__544 (
            .O(N__3465),
            .I(N__3454));
    CascadeMux I__543 (
            .O(N__3464),
            .I(N__3451));
    InMux I__542 (
            .O(N__3461),
            .I(N__3445));
    InMux I__541 (
            .O(N__3460),
            .I(N__3442));
    InMux I__540 (
            .O(N__3457),
            .I(N__3435));
    InMux I__539 (
            .O(N__3454),
            .I(N__3435));
    InMux I__538 (
            .O(N__3451),
            .I(N__3435));
    InMux I__537 (
            .O(N__3450),
            .I(N__3432));
    InMux I__536 (
            .O(N__3449),
            .I(N__3427));
    InMux I__535 (
            .O(N__3448),
            .I(N__3427));
    LocalMux I__534 (
            .O(N__3445),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__533 (
            .O(N__3442),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__532 (
            .O(N__3435),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__531 (
            .O(N__3432),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__530 (
            .O(N__3427),
            .I(\U409_TICK.TICK503_10 ));
    InMux I__529 (
            .O(N__3416),
            .I(N__3413));
    LocalMux I__528 (
            .O(N__3413),
            .I(N__3410));
    Odrv4 I__527 (
            .O(N__3410),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__526 (
            .O(N__3407),
            .I(N__3403));
    InMux I__525 (
            .O(N__3406),
            .I(N__3400));
    LocalMux I__524 (
            .O(N__3403),
            .I(N__3397));
    LocalMux I__523 (
            .O(N__3400),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    Odrv4 I__522 (
            .O(N__3397),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__521 (
            .O(N__3392),
            .I(N__3386));
    InMux I__520 (
            .O(N__3391),
            .I(N__3386));
    LocalMux I__519 (
            .O(N__3386),
            .I(N__3383));
    Odrv4 I__518 (
            .O(N__3383),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ));
    CascadeMux I__517 (
            .O(N__3380),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_ ));
    CascadeMux I__516 (
            .O(N__3377),
            .I(N__3374));
    InMux I__515 (
            .O(N__3374),
            .I(N__3368));
    InMux I__514 (
            .O(N__3373),
            .I(N__3368));
    LocalMux I__513 (
            .O(N__3368),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    InMux I__512 (
            .O(N__3365),
            .I(N__3362));
    LocalMux I__511 (
            .O(N__3362),
            .I(\U409_TICK.TICK503_11 ));
    InMux I__510 (
            .O(N__3359),
            .I(N__3355));
    InMux I__509 (
            .O(N__3358),
            .I(N__3352));
    LocalMux I__508 (
            .O(N__3355),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__507 (
            .O(N__3352),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    CascadeMux I__506 (
            .O(N__3347),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    InMux I__505 (
            .O(N__3344),
            .I(N__3341));
    LocalMux I__504 (
            .O(N__3341),
            .I(N__3337));
    InMux I__503 (
            .O(N__3340),
            .I(N__3334));
    Odrv4 I__502 (
            .O(N__3337),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__501 (
            .O(N__3334),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    CascadeMux I__500 (
            .O(N__3329),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    InMux I__499 (
            .O(N__3326),
            .I(N__3323));
    LocalMux I__498 (
            .O(N__3323),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    CascadeMux I__497 (
            .O(N__3320),
            .I(N__3316));
    CascadeMux I__496 (
            .O(N__3319),
            .I(N__3313));
    InMux I__495 (
            .O(N__3316),
            .I(N__3307));
    InMux I__494 (
            .O(N__3313),
            .I(N__3307));
    InMux I__493 (
            .O(N__3312),
            .I(N__3304));
    LocalMux I__492 (
            .O(N__3307),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__491 (
            .O(N__3304),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    CascadeMux I__490 (
            .O(N__3299),
            .I(N__3293));
    InMux I__489 (
            .O(N__3298),
            .I(N__3286));
    InMux I__488 (
            .O(N__3297),
            .I(N__3286));
    InMux I__487 (
            .O(N__3296),
            .I(N__3286));
    InMux I__486 (
            .O(N__3293),
            .I(N__3283));
    LocalMux I__485 (
            .O(N__3286),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__484 (
            .O(N__3283),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__483 (
            .O(N__3278),
            .I(N__3275));
    LocalMux I__482 (
            .O(N__3275),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    CascadeMux I__481 (
            .O(N__3272),
            .I(N__3269));
    InMux I__480 (
            .O(N__3269),
            .I(N__3265));
    InMux I__479 (
            .O(N__3268),
            .I(N__3262));
    LocalMux I__478 (
            .O(N__3265),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__477 (
            .O(N__3262),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    CascadeMux I__476 (
            .O(N__3257),
            .I(N__3254));
    InMux I__475 (
            .O(N__3254),
            .I(N__3251));
    LocalMux I__474 (
            .O(N__3251),
            .I(N__3247));
    InMux I__473 (
            .O(N__3250),
            .I(N__3244));
    Odrv4 I__472 (
            .O(N__3247),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__471 (
            .O(N__3244),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    CascadeMux I__470 (
            .O(N__3239),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    InMux I__469 (
            .O(N__3236),
            .I(N__3233));
    LocalMux I__468 (
            .O(N__3233),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__467 (
            .O(N__3230),
            .I(N__3226));
    InMux I__466 (
            .O(N__3229),
            .I(N__3223));
    LocalMux I__465 (
            .O(N__3226),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__464 (
            .O(N__3223),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    InMux I__463 (
            .O(N__3218),
            .I(N__3215));
    LocalMux I__462 (
            .O(N__3215),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__461 (
            .O(N__3212),
            .I(N__3208));
    InMux I__460 (
            .O(N__3211),
            .I(N__3205));
    LocalMux I__459 (
            .O(N__3208),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__458 (
            .O(N__3205),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    InMux I__457 (
            .O(N__3200),
            .I(N__3197));
    LocalMux I__456 (
            .O(N__3197),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__455 (
            .O(N__3194),
            .I(N__3190));
    InMux I__454 (
            .O(N__3193),
            .I(N__3187));
    LocalMux I__453 (
            .O(N__3190),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__452 (
            .O(N__3187),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__451 (
            .O(N__3182),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__450 (
            .O(N__3179),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__449 (
            .O(N__3176),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__448 (
            .O(N__3173),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__447 (
            .O(N__3170),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__446 (
            .O(N__3167),
            .I(N__3163));
    InMux I__445 (
            .O(N__3166),
            .I(N__3160));
    LocalMux I__444 (
            .O(N__3163),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__443 (
            .O(N__3160),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    InMux I__442 (
            .O(N__3155),
            .I(N__3151));
    InMux I__441 (
            .O(N__3154),
            .I(N__3148));
    LocalMux I__440 (
            .O(N__3151),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__439 (
            .O(N__3148),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__438 (
            .O(N__3143),
            .I(N__3139));
    InMux I__437 (
            .O(N__3142),
            .I(N__3136));
    LocalMux I__436 (
            .O(N__3139),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__435 (
            .O(N__3136),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__434 (
            .O(N__3131),
            .I(N__3127));
    InMux I__433 (
            .O(N__3130),
            .I(N__3124));
    LocalMux I__432 (
            .O(N__3127),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__431 (
            .O(N__3124),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    InMux I__430 (
            .O(N__3119),
            .I(N__3115));
    InMux I__429 (
            .O(N__3118),
            .I(N__3112));
    LocalMux I__428 (
            .O(N__3115),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__427 (
            .O(N__3112),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    CascadeMux I__426 (
            .O(N__3107),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    InMux I__425 (
            .O(N__3104),
            .I(N__3101));
    LocalMux I__424 (
            .O(N__3101),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__423 (
            .O(N__3098),
            .I(N__3094));
    InMux I__422 (
            .O(N__3097),
            .I(N__3091));
    LocalMux I__421 (
            .O(N__3094),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__420 (
            .O(N__3091),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__419 (
            .O(N__3086),
            .I(N__3082));
    InMux I__418 (
            .O(N__3085),
            .I(N__3079));
    LocalMux I__417 (
            .O(N__3082),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__416 (
            .O(N__3079),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__415 (
            .O(N__3074),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    InMux I__414 (
            .O(N__3071),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__413 (
            .O(N__3068),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    InMux I__412 (
            .O(N__3065),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__411 (
            .O(N__3062),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__410 (
            .O(N__3059),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__409 (
            .O(N__3056),
            .I(bfn_8_6_0_));
    InMux I__408 (
            .O(N__3053),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__407 (
            .O(N__3050),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    CascadeMux I__406 (
            .O(N__3047),
            .I(N__3044));
    InMux I__405 (
            .O(N__3044),
            .I(N__3038));
    InMux I__404 (
            .O(N__3043),
            .I(N__3038));
    LocalMux I__403 (
            .O(N__3038),
            .I(N__3034));
    InMux I__402 (
            .O(N__3037),
            .I(N__3031));
    Span4Mux_v I__401 (
            .O(N__3034),
            .I(N__3026));
    LocalMux I__400 (
            .O(N__3031),
            .I(N__3026));
    Span4Mux_v I__399 (
            .O(N__3026),
            .I(N__3023));
    Odrv4 I__398 (
            .O(N__3023),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEm_6 ));
    CascadeMux I__397 (
            .O(N__3020),
            .I(N__3017));
    InMux I__396 (
            .O(N__3017),
            .I(N__3014));
    LocalMux I__395 (
            .O(N__3014),
            .I(N__3010));
    InMux I__394 (
            .O(N__3013),
            .I(N__3007));
    Span4Mux_v I__393 (
            .O(N__3010),
            .I(N__3004));
    LocalMux I__392 (
            .O(N__3007),
            .I(N__3001));
    Span4Mux_v I__391 (
            .O(N__3004),
            .I(N__2994));
    Span4Mux_v I__390 (
            .O(N__3001),
            .I(N__2994));
    InMux I__389 (
            .O(N__3000),
            .I(N__2991));
    InMux I__388 (
            .O(N__2999),
            .I(N__2988));
    Sp12to4 I__387 (
            .O(N__2994),
            .I(N__2981));
    LocalMux I__386 (
            .O(N__2991),
            .I(N__2981));
    LocalMux I__385 (
            .O(N__2988),
            .I(N__2981));
    Odrv12 I__384 (
            .O(N__2981),
            .I(A_c_20));
    InMux I__383 (
            .O(N__2978),
            .I(N__2975));
    LocalMux I__382 (
            .O(N__2975),
            .I(N__2972));
    Odrv12 I__381 (
            .O(N__2972),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_0 ));
    InMux I__380 (
            .O(N__2969),
            .I(N__2966));
    LocalMux I__379 (
            .O(N__2966),
            .I(N__2963));
    Span4Mux_v I__378 (
            .O(N__2963),
            .I(N__2960));
    Span4Mux_v I__377 (
            .O(N__2960),
            .I(N__2957));
    IoSpan4Mux I__376 (
            .O(N__2957),
            .I(N__2954));
    Odrv4 I__375 (
            .O(N__2954),
            .I(TT_c_1));
    InMux I__374 (
            .O(N__2951),
            .I(N__2948));
    LocalMux I__373 (
            .O(N__2948),
            .I(N__2945));
    Span4Mux_h I__372 (
            .O(N__2945),
            .I(N__2942));
    Span4Mux_v I__371 (
            .O(N__2942),
            .I(N__2939));
    Span4Mux_v I__370 (
            .O(N__2939),
            .I(N__2936));
    Odrv4 I__369 (
            .O(N__2936),
            .I(TT_c_0));
    InMux I__368 (
            .O(N__2933),
            .I(N__2930));
    LocalMux I__367 (
            .O(N__2930),
            .I(N__2927));
    Odrv4 I__366 (
            .O(N__2927),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9 ));
    InMux I__365 (
            .O(N__2924),
            .I(N__2921));
    LocalMux I__364 (
            .O(N__2921),
            .I(N__2918));
    Span12Mux_v I__363 (
            .O(N__2918),
            .I(N__2915));
    Odrv12 I__362 (
            .O(N__2915),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_1Z0Z_0 ));
    CascadeMux I__361 (
            .O(N__2912),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEm_cascade_ ));
    IoInMux I__360 (
            .O(N__2909),
            .I(N__2906));
    LocalMux I__359 (
            .O(N__2906),
            .I(N__2903));
    Span12Mux_s9_v I__358 (
            .O(N__2903),
            .I(N__2900));
    Odrv12 I__357 (
            .O(N__2900),
            .I(PORTSIZE_0_i));
    InMux I__356 (
            .O(N__2897),
            .I(N__2894));
    LocalMux I__355 (
            .O(N__2894),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEm_3 ));
    InMux I__354 (
            .O(N__2891),
            .I(N__2886));
    InMux I__353 (
            .O(N__2890),
            .I(N__2883));
    InMux I__352 (
            .O(N__2889),
            .I(N__2880));
    LocalMux I__351 (
            .O(N__2886),
            .I(N__2877));
    LocalMux I__350 (
            .O(N__2883),
            .I(N__2872));
    LocalMux I__349 (
            .O(N__2880),
            .I(N__2872));
    Span12Mux_h I__348 (
            .O(N__2877),
            .I(N__2869));
    Span12Mux_h I__347 (
            .O(N__2872),
            .I(N__2866));
    Span12Mux_v I__346 (
            .O(N__2869),
            .I(N__2863));
    Span12Mux_v I__345 (
            .O(N__2866),
            .I(N__2860));
    Odrv12 I__344 (
            .O(N__2863),
            .I(A_c_19));
    Odrv12 I__343 (
            .O(N__2860),
            .I(A_c_19));
    InMux I__342 (
            .O(N__2855),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    CascadeMux I__341 (
            .O(N__2852),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_ ));
    InMux I__340 (
            .O(N__2849),
            .I(N__2846));
    LocalMux I__339 (
            .O(N__2846),
            .I(N__2843));
    Span4Mux_v I__338 (
            .O(N__2843),
            .I(N__2838));
    InMux I__337 (
            .O(N__2842),
            .I(N__2833));
    InMux I__336 (
            .O(N__2841),
            .I(N__2833));
    Span4Mux_v I__335 (
            .O(N__2838),
            .I(N__2828));
    LocalMux I__334 (
            .O(N__2833),
            .I(N__2828));
    Span4Mux_v I__333 (
            .O(N__2828),
            .I(N__2825));
    Span4Mux_v I__332 (
            .O(N__2825),
            .I(N__2822));
    Span4Mux_h I__331 (
            .O(N__2822),
            .I(N__2819));
    Odrv4 I__330 (
            .O(N__2819),
            .I(A_c_26));
    InMux I__329 (
            .O(N__2816),
            .I(N__2813));
    LocalMux I__328 (
            .O(N__2813),
            .I(N__2810));
    Span4Mux_v I__327 (
            .O(N__2810),
            .I(N__2805));
    InMux I__326 (
            .O(N__2809),
            .I(N__2800));
    InMux I__325 (
            .O(N__2808),
            .I(N__2800));
    Sp12to4 I__324 (
            .O(N__2805),
            .I(N__2795));
    LocalMux I__323 (
            .O(N__2800),
            .I(N__2795));
    Odrv12 I__322 (
            .O(N__2795),
            .I(A_c_27));
    InMux I__321 (
            .O(N__2792),
            .I(N__2789));
    LocalMux I__320 (
            .O(N__2789),
            .I(N__2785));
    CascadeMux I__319 (
            .O(N__2788),
            .I(N__2781));
    Span4Mux_v I__318 (
            .O(N__2785),
            .I(N__2778));
    InMux I__317 (
            .O(N__2784),
            .I(N__2773));
    InMux I__316 (
            .O(N__2781),
            .I(N__2773));
    Sp12to4 I__315 (
            .O(N__2778),
            .I(N__2768));
    LocalMux I__314 (
            .O(N__2773),
            .I(N__2768));
    Odrv12 I__313 (
            .O(N__2768),
            .I(A_c_25));
    InMux I__312 (
            .O(N__2765),
            .I(N__2760));
    InMux I__311 (
            .O(N__2764),
            .I(N__2755));
    InMux I__310 (
            .O(N__2763),
            .I(N__2755));
    LocalMux I__309 (
            .O(N__2760),
            .I(N__2750));
    LocalMux I__308 (
            .O(N__2755),
            .I(N__2750));
    Span4Mux_v I__307 (
            .O(N__2750),
            .I(N__2747));
    Span4Mux_v I__306 (
            .O(N__2747),
            .I(N__2744));
    Sp12to4 I__305 (
            .O(N__2744),
            .I(N__2741));
    Odrv12 I__304 (
            .O(N__2741),
            .I(A_c_24));
    InMux I__303 (
            .O(N__2738),
            .I(N__2735));
    LocalMux I__302 (
            .O(N__2735),
            .I(N__2732));
    Odrv4 I__301 (
            .O(N__2732),
            .I(\U409_CIA.g0Z0Z_10 ));
    InMux I__300 (
            .O(N__2729),
            .I(N__2720));
    InMux I__299 (
            .O(N__2728),
            .I(N__2720));
    InMux I__298 (
            .O(N__2727),
            .I(N__2720));
    LocalMux I__297 (
            .O(N__2720),
            .I(N__2717));
    Span4Mux_v I__296 (
            .O(N__2717),
            .I(N__2714));
    Sp12to4 I__295 (
            .O(N__2714),
            .I(N__2711));
    Odrv12 I__294 (
            .O(N__2711),
            .I(A_c_31));
    InMux I__293 (
            .O(N__2708),
            .I(N__2699));
    InMux I__292 (
            .O(N__2707),
            .I(N__2699));
    InMux I__291 (
            .O(N__2706),
            .I(N__2699));
    LocalMux I__290 (
            .O(N__2699),
            .I(N__2696));
    Span4Mux_v I__289 (
            .O(N__2696),
            .I(N__2693));
    Span4Mux_v I__288 (
            .O(N__2693),
            .I(N__2690));
    Sp12to4 I__287 (
            .O(N__2690),
            .I(N__2687));
    Odrv12 I__286 (
            .O(N__2687),
            .I(A_c_28));
    InMux I__285 (
            .O(N__2684),
            .I(N__2680));
    CascadeMux I__284 (
            .O(N__2683),
            .I(N__2677));
    LocalMux I__283 (
            .O(N__2680),
            .I(N__2673));
    InMux I__282 (
            .O(N__2677),
            .I(N__2668));
    InMux I__281 (
            .O(N__2676),
            .I(N__2668));
    Span4Mux_h I__280 (
            .O(N__2673),
            .I(N__2663));
    LocalMux I__279 (
            .O(N__2668),
            .I(N__2663));
    Span4Mux_v I__278 (
            .O(N__2663),
            .I(N__2660));
    Span4Mux_h I__277 (
            .O(N__2660),
            .I(N__2657));
    Odrv4 I__276 (
            .O(N__2657),
            .I(A_c_30));
    CascadeMux I__275 (
            .O(N__2654),
            .I(N__2650));
    CascadeMux I__274 (
            .O(N__2653),
            .I(N__2646));
    InMux I__273 (
            .O(N__2650),
            .I(N__2639));
    InMux I__272 (
            .O(N__2649),
            .I(N__2639));
    InMux I__271 (
            .O(N__2646),
            .I(N__2639));
    LocalMux I__270 (
            .O(N__2639),
            .I(N__2636));
    Span4Mux_h I__269 (
            .O(N__2636),
            .I(N__2633));
    Span4Mux_v I__268 (
            .O(N__2633),
            .I(N__2630));
    Odrv4 I__267 (
            .O(N__2630),
            .I(A_c_29));
    InMux I__266 (
            .O(N__2627),
            .I(N__2624));
    LocalMux I__265 (
            .O(N__2624),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ));
    InMux I__264 (
            .O(N__2621),
            .I(N__2618));
    LocalMux I__263 (
            .O(N__2618),
            .I(\U409_CIA.g0Z0Z_8 ));
    CascadeMux I__262 (
            .O(N__2615),
            .I(N__2612));
    InMux I__261 (
            .O(N__2612),
            .I(N__2609));
    LocalMux I__260 (
            .O(N__2609),
            .I(N__2605));
    InMux I__259 (
            .O(N__2608),
            .I(N__2602));
    Span4Mux_h I__258 (
            .O(N__2605),
            .I(N__2597));
    LocalMux I__257 (
            .O(N__2602),
            .I(N__2597));
    Span4Mux_v I__256 (
            .O(N__2597),
            .I(N__2594));
    Span4Mux_h I__255 (
            .O(N__2594),
            .I(N__2591));
    Span4Mux_v I__254 (
            .O(N__2591),
            .I(N__2588));
    Odrv4 I__253 (
            .O(N__2588),
            .I(A_c_16));
    InMux I__252 (
            .O(N__2585),
            .I(N__2582));
    LocalMux I__251 (
            .O(N__2582),
            .I(\U409_CIA.g0Z0Z_11 ));
    InMux I__250 (
            .O(N__2579),
            .I(N__2576));
    LocalMux I__249 (
            .O(N__2576),
            .I(N__2573));
    Span4Mux_h I__248 (
            .O(N__2573),
            .I(N__2570));
    Odrv4 I__247 (
            .O(N__2570),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8 ));
    InMux I__246 (
            .O(N__2567),
            .I(N__2564));
    LocalMux I__245 (
            .O(N__2564),
            .I(N__2561));
    Odrv12 I__244 (
            .O(N__2561),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7 ));
    CascadeMux I__243 (
            .O(N__2558),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEm_3_cascade_ ));
    CascadeMux I__242 (
            .O(N__2555),
            .I(N__2551));
    InMux I__241 (
            .O(N__2554),
            .I(N__2548));
    InMux I__240 (
            .O(N__2551),
            .I(N__2545));
    LocalMux I__239 (
            .O(N__2548),
            .I(N__2540));
    LocalMux I__238 (
            .O(N__2545),
            .I(N__2540));
    Span4Mux_v I__237 (
            .O(N__2540),
            .I(N__2537));
    Span4Mux_h I__236 (
            .O(N__2537),
            .I(N__2534));
    Span4Mux_v I__235 (
            .O(N__2534),
            .I(N__2531));
    Span4Mux_v I__234 (
            .O(N__2531),
            .I(N__2528));
    Odrv4 I__233 (
            .O(N__2528),
            .I(A_c_18));
    InMux I__232 (
            .O(N__2525),
            .I(N__2519));
    InMux I__231 (
            .O(N__2524),
            .I(N__2519));
    LocalMux I__230 (
            .O(N__2519),
            .I(N__2516));
    Sp12to4 I__229 (
            .O(N__2516),
            .I(N__2513));
    Span12Mux_v I__228 (
            .O(N__2513),
            .I(N__2510));
    Odrv12 I__227 (
            .O(N__2510),
            .I(A_c_17));
    CascadeMux I__226 (
            .O(N__2507),
            .I(\U409_CIA.g0Z0Z_2_cascade_ ));
    ClkMux I__225 (
            .O(N__2504),
            .I(N__2474));
    ClkMux I__224 (
            .O(N__2503),
            .I(N__2474));
    ClkMux I__223 (
            .O(N__2502),
            .I(N__2474));
    ClkMux I__222 (
            .O(N__2501),
            .I(N__2474));
    ClkMux I__221 (
            .O(N__2500),
            .I(N__2474));
    ClkMux I__220 (
            .O(N__2499),
            .I(N__2474));
    ClkMux I__219 (
            .O(N__2498),
            .I(N__2474));
    ClkMux I__218 (
            .O(N__2497),
            .I(N__2474));
    ClkMux I__217 (
            .O(N__2496),
            .I(N__2474));
    ClkMux I__216 (
            .O(N__2495),
            .I(N__2474));
    GlobalMux I__215 (
            .O(N__2474),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.TACK_EN_iC  (
            .O(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .I(N__2504));
    INV \INVU409_TRANSFER_ACK.TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .I(N__2503));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .I(N__2502));
    INV \INVU409_TRANSFER_ACK.LASTCLK_0C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .I(N__2498));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .I(N__2495));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__2501));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .I(N__2500));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .I(N__2497));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .I(N__2499));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .I(N__2496));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_7_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_1_7_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_1_7_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_1_7_0  (
            .in0(N__2608),
            .in1(N__2889),
            .in2(N__2555),
            .in3(N__2524),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_11_LC_1_7_2 .C_ON=1'b0;
    defparam \U409_CIA.g0_11_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_11_LC_1_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.g0_11_LC_1_7_2  (
            .in0(N__4384),
            .in1(N__4296),
            .in2(N__3020),
            .in3(N__2554),
            .lcout(\U409_CIA.g0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_8_LC_1_7_5 .C_ON=1'b0;
    defparam \U409_CIA.g0_8_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_8_LC_1_7_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_CIA.g0_8_LC_1_7_5  (
            .in0(N__2525),
            .in1(N__2849),
            .in2(_gnd_net_),
            .in3(N__4468),
            .lcout(\U409_CIA.g0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_2_LC_1_15_0 .C_ON=1'b0;
    defparam \U409_CIA.g0_2_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_2_LC_1_15_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_CIA.g0_2_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__2684),
            .in2(_gnd_net_),
            .in3(N__2792),
            .lcout(),
            .ltout(\U409_CIA.g0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_13_LC_1_15_1 .C_ON=1'b0;
    defparam \U409_CIA.g0_13_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_13_LC_1_15_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_CIA.g0_13_LC_1_15_1  (
            .in0(N__2765),
            .in1(N__2816),
            .in2(N__2507),
            .in3(N__2738),
            .lcout(\U409_CIA.g0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_16_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_16_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_16_2  (
            .in0(N__2764),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2784),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_16_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_16_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_16_3  (
            .in0(N__2842),
            .in1(N__2809),
            .in2(N__2852),
            .in3(N__2627),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_1_16_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_1_16_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_1_16_5  (
            .in0(N__2841),
            .in1(N__2808),
            .in2(N__2788),
            .in3(N__2763),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_10_LC_1_17_3 .C_ON=1'b0;
    defparam \U409_CIA.g0_10_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_10_LC_1_17_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_CIA.g0_10_LC_1_17_3  (
            .in0(N__2708),
            .in1(N__6152),
            .in2(N__2654),
            .in3(N__2729),
            .lcout(\U409_CIA.g0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_1_17_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_1_17_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_1_17_5  (
            .in0(N__2706),
            .in1(N__2727),
            .in2(N__2653),
            .in3(N__2676),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_6  (
            .in0(N__2728),
            .in1(N__2707),
            .in2(N__2683),
            .in3(N__2649),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_14_LC_2_7_5 .C_ON=1'b0;
    defparam \U409_CIA.g0_14_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_14_LC_2_7_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.g0_14_LC_2_7_5  (
            .in0(N__2890),
            .in1(N__2621),
            .in2(N__2615),
            .in3(N__2585),
            .lcout(\U409_CIA.g0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_LC_3_16_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_LC_3_16_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_LC_3_16_3  (
            .in0(N__2579),
            .in1(N__2933),
            .in2(_gnd_net_),
            .in3(N__2567),
            .lcout(AUTOVECTORm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.HIROM_0_LC_5_11_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.HIROM_0_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.HIROM_0_LC_5_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.HIROM_0_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__4282),
            .in2(_gnd_net_),
            .in3(N__3013),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEm_3 ),
            .ltout(\U409_ADDRESS_DECODE.CIA_SPACEm_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_0_LC_5_11_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_0_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_0_LC_5_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_0_LC_5_11_2  (
            .in0(N__4459),
            .in1(N__4366),
            .in2(N__2558),
            .in3(N__3037),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_1_0_LC_5_12_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_1_0_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_1_0_LC_5_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_1_0_LC_5_12_4  (
            .in0(N__4365),
            .in1(N__2999),
            .in2(N__4292),
            .in3(N__3043),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACE_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_5_12_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_5_12_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_5_12_7  (
            .in0(N__4458),
            .in1(N__4281),
            .in2(N__3047),
            .in3(N__3000),
            .lcout(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_5_16_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_5_16_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_5_16_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_5_16_4  (
            .in0(N__2978),
            .in1(N__2969),
            .in2(N__6151),
            .in3(N__2951),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_17_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_17_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_17_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_17_4  (
            .in0(N__2924),
            .in1(N__4457),
            .in2(N__5658),
            .in3(N__6147),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.CIA_SPACEm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_5_17_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_5_17_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_5_17_5  (
            .in0(N__5644),
            .in1(N__4367),
            .in2(N__2912),
            .in3(N__3636),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.HIROM_LC_6_11_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_6_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.HIROM_LC_6_11_3  (
            .in0(N__2897),
            .in1(N__4371),
            .in2(N__4460),
            .in3(N__2891),
            .lcout(\U409_ADDRESS_DECODE.HIROMZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_8_5_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_8_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__3312),
            .in2(N__3299),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_5_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_8_5_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_8_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_8_5_1  (
            .in0(_gnd_net_),
            .in1(N__3154),
            .in2(_gnd_net_),
            .in3(N__2855),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__5127),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_8_5_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_8_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(N__3085),
            .in2(_gnd_net_),
            .in3(N__3074),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__5127),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_8_5_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_8_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(N__3118),
            .in2(_gnd_net_),
            .in3(N__3071),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__5127),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_8_5_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_8_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_8_5_4  (
            .in0(_gnd_net_),
            .in1(N__3097),
            .in2(_gnd_net_),
            .in3(N__3068),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_8_5_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_8_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(N__3250),
            .in2(_gnd_net_),
            .in3(N__3065),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_8_5_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_8_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_8_5_6  (
            .in0(_gnd_net_),
            .in1(N__3130),
            .in2(_gnd_net_),
            .in3(N__3062),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__5127),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_8_5_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_8_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_8_5_7  (
            .in0(_gnd_net_),
            .in1(N__3142),
            .in2(_gnd_net_),
            .in3(N__3059),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__5127),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_8_6_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_8_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__3211),
            .in2(_gnd_net_),
            .in3(N__3056),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_8_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_8_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__3340),
            .in2(_gnd_net_),
            .in3(N__3053),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__5129),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_8_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_8_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(N__3407),
            .in2(_gnd_net_),
            .in3(N__3050),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_8_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_8_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__3358),
            .in2(_gnd_net_),
            .in3(N__3182),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__5129),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_8_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_8_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__3193),
            .in2(_gnd_net_),
            .in3(N__3179),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_8_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_8_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(N__3268),
            .in2(_gnd_net_),
            .in3(N__3176),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_8_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_8_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(N__3229),
            .in2(_gnd_net_),
            .in3(N__3173),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_8_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_8_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(N__3167),
            .in2(_gnd_net_),
            .in3(N__3170),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5129),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_9_5_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_9_5_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_9_5_0  (
            .in0(N__3166),
            .in1(N__3155),
            .in2(N__3319),
            .in3(N__3143),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_9_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_9_5_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_9_5_1  (
            .in0(N__3230),
            .in1(N__3131),
            .in2(N__3272),
            .in3(N__3119),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_9_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_9_5_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_9_5_2  (
            .in0(N__3501),
            .in1(N__3529),
            .in2(N__3107),
            .in3(N__3104),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_9_5_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_9_5_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_9_5_3  (
            .in0(N__3098),
            .in1(N__3086),
            .in2(_gnd_net_),
            .in3(N__3296),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_9_5_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_9_5_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_9_5_4  (
            .in0(N__3365),
            .in1(N__3359),
            .in2(N__3347),
            .in3(N__3344),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_9_5_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_9_5_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_9_5_5  (
            .in0(N__3449),
            .in1(N__3500),
            .in2(N__3329),
            .in3(N__3326),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_9_5_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_9_5_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_9_5_6  (
            .in0(N__3297),
            .in1(_gnd_net_),
            .in2(N__3320),
            .in3(_gnd_net_),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_9_5_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_9_5_7 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_9_5_7  (
            .in0(N__3448),
            .in1(N__3298),
            .in2(N__3544),
            .in3(N__3502),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_9_6_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_9_6_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_9_6_0  (
            .in0(N__3546),
            .in1(N__3497),
            .in2(N__3465),
            .in3(N__3278),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5128),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_9_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_9_6_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_9_6_1  (
            .in0(N__3406),
            .in1(N__3212),
            .in2(N__3257),
            .in3(N__3194),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_9_6_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_9_6_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_9_6_2  (
            .in0(N__3547),
            .in1(N__3460),
            .in2(N__3239),
            .in3(N__3236),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5128),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_9_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_9_6_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_9_6_4  (
            .in0(N__3548),
            .in1(N__3498),
            .in2(N__3466),
            .in3(N__3218),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5128),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_9_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_9_6_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_9_6_6  (
            .in0(N__3545),
            .in1(N__3496),
            .in2(N__3464),
            .in3(N__3200),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5128),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_10_5_3 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_10_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_10_5_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK50_LC_10_5_3  (
            .in0(N__3450),
            .in1(N__3559),
            .in2(N__3506),
            .in3(N__3543),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_10_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_10_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_10_6_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_10_6_4  (
            .in0(N__3542),
            .in1(N__3499),
            .in2(N__3467),
            .in3(N__3416),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5125),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_7_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_7_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_7_6 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_7_6  (
            .in0(N__3747),
            .in1(N__3392),
            .in2(N__3698),
            .in3(N__3780),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__5947));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_7_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_7_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_7_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_7_7  (
            .in0(N__3391),
            .in1(N__3748),
            .in2(_gnd_net_),
            .in3(N__3693),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__5947));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_8_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_8_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_8_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_8_2  (
            .in0(N__3863),
            .in1(N__3827),
            .in2(_gnd_net_),
            .in3(N__3688),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__5948));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_8_3 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_8_3 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(N__3373),
            .in2(N__3697),
            .in3(N__3802),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__5948));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_8_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_8_4 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_8_4  (
            .in0(N__3801),
            .in1(N__3847),
            .in2(N__3377),
            .in3(N__3692),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__5948));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_9_5  (
            .in0(N__3919),
            .in1(N__3943),
            .in2(N__3983),
            .in3(N__3826),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_9_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__3781),
            .in2(N__3380),
            .in3(N__3749),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_10_12_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_10_12_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_10_12_0  (
            .in0(N__5675),
            .in1(N__3637),
            .in2(_gnd_net_),
            .in3(N__4385),
            .lcout(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_10_17_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_10_17_3 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_10_17_3  (
            .in0(N__3644),
            .in1(N__5674),
            .in2(_gnd_net_),
            .in3(N__4392),
            .lcout(U409_ADDRESS_DECODE_un1_nREGSPACE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_11_5_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_11_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_11_5_0  (
            .in0(_gnd_net_),
            .in1(N__4542),
            .in2(N__4739),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_11_5_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_11_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__4558),
            .in2(_gnd_net_),
            .in3(N__3590),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__5120),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_11_5_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_11_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(N__4693),
            .in2(_gnd_net_),
            .in3(N__3587),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__5120),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_11_5_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_11_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__4750),
            .in2(_gnd_net_),
            .in3(N__3584),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_11_5_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_11_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_11_5_4  (
            .in0(_gnd_net_),
            .in1(N__4762),
            .in2(_gnd_net_),
            .in3(N__3581),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__5120),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_11_5_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_11_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_11_5_5  (
            .in0(_gnd_net_),
            .in1(N__4504),
            .in2(_gnd_net_),
            .in3(N__3578),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_11_5_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_11_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_11_5_6  (
            .in0(_gnd_net_),
            .in1(N__4810),
            .in2(_gnd_net_),
            .in3(N__3575),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__5120),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_11_5_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_11_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_11_5_7  (
            .in0(_gnd_net_),
            .in1(N__5146),
            .in2(_gnd_net_),
            .in3(N__3671),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_11_6_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_11_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__4774),
            .in2(_gnd_net_),
            .in3(N__3668),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_11_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_11_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__4828),
            .in2(_gnd_net_),
            .in3(N__3665),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__5123),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_11_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_11_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__4708),
            .in2(_gnd_net_),
            .in3(N__3662),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__5123),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_11_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_11_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__4570),
            .in2(_gnd_net_),
            .in3(N__3659),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__5123),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_11_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_11_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(N__4840),
            .in2(_gnd_net_),
            .in3(N__3656),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__5123),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_11_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_11_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__4672),
            .in2(_gnd_net_),
            .in3(N__3653),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_11_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_11_6_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4799),
            .in3(N__3650),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_11_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_11_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(N__4529),
            .in2(_gnd_net_),
            .in3(N__3647),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5123),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.LOWROM_LC_11_7_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.LOWROM_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.LOWROM_LC_11_7_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_ADDRESS_DECODE.LOWROM_LC_11_7_0  (
            .in0(N__4301),
            .in1(N__4394),
            .in2(N__5600),
            .in3(N__4472),
            .lcout(\U409_ADDRESS_DECODE.LOWROMZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_11_7_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_11_7_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_11_7_2  (
            .in0(N__5273),
            .in1(N__5195),
            .in2(N__3872),
            .in3(N__5236),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5126),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_7_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_7_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_7_6  (
            .in0(N__3982),
            .in1(N__3920),
            .in2(_gnd_net_),
            .in3(N__3944),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_11_7_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_11_7_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_11_7_7  (
            .in0(N__3746),
            .in1(N__3824),
            .in2(N__3782),
            .in3(N__3843),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_11_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_11_8_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_11_8_0  (
            .in0(N__3797),
            .in1(N__3969),
            .in2(N__3713),
            .in3(N__3854),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_8_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_8_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__3940),
            .in2(_gnd_net_),
            .in3(N__3917),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_11_8_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_11_8_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_11_8_2  (
            .in0(N__3848),
            .in1(N__3825),
            .in2(N__3803),
            .in3(N__3968),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_11_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_11_8_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_11_8_3  (
            .in0(N__3776),
            .in1(N__3745),
            .in2(N__3716),
            .in3(N__3709),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_8_4 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_8_4  (
            .in0(N__4151),
            .in1(N__4110),
            .in2(N__3701),
            .in3(N__3891),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_8_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_8_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_8_5 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_8_5  (
            .in0(N__3971),
            .in1(_gnd_net_),
            .in2(N__3986),
            .in3(N__3941),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__5943));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_8_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_8_6 .LUT_INIT=16'b0001000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_8_6  (
            .in0(N__4150),
            .in1(N__3970),
            .in2(N__4114),
            .in3(N__3892),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__5943));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_8_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_8_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_8_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_8_7  (
            .in0(N__3972),
            .in1(N__3918),
            .in2(_gnd_net_),
            .in3(N__3942),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__5943));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_9_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_9_4 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_9_4  (
            .in0(N__4867),
            .in1(N__3899),
            .in2(_gnd_net_),
            .in3(N__3893),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .ce(),
            .sr(N__5936));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_11_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_11_10_0 .LUT_INIT=16'b1111011100000111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_11_10_0  (
            .in0(N__4903),
            .in1(N__4923),
            .in2(N__4976),
            .in3(N__4480),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.m9_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_10_1 .LUT_INIT=16'b0000001010001010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_10_1  (
            .in0(N__6106),
            .in1(N__4954),
            .in2(N__3878),
            .in3(N__4487),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_11_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_11_10_2 .LUT_INIT=16'b0000001001010111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_11_10_2  (
            .in0(N__4952),
            .in1(N__4924),
            .in2(N__4907),
            .in3(N__4481),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_10_3 .LUT_INIT=16'b0010101000001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_10_3  (
            .in0(N__6107),
            .in1(N__4974),
            .in2(N__3875),
            .in3(N__4953),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_11_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_11_10_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_11_10_4  (
            .in0(N__4951),
            .in1(N__4877),
            .in2(N__4105),
            .in3(N__4891),
            .lcout(\U409_TRANSFER_ACK.N_105 ),
            .ltout(\U409_TRANSFER_ACK.N_105_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_11_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_11_10_5 .LUT_INIT=16'b0000001101000111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_11_10_5  (
            .in0(N__4922),
            .in1(N__4973),
            .in2(N__4490),
            .in3(N__4902),
            .lcout(\U409_TRANSFER_ACK.m9_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__4876),
            .in2(_gnd_net_),
            .in3(N__4890),
            .lcout(\U409_TRANSFER_ACK.N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_11_10_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_11_10_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_11_10_7  (
            .in0(N__4464),
            .in1(N__4393),
            .in2(_gnd_net_),
            .in3(N__4300),
            .lcout(\U409_ADDRESS_DECODE.un5_nRAMSPACEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_LC_11_11_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_LC_11_11_0 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_LC_11_11_0  (
            .in0(N__5683),
            .in1(N__4228),
            .in2(N__4214),
            .in3(N__6108),
            .lcout(ROMENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_11_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_11_12_2 .LUT_INIT=16'b0111011101111111;
    LogicCell40 \U409_ADDRESS_DECODE.ROMENm_i_LC_11_12_2  (
            .in0(N__6109),
            .in1(N__5676),
            .in2(N__4232),
            .in3(N__4213),
            .lcout(ROMENm_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_11_13_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_11_13_0 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_11_13_0  (
            .in0(N__4166),
            .in1(N__4138),
            .in2(N__4106),
            .in3(N__4049),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_12_4_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_12_4_4 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_12_4_4  (
            .in0(N__4025),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4660),
            .lcout(U409_ADDRESS_DECODE_un1_nCIACS0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_12_4_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_12_4_6 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_12_4_6  (
            .in0(_gnd_net_),
            .in1(N__4646),
            .in2(_gnd_net_),
            .in3(N__4661),
            .lcout(U409_ADDRESS_DECODE_un1_nCIACS1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_12_4_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_12_4_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_12_4_7 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_12_4_7  (
            .in0(N__5711),
            .in1(N__5673),
            .in2(_gnd_net_),
            .in3(N__5589),
            .lcout(U409_ADDRESS_DECODE_un1_nRAMSPACE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_12_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_12_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_12_5_2  (
            .in0(N__4546),
            .in1(N__4738),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5119),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_12_5_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_12_5_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_12_5_4  (
            .in0(N__5233),
            .in1(N__5266),
            .in2(N__5202),
            .in3(N__4601),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5119),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_12_5_5 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_12_5_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \U409_TICK.TICK60_LC_12_5_5  (
            .in0(N__5265),
            .in1(N__5235),
            .in2(N__5204),
            .in3(N__4582),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5119),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_12_5_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_12_5_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_12_5_6  (
            .in0(N__4571),
            .in1(N__4559),
            .in2(N__4547),
            .in3(N__4528),
            .lcout(\U409_TICK.TICK603_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_12_5_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_12_5_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_12_5_7  (
            .in0(N__5264),
            .in1(N__5234),
            .in2(N__4517),
            .in3(N__5192),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5119),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_12_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_12_6_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_12_6_1  (
            .in0(N__5147),
            .in1(N__4775),
            .in2(N__4508),
            .in3(N__4673),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_12_6_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_12_6_2 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_12_6_2  (
            .in0(N__4737),
            .in1(N__5232),
            .in2(N__4493),
            .in3(N__5269),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5121),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_12_6_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_12_6_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_12_6_3  (
            .in0(N__4841),
            .in1(N__4829),
            .in2(N__4817),
            .in3(N__4798),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(\U409_TICK.TICK603_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_12_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_12_6_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_12_6_4  (
            .in0(N__5193),
            .in1(N__5268),
            .in2(N__4784),
            .in3(N__4781),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5121),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_12_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_12_6_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_12_6_5  (
            .in0(N__4763),
            .in1(N__4751),
            .in2(_gnd_net_),
            .in3(N__4736),
            .lcout(),
            .ltout(\U409_TICK.TICK603_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_12_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_12_6_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_12_6_6  (
            .in0(N__4715),
            .in1(N__4709),
            .in2(N__4697),
            .in3(N__4694),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_12_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_12_6_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_12_6_7  (
            .in0(N__5231),
            .in1(N__5194),
            .in2(N__4682),
            .in3(N__4679),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5121),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_12_7_1 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_12_7_1 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_12_7_1  (
            .in0(N__4990),
            .in1(N__5071),
            .in2(N__5054),
            .in3(N__5029),
            .lcout(CIA_ENABLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_HOLD_LC_12_7_2 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_LC_12_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_HOLD_LC_12_7_2 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U409_CIA.CIA_HOLD_LC_12_7_2  (
            .in0(N__5070),
            .in1(N__5049),
            .in2(N__5030),
            .in3(N__4989),
            .lcout(\U409_CIA.CIA_HOLDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5387),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_12_8_4 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_12_8_4 .LUT_INIT=16'b0100010000100010;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_12_8_4  (
            .in0(N__5866),
            .in1(N__5482),
            .in2(_gnd_net_),
            .in3(N__5444),
            .lcout(),
            .ltout(\U409_CIA.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_12_8_5 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_12_8_5 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \U409_CIA.VMA_LC_12_8_5  (
            .in0(N__5048),
            .in1(N__5867),
            .in2(N__4649),
            .in3(N__5762),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5385),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_9_5 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_9_5  (
            .in0(N__5078),
            .in1(N__5053),
            .in2(N__5025),
            .in3(N__4994),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__5742));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_12_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_12_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5410),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__5749));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_12_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_12_10_4 .LUT_INIT=16'b0100011101000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_12_10_4  (
            .in0(N__4975),
            .in1(N__4955),
            .in2(N__4934),
            .in3(N__4853),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__5749));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4925),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__5749));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_12_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_12_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_12_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4892),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__5749));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_12_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_12_11_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(N__4868),
            .in2(_gnd_net_),
            .in3(N__4852),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_12_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_12_0 .LUT_INIT=16'b0101010110100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_12_0  (
            .in0(N__5348),
            .in1(_gnd_net_),
            .in2(N__5306),
            .in3(N__5327),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__5750));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_12_1 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_12_1  (
            .in0(N__5325),
            .in1(N__5304),
            .in2(N__5368),
            .in3(N__5346),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__5750));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_12_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_12_12_3 .LUT_INIT=16'b1111101100101010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_12_12_3  (
            .in0(N__5279),
            .in1(N__5354),
            .in2(N__5369),
            .in3(N__5528),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__5750));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_12_5 .LUT_INIT=16'b0001000111001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_12_5  (
            .in0(N__5326),
            .in1(N__5300),
            .in2(_gnd_net_),
            .in3(N__5347),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__5750));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_13_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_13_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_13_0  (
            .in0(N__5323),
            .in1(N__5344),
            .in2(_gnd_net_),
            .in3(N__5296),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_1_LC_12_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_1_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_1_LC_12_13_5 .LUT_INIT=16'b0000100000001000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_1_LC_12_13_5  (
            .in0(N__5345),
            .in1(N__5324),
            .in2(N__5305),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_13_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_13_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_13_5_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_13_5_2  (
            .in0(N__5267),
            .in1(N__5237),
            .in2(N__5203),
            .in3(N__5156),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5118),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_13_7_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_13_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__5439),
            .in2(N__5483),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_13_7_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_13_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__5780),
            .in2(_gnd_net_),
            .in3(N__5087),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__5386),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_13_7_2 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_13_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__5861),
            .in2(_gnd_net_),
            .in3(N__5084),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_13_7_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_13_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__5803),
            .in2(_gnd_net_),
            .in3(N__5081),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__5386),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_13_7_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_13_7_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(N__5829),
            .in2(_gnd_net_),
            .in3(N__5507),
            .lcout(),
            .ltout(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_13_7_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_13_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_13_7_5 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_13_7_5  (
            .in0(N__5862),
            .in1(N__5501),
            .in2(N__5504),
            .in3(N__5477),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5386),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_13_7_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_13_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_13_7_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_13_7_6  (
            .in0(N__5476),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5386),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_13_7_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_13_7_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_13_7_7  (
            .in0(N__5440),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5478),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5386),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_13_8_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_13_8_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_13_8_0  (
            .in0(N__5442),
            .in1(N__5782),
            .in2(N__5831),
            .in3(N__5804),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_13_8_1 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_13_8_1 .LUT_INIT=16'b0010011001100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_13_8_1  (
            .in0(N__5865),
            .in1(N__5495),
            .in2(N__5489),
            .in3(N__5481),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5384),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_2_LC_13_8_3 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_13_8_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_CIA.CLKCIA_RNO_2_LC_13_8_3  (
            .in0(N__5863),
            .in1(N__5479),
            .in2(_gnd_net_),
            .in3(N__5441),
            .lcout(),
            .ltout(\U409_CIA.N_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_0_LC_13_8_4 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_13_8_4 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \U409_CIA.CLKCIA_RNO_0_LC_13_8_4  (
            .in0(_gnd_net_),
            .in1(N__5403),
            .in2(N__5486),
            .in3(N__5761),
            .lcout(),
            .ltout(\U409_CIA.CLKCIAZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_LC_13_8_5 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLKCIA_LC_13_8_5 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \U409_CIA.CLKCIA_LC_13_8_5  (
            .in0(N__5837),
            .in1(N__5480),
            .in2(N__5447),
            .in3(N__5443),
            .lcout(CLKCIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5384),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_1_LC_13_8_6 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_13_8_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CLKCIA_RNO_1_LC_13_8_6  (
            .in0(N__5802),
            .in1(N__5783),
            .in2(N__5830),
            .in3(N__5864),
            .lcout(\U409_CIA.CLKCIA6_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_13_8_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_13_8_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_13_8_7  (
            .in0(N__5822),
            .in1(N__5801),
            .in2(_gnd_net_),
            .in3(N__5781),
            .lcout(\U409_CIA.CLKCIA8_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_13_9_2.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_13_9_2.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_13_9_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_13_9_2 (
            .in0(N__6089),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_13_11_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_13_11_1 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_13_11_1  (
            .in0(N__5723),
            .in1(N__5710),
            .in2(N__5687),
            .in3(N__5593),
            .lcout(nBUFEN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_13_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_13_12_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_13_12_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_13_12_0  (
            .in0(N__6185),
            .in1(_gnd_net_),
            .in2(N__6125),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_13_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_13_12_1 .LUT_INIT=16'b0000101011101010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_13_12_1  (
            .in0(N__5539),
            .in1(N__6199),
            .in2(N__6126),
            .in3(N__6173),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_13_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_13_12_2 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_13_12_2  (
            .in0(N__6183),
            .in1(N__5527),
            .in2(N__6200),
            .in3(N__5516),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_13_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_13_12_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_13_12_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5510),
            .in3(N__6112),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_13_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_13_12_5 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_13_12_5  (
            .in0(N__6116),
            .in1(N__6198),
            .in2(_gnd_net_),
            .in3(N__6184),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_14_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_14_12_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_14_12_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_LC_14_12_0  (
            .in0(N__6110),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6172),
            .lcout(TACK_EN_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .ce(N__6161),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_15_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_15_11_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_15_11_6  (
            .in0(N__6111),
            .in1(N__5983),
            .in2(_gnd_net_),
            .in3(N__5969),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_iobuf_RNO_LC_19_18_0.C_ON=1'b0;
    defparam TACKn_iobuf_RNO_LC_19_18_0.SEQ_MODE=4'b0000;
    defparam TACKn_iobuf_RNO_LC_19_18_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 TACKn_iobuf_RNO_LC_19_18_0 (
            .in0(N__5900),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_365_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 18 2024 19:21:53

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RAMENn : out std_logic;
    RASn : out std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__10191\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_OUT_i_i\ : std_logic;
signal \bfn_6_8_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \N_71_cascade_\ : std_logic;
signal \N_736_i\ : std_logic;
signal \U712_REG_SM.UDS_OUT_2_0_a2_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_82\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUUBEn_iZ0Z_0\ : std_logic;
signal \N_55_i\ : std_logic;
signal \U712_BYTE_ENABLE.LLBE_0_cascade_\ : std_logic;
signal \CLLBEn_c\ : std_logic;
signal \A_c_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \U712_BYTE_ENABLE.N_79_cascade_\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_iZ0Z_0_cascade_\ : std_logic;
signal \N_54_i\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_REG_SM.N_163_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_178_cascade_\ : std_logic;
signal \U712_REG_SM.N_163_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_45_0_0_en_cascade_\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \U712_CYCLE_TERM.N_45_0_0_en_0\ : std_logic;
signal \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1\ : std_logic;
signal \U712_BYTE_ENABLE.LMBE_0\ : std_logic;
signal \CLMBEn_c\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_175_cascade_\ : std_logic;
signal \U712_REG_SM.N_175_0_0\ : std_logic;
signal \U712_REG_SM.DS_EN_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_REG_SM.N_175\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.N_156_0\ : std_logic;
signal \U712_REG_SM.N_156_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_166_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_1\ : std_logic;
signal \U712_REG_SM.N_148_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_164_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_181\ : std_logic;
signal \U712_REG_SM.DS_EN_7_0_cascade_\ : std_logic;
signal \C1_c\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.LDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_LDSn_i\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\ : std_logic;
signal \A_c_10\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_\ : std_logic;
signal \A_c_12\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_CHIP_RAM.N_61_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_101_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_a2_0_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_68_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_108\ : std_logic;
signal \U712_CHIP_RAM.N_109\ : std_logic;
signal \U712_CHIP_RAM.N_108_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0\ : std_logic;
signal \U712_CHIP_RAM.N_65_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_114\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_0_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\ : std_logic;
signal \U712_REG_SM.N_148_0\ : std_logic;
signal \U712_REG_SM.N_151_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_160_0\ : std_logic;
signal \U712_REG_SM.N_147_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_161_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_161_0_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \U712_REG_SM.N_187_cascade_\ : std_logic;
signal \U712_REG_SM.N_183\ : std_logic;
signal \U712_REG_SM.N_147_0\ : std_logic;
signal \U712_REG_SM.N_153_0\ : std_logic;
signal \U712_REG_SM.N_174\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \CLK40_OUT_i_i\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_187\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.DS_ENZ0\ : std_logic;
signal \U712_REG_SM.UDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_UDSn_i\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \DRDDIR_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_32\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.N_34\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_58_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_97_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \U712_CHIP_RAM.N_421_tz\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_68\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_52_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_61\ : std_logic;
signal \U712_CHIP_RAM.N_90_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_69\ : std_logic;
signal \U712_CHIP_RAM.N_57\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_7\ : std_logic;
signal \U712_REG_SM.N_151_0\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_1\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_0\ : std_logic;
signal \U712_REG_SM.N_159_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_165\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_REG_SM.C1_SYNC_RNIPBP14Z0Z_2\ : std_logic;
signal \U712_REG_SM.N_180_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.N_31\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_4_cascade_\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.N_35\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.un6_CPU_CYCLE_START\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_52\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER35\ : std_logic;
signal \U712_CHIP_RAM.N_46_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_116\ : std_logic;
signal \U712_CHIP_RAM.N_116_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER39\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_46\ : std_logic;
signal \U712_CHIP_RAM.N_96\ : std_logic;
signal \U712_CHIP_RAM.N_124\ : std_logic;
signal \U712_CHIP_RAM.N_96_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_72\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_65\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_5\ : std_logic;
signal \U712_REG_SM.N_159_0\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \CLK40_OUT_i\ : std_logic;
signal \U712_CYCLE_TERM.N_49_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_5_cascade_\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_36\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.N_33\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_6_cascade_\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.N_37\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_7\ : std_logic;
signal \U712_CHIP_RAM.N_38\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\ : std_logic;
signal \CASn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    CLK_EN <= \CLK_EN_wire\;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    LDSn <= \LDSn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_OUT_i\,
            REFERENCECLK => \N__3644\,
            RESETB => \N__6770\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_OUT\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10191\,
            DIN => \N__10190\,
            DOUT => \N__10189\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10191\,
            PADOUT => \N__10190\,
            PADIN => \N__10189\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4127\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10182\,
            DIN => \N__10181\,
            DOUT => \N__10180\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10182\,
            PADOUT => \N__10181\,
            PADIN => \N__10180\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10173\,
            DIN => \N__10172\,
            DOUT => \N__10171\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10173\,
            PADOUT => \N__10172\,
            PADIN => \N__10171\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8876\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10164\,
            DIN => \N__10163\,
            DOUT => \N__10162\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10164\,
            PADOUT => \N__10163\,
            PADIN => \N__10162\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5009\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10155\,
            DIN => \N__10154\,
            DOUT => \N__10153\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10155\,
            PADOUT => \N__10154\,
            PADIN => \N__10153\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10146\,
            DIN => \N__10145\,
            DOUT => \N__10144\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10146\,
            PADOUT => \N__10145\,
            PADIN => \N__10144\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10137\,
            DIN => \N__10136\,
            DOUT => \N__10135\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10137\,
            PADOUT => \N__10136\,
            PADIN => \N__10135\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10128\,
            DIN => \N__10127\,
            DOUT => \N__10126\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10128\,
            PADOUT => \N__10127\,
            PADIN => \N__10126\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10119\,
            DIN => \N__10118\,
            DOUT => \N__10117\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10119\,
            PADOUT => \N__10118\,
            PADIN => \N__10117\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10110\,
            DIN => \N__10109\,
            DOUT => \N__10108\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10110\,
            PADOUT => \N__10109\,
            PADIN => \N__10108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10101\,
            DIN => \N__10100\,
            DOUT => \N__10099\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10101\,
            PADOUT => \N__10100\,
            PADIN => \N__10099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8075\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10092\,
            DIN => \N__10091\,
            DOUT => \N__10090\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10092\,
            PADOUT => \N__10091\,
            PADIN => \N__10090\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5359\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10083\,
            DIN => \N__10082\,
            DOUT => \N__10081\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10083\,
            PADOUT => \N__10082\,
            PADIN => \N__10081\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10074\,
            DIN => \N__10073\,
            DOUT => \N__10072\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10074\,
            PADOUT => \N__10073\,
            PADIN => \N__10072\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10065\,
            DIN => \N__10064\,
            DOUT => \N__10063\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10065\,
            PADOUT => \N__10064\,
            PADIN => \N__10063\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4142\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10056\,
            DIN => \N__10055\,
            DOUT => \N__10054\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10056\,
            PADOUT => \N__10055\,
            PADIN => \N__10054\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10047\,
            DIN => \N__10046\,
            DOUT => \N__10045\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10047\,
            PADOUT => \N__10046\,
            PADIN => \N__10045\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10038\,
            DIN => \N__10037\,
            DOUT => \N__10036\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10038\,
            PADOUT => \N__10037\,
            PADIN => \N__10036\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5969\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10029\,
            DIN => \N__10028\,
            DOUT => \N__10027\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10029\,
            PADOUT => \N__10028\,
            PADIN => \N__10027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10020\,
            DIN => \N__10019\,
            DOUT => \N__10018\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10020\,
            PADOUT => \N__10019\,
            PADIN => \N__10018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8771\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10011\,
            DIN => \N__10010\,
            DOUT => \N__10009\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10011\,
            PADOUT => \N__10010\,
            PADIN => \N__10009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10002\,
            DIN => \N__10001\,
            DOUT => \N__10000\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10002\,
            PADOUT => \N__10001\,
            PADIN => \N__10000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9993\,
            DIN => \N__9992\,
            DOUT => \N__9991\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9993\,
            PADOUT => \N__9992\,
            PADIN => \N__9991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9984\,
            DIN => \N__9983\,
            DOUT => \N__9982\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9984\,
            PADOUT => \N__9983\,
            PADIN => \N__9982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9975\,
            DIN => \N__9974\,
            DOUT => \N__9973\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9975\,
            PADOUT => \N__9974\,
            PADIN => \N__9973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9966\,
            DIN => \N__9965\,
            DOUT => \N__9964\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9966\,
            PADOUT => \N__9965\,
            PADIN => \N__9964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5630\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9957\,
            DIN => \N__9956\,
            DOUT => \N__9955\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9957\,
            PADOUT => \N__9956\,
            PADIN => \N__9955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9948\,
            DIN => \N__9947\,
            DOUT => \N__9946\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9948\,
            PADOUT => \N__9947\,
            PADIN => \N__9946\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9939\,
            DIN => \N__9938\,
            DOUT => \N__9937\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9939\,
            PADOUT => \N__9938\,
            PADIN => \N__9937\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9930\,
            DIN => \N__9929\,
            DOUT => \N__9928\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9930\,
            PADOUT => \N__9929\,
            PADIN => \N__9928\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9921\,
            DIN => \N__9920\,
            DOUT => \N__9919\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9921\,
            PADOUT => \N__9920\,
            PADIN => \N__9919\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9912\,
            DIN => \N__9911\,
            DOUT => \N__9910\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9912\,
            PADOUT => \N__9911\,
            PADIN => \N__9910\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7595\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9903\,
            DIN => \N__9902\,
            DOUT => \N__9901\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9903\,
            PADOUT => \N__9902\,
            PADIN => \N__9901\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9894\,
            DIN => \N__9893\,
            DOUT => \N__9892\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9894\,
            PADOUT => \N__9893\,
            PADIN => \N__9892\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9885\,
            DIN => \N__9884\,
            DOUT => \N__9883\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9885\,
            PADOUT => \N__9884\,
            PADIN => \N__9883\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9876\,
            DIN => \N__9875\,
            DOUT => \N__9874\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9876\,
            PADOUT => \N__9875\,
            PADIN => \N__9874\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9867\,
            DIN => \N__9866\,
            DOUT => \N__9865\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9867\,
            PADOUT => \N__9866\,
            PADIN => \N__9865\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4796\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9858\,
            DIN => \N__9857\,
            DOUT => \N__9856\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9858\,
            PADOUT => \N__9857\,
            PADIN => \N__9856\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4448\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9849\,
            DIN => \N__9848\,
            DOUT => \N__9847\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9849\,
            PADOUT => \N__9848\,
            PADIN => \N__9847\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9840\,
            DIN => \N__9839\,
            DOUT => \N__9838\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9840\,
            PADOUT => \N__9839\,
            PADIN => \N__9838\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8843\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9831\,
            DIN => \N__9830\,
            DOUT => \N__9829\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9831\,
            PADOUT => \N__9830\,
            PADIN => \N__9829\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9822\,
            DIN => \N__9821\,
            DOUT => \N__9820\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9822\,
            PADOUT => \N__9821\,
            PADIN => \N__9820\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9813\,
            DIN => \N__9812\,
            DOUT => \N__9811\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9813\,
            PADOUT => \N__9812\,
            PADIN => \N__9811\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3665\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9804\,
            DIN => \N__9803\,
            DOUT => \N__9802\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9804\,
            PADOUT => \N__9803\,
            PADIN => \N__9802\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9795\,
            DIN => \N__9794\,
            DOUT => \N__9793\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9795\,
            PADOUT => \N__9794\,
            PADIN => \N__9793\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5147\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9786\,
            DIN => \N__9785\,
            DOUT => \N__9784\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9786\,
            PADOUT => \N__9785\,
            PADIN => \N__9784\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4958\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9777\,
            DIN => \N__9776\,
            DOUT => \N__9775\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9777\,
            PADOUT => \N__9776\,
            PADIN => \N__9775\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9768\,
            DIN => \N__9767\,
            DOUT => \N__9766\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9768\,
            PADOUT => \N__9767\,
            PADIN => \N__9766\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9759\,
            DIN => \N__9758\,
            DOUT => \N__9757\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9759\,
            PADOUT => \N__9758\,
            PADIN => \N__9757\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9750\,
            DIN => \N__9749\,
            DOUT => \N__9748\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9750\,
            PADOUT => \N__9749\,
            PADIN => \N__9748\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7931\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9741\,
            DIN => \N__9740\,
            DOUT => \N__9739\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9741\,
            PADOUT => \N__9740\,
            PADIN => \N__9739\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9732\,
            DIN => \N__9731\,
            DOUT => \N__9730\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9732\,
            PADOUT => \N__9731\,
            PADIN => \N__9730\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5948\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9723\,
            DIN => \N__9722\,
            DOUT => \N__9721\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9723\,
            PADOUT => \N__9722\,
            PADIN => \N__9721\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6791\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9714\,
            DIN => \N__9713\,
            DOUT => \N__9712\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9714\,
            PADOUT => \N__9713\,
            PADIN => \N__9712\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4082\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9705\,
            DIN => \N__9704\,
            DOUT => \N__9703\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9705\,
            PADOUT => \N__9704\,
            PADIN => \N__9703\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8447\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9696\,
            DIN => \N__9695\,
            DOUT => \N__9694\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9696\,
            PADOUT => \N__9695\,
            PADIN => \N__9694\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5143\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9687\,
            DIN => \N__9686\,
            DOUT => \N__9685\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9687\,
            PADOUT => \N__9686\,
            PADIN => \N__9685\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9678\,
            DIN => \N__9677\,
            DOUT => \N__9676\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9678\,
            PADOUT => \N__9677\,
            PADIN => \N__9676\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9669\,
            DIN => \N__9668\,
            DOUT => \N__9667\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9669\,
            PADOUT => \N__9668\,
            PADIN => \N__9667\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4166\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9660\,
            DIN => \N__9659\,
            DOUT => \N__9658\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9660\,
            PADOUT => \N__9659\,
            PADIN => \N__9658\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8864\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9651\,
            DIN => \N__9650\,
            DOUT => \N__9649\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9651\,
            PADOUT => \N__9650\,
            PADIN => \N__9649\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5045\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9642\,
            DIN => \N__9641\,
            DOUT => \N__9640\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9642\,
            PADOUT => \N__9641\,
            PADIN => \N__9640\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3884\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9633\,
            DIN => \N__9632\,
            DOUT => \N__9631\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9633\,
            PADOUT => \N__9632\,
            PADIN => \N__9631\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9624\,
            DIN => \N__9623\,
            DOUT => \N__9622\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9624\,
            PADOUT => \N__9623\,
            PADIN => \N__9622\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9615\,
            DIN => \N__9614\,
            DOUT => \N__9613\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9615\,
            PADOUT => \N__9614\,
            PADIN => \N__9613\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9606\,
            DIN => \N__9605\,
            DOUT => \N__9604\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9606\,
            PADOUT => \N__9605\,
            PADIN => \N__9604\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9597\,
            DIN => \N__9596\,
            DOUT => \N__9595\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9597\,
            PADOUT => \N__9596\,
            PADIN => \N__9595\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4979\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9588\,
            DIN => \N__9587\,
            DOUT => \N__9586\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9588\,
            PADOUT => \N__9587\,
            PADIN => \N__9586\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9579\,
            DIN => \N__9578\,
            DOUT => \N__9577\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9579\,
            PADOUT => \N__9578\,
            PADIN => \N__9577\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3797\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9570\,
            DIN => \N__9569\,
            DOUT => \N__9568\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9570\,
            PADOUT => \N__9569\,
            PADIN => \N__9568\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3836\,
            DIN0 => OPEN,
            DOUT0 => \N__4817\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9561\,
            DIN => \N__9560\,
            DOUT => \N__9559\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9561\,
            PADOUT => \N__9560\,
            PADIN => \N__9559\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6755\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9552\,
            DIN => \N__9551\,
            DOUT => \N__9550\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9552\,
            PADOUT => \N__9551\,
            PADIN => \N__9550\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9543\,
            DIN => \N__9542\,
            DOUT => \N__9541\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9543\,
            PADOUT => \N__9542\,
            PADIN => \N__9541\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9534\,
            DIN => \N__9533\,
            DOUT => \N__9532\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9534\,
            PADOUT => \N__9533\,
            PADIN => \N__9532\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8696\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9525\,
            DIN => \N__9524\,
            DOUT => \N__9523\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9525\,
            PADOUT => \N__9524\,
            PADIN => \N__9523\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9516\,
            DIN => \N__9515\,
            DOUT => \N__9514\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9516\,
            PADOUT => \N__9515\,
            PADIN => \N__9514\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9507\,
            DIN => \N__9506\,
            DOUT => \N__9505\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9507\,
            PADOUT => \N__9506\,
            PADIN => \N__9505\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9498\,
            DIN => \N__9497\,
            DOUT => \N__9496\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9498\,
            PADOUT => \N__9497\,
            PADIN => \N__9496\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9489\,
            DIN => \N__9488\,
            DOUT => \N__9487\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9489\,
            PADOUT => \N__9488\,
            PADIN => \N__9487\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6737\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9480\,
            DIN => \N__9479\,
            DOUT => \N__9478\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9480\,
            PADOUT => \N__9479\,
            PADIN => \N__9478\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5063\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2252\ : InMux
    port map (
            O => \N__9461\,
            I => \N__9446\
        );

    \I__2251\ : InMux
    port map (
            O => \N__9460\,
            I => \N__9443\
        );

    \I__2250\ : InMux
    port map (
            O => \N__9459\,
            I => \N__9440\
        );

    \I__2249\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9437\
        );

    \I__2248\ : InMux
    port map (
            O => \N__9457\,
            I => \N__9434\
        );

    \I__2247\ : InMux
    port map (
            O => \N__9456\,
            I => \N__9431\
        );

    \I__2246\ : InMux
    port map (
            O => \N__9455\,
            I => \N__9428\
        );

    \I__2245\ : InMux
    port map (
            O => \N__9454\,
            I => \N__9425\
        );

    \I__2244\ : InMux
    port map (
            O => \N__9453\,
            I => \N__9418\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9452\,
            I => \N__9418\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9451\,
            I => \N__9418\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9450\,
            I => \N__9415\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9412\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__9446\,
            I => \N__9405\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__9443\,
            I => \N__9399\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__9440\,
            I => \N__9390\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__9437\,
            I => \N__9387\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__9434\,
            I => \N__9381\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__9431\,
            I => \N__9378\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__9428\,
            I => \N__9375\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__9425\,
            I => \N__9371\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9418\,
            I => \N__9362\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__9415\,
            I => \N__9357\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__9412\,
            I => \N__9352\
        );

    \I__2228\ : SRMux
    port map (
            O => \N__9411\,
            I => \N__9275\
        );

    \I__2227\ : SRMux
    port map (
            O => \N__9410\,
            I => \N__9275\
        );

    \I__2226\ : SRMux
    port map (
            O => \N__9409\,
            I => \N__9275\
        );

    \I__2225\ : SRMux
    port map (
            O => \N__9408\,
            I => \N__9275\
        );

    \I__2224\ : Glb2LocalMux
    port map (
            O => \N__9405\,
            I => \N__9275\
        );

    \I__2223\ : SRMux
    port map (
            O => \N__9404\,
            I => \N__9275\
        );

    \I__2222\ : SRMux
    port map (
            O => \N__9403\,
            I => \N__9275\
        );

    \I__2221\ : SRMux
    port map (
            O => \N__9402\,
            I => \N__9275\
        );

    \I__2220\ : Glb2LocalMux
    port map (
            O => \N__9399\,
            I => \N__9275\
        );

    \I__2219\ : SRMux
    port map (
            O => \N__9398\,
            I => \N__9275\
        );

    \I__2218\ : SRMux
    port map (
            O => \N__9397\,
            I => \N__9275\
        );

    \I__2217\ : SRMux
    port map (
            O => \N__9396\,
            I => \N__9275\
        );

    \I__2216\ : SRMux
    port map (
            O => \N__9395\,
            I => \N__9275\
        );

    \I__2215\ : SRMux
    port map (
            O => \N__9394\,
            I => \N__9275\
        );

    \I__2214\ : SRMux
    port map (
            O => \N__9393\,
            I => \N__9275\
        );

    \I__2213\ : Glb2LocalMux
    port map (
            O => \N__9390\,
            I => \N__9275\
        );

    \I__2212\ : Glb2LocalMux
    port map (
            O => \N__9387\,
            I => \N__9275\
        );

    \I__2211\ : SRMux
    port map (
            O => \N__9386\,
            I => \N__9275\
        );

    \I__2210\ : SRMux
    port map (
            O => \N__9385\,
            I => \N__9275\
        );

    \I__2209\ : SRMux
    port map (
            O => \N__9384\,
            I => \N__9275\
        );

    \I__2208\ : Glb2LocalMux
    port map (
            O => \N__9381\,
            I => \N__9275\
        );

    \I__2207\ : Glb2LocalMux
    port map (
            O => \N__9378\,
            I => \N__9275\
        );

    \I__2206\ : Glb2LocalMux
    port map (
            O => \N__9375\,
            I => \N__9275\
        );

    \I__2205\ : SRMux
    port map (
            O => \N__9374\,
            I => \N__9275\
        );

    \I__2204\ : Glb2LocalMux
    port map (
            O => \N__9371\,
            I => \N__9275\
        );

    \I__2203\ : SRMux
    port map (
            O => \N__9370\,
            I => \N__9275\
        );

    \I__2202\ : SRMux
    port map (
            O => \N__9369\,
            I => \N__9275\
        );

    \I__2201\ : SRMux
    port map (
            O => \N__9368\,
            I => \N__9275\
        );

    \I__2200\ : SRMux
    port map (
            O => \N__9367\,
            I => \N__9275\
        );

    \I__2199\ : SRMux
    port map (
            O => \N__9366\,
            I => \N__9275\
        );

    \I__2198\ : SRMux
    port map (
            O => \N__9365\,
            I => \N__9275\
        );

    \I__2197\ : Glb2LocalMux
    port map (
            O => \N__9362\,
            I => \N__9275\
        );

    \I__2196\ : SRMux
    port map (
            O => \N__9361\,
            I => \N__9275\
        );

    \I__2195\ : SRMux
    port map (
            O => \N__9360\,
            I => \N__9275\
        );

    \I__2194\ : Glb2LocalMux
    port map (
            O => \N__9357\,
            I => \N__9275\
        );

    \I__2193\ : SRMux
    port map (
            O => \N__9356\,
            I => \N__9275\
        );

    \I__2192\ : SRMux
    port map (
            O => \N__9355\,
            I => \N__9275\
        );

    \I__2191\ : Glb2LocalMux
    port map (
            O => \N__9352\,
            I => \N__9275\
        );

    \I__2190\ : GlobalMux
    port map (
            O => \N__9275\,
            I => \N__9272\
        );

    \I__2189\ : gio2CtrlBuf
    port map (
            O => \N__9272\,
            I => \RESETn_c_i_g\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__9269\,
            I => \N__9260\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9268\,
            I => \N__9256\
        );

    \I__2186\ : InMux
    port map (
            O => \N__9267\,
            I => \N__9253\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9266\,
            I => \N__9250\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__9265\,
            I => \N__9246\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9264\,
            I => \N__9238\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9238\
        );

    \I__2181\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9233\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9259\,
            I => \N__9233\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9256\,
            I => \N__9228\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9253\,
            I => \N__9228\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__9250\,
            I => \N__9225\
        );

    \I__2176\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9222\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9246\,
            I => \N__9216\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9245\,
            I => \N__9216\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9244\,
            I => \N__9211\
        );

    \I__2172\ : InMux
    port map (
            O => \N__9243\,
            I => \N__9211\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9238\,
            I => \N__9208\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9233\,
            I => \N__9204\
        );

    \I__2169\ : Span4Mux_v
    port map (
            O => \N__9228\,
            I => \N__9199\
        );

    \I__2168\ : Span4Mux_v
    port map (
            O => \N__9225\,
            I => \N__9199\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9222\,
            I => \N__9196\
        );

    \I__2166\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9193\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9216\,
            I => \N__9190\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9211\,
            I => \N__9187\
        );

    \I__2163\ : Span12Mux_v
    port map (
            O => \N__9208\,
            I => \N__9184\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9207\,
            I => \N__9181\
        );

    \I__2161\ : Span4Mux_v
    port map (
            O => \N__9204\,
            I => \N__9174\
        );

    \I__2160\ : Span4Mux_h
    port map (
            O => \N__9199\,
            I => \N__9174\
        );

    \I__2159\ : Span4Mux_v
    port map (
            O => \N__9196\,
            I => \N__9174\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__9193\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__9190\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__9187\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2155\ : Odrv12
    port map (
            O => \N__9184\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9181\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__9174\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__9161\,
            I => \N__9152\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9160\,
            I => \N__9148\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9159\,
            I => \N__9145\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__9158\,
            I => \N__9141\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__9157\,
            I => \N__9138\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__9156\,
            I => \N__9135\
        );

    \I__2146\ : InMux
    port map (
            O => \N__9155\,
            I => \N__9129\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9152\,
            I => \N__9126\
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__9151\,
            I => \N__9122\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9148\,
            I => \N__9119\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9145\,
            I => \N__9116\
        );

    \I__2141\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9113\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9141\,
            I => \N__9106\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9138\,
            I => \N__9106\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9106\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9103\
        );

    \I__2136\ : InMux
    port map (
            O => \N__9133\,
            I => \N__9099\
        );

    \I__2135\ : CascadeMux
    port map (
            O => \N__9132\,
            I => \N__9094\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9129\,
            I => \N__9089\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__9126\,
            I => \N__9089\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__9125\,
            I => \N__9086\
        );

    \I__2131\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9083\
        );

    \I__2130\ : Span4Mux_v
    port map (
            O => \N__9119\,
            I => \N__9078\
        );

    \I__2129\ : Span4Mux_v
    port map (
            O => \N__9116\,
            I => \N__9078\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__9113\,
            I => \N__9073\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__9106\,
            I => \N__9073\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__9103\,
            I => \N__9070\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9067\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9099\,
            I => \N__9064\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9098\,
            I => \N__9061\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9058\
        );

    \I__2121\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9055\
        );

    \I__2120\ : Span4Mux_v
    port map (
            O => \N__9089\,
            I => \N__9052\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9049\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9083\,
            I => \N__9046\
        );

    \I__2117\ : Span4Mux_h
    port map (
            O => \N__9078\,
            I => \N__9039\
        );

    \I__2116\ : Span4Mux_v
    port map (
            O => \N__9073\,
            I => \N__9039\
        );

    \I__2115\ : Span4Mux_v
    port map (
            O => \N__9070\,
            I => \N__9039\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__9067\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__9064\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__9061\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__9058\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9055\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2109\ : Odrv4
    port map (
            O => \N__9052\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__9049\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2107\ : Odrv12
    port map (
            O => \N__9046\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__9039\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__9020\,
            I => \N__9012\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9019\,
            I => \N__9004\
        );

    \I__2103\ : InMux
    port map (
            O => \N__9018\,
            I => \N__9001\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9017\,
            I => \N__8996\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9016\,
            I => \N__8996\
        );

    \I__2100\ : InMux
    port map (
            O => \N__9015\,
            I => \N__8993\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9012\,
            I => \N__8988\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9011\,
            I => \N__8988\
        );

    \I__2097\ : InMux
    port map (
            O => \N__9010\,
            I => \N__8983\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9009\,
            I => \N__8983\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9008\,
            I => \N__8978\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9007\,
            I => \N__8978\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__9004\,
            I => \N__8973\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__9001\,
            I => \N__8973\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__8996\,
            I => \N__8965\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__8993\,
            I => \N__8965\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__8988\,
            I => \N__8956\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__8983\,
            I => \N__8956\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__8978\,
            I => \N__8956\
        );

    \I__2086\ : Span4Mux_h
    port map (
            O => \N__8973\,
            I => \N__8956\
        );

    \I__2085\ : InMux
    port map (
            O => \N__8972\,
            I => \N__8953\
        );

    \I__2084\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8950\
        );

    \I__2083\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8947\
        );

    \I__2082\ : Span4Mux_h
    port map (
            O => \N__8965\,
            I => \N__8944\
        );

    \I__2081\ : Span4Mux_h
    port map (
            O => \N__8956\,
            I => \N__8939\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__8953\,
            I => \N__8939\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__8950\,
            I => \N__8936\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__8947\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2077\ : Odrv4
    port map (
            O => \N__8944\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__8939\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__8936\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2074\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8921\
        );

    \I__2073\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8921\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__8921\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__2071\ : InMux
    port map (
            O => \N__8918\,
            I => \N__8915\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__8915\,
            I => \N__8911\
        );

    \I__2069\ : InMux
    port map (
            O => \N__8914\,
            I => \N__8908\
        );

    \I__2068\ : Span4Mux_h
    port map (
            O => \N__8911\,
            I => \N__8903\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__8908\,
            I => \N__8903\
        );

    \I__2066\ : Span4Mux_v
    port map (
            O => \N__8903\,
            I => \N__8900\
        );

    \I__2065\ : Sp12to4
    port map (
            O => \N__8900\,
            I => \N__8897\
        );

    \I__2064\ : Span12Mux_h
    port map (
            O => \N__8897\,
            I => \N__8894\
        );

    \I__2063\ : Odrv12
    port map (
            O => \N__8894\,
            I => \DRA_c_8\
        );

    \I__2062\ : CEMux
    port map (
            O => \N__8891\,
            I => \N__8888\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__8888\,
            I => \N__8884\
        );

    \I__2060\ : CEMux
    port map (
            O => \N__8887\,
            I => \N__8881\
        );

    \I__2059\ : Odrv12
    port map (
            O => \N__8884\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__8881\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__2057\ : IoInMux
    port map (
            O => \N__8876\,
            I => \N__8873\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__8873\,
            I => \N__8870\
        );

    \I__2055\ : Span12Mux_s8_v
    port map (
            O => \N__8870\,
            I => \N__8867\
        );

    \I__2054\ : Odrv12
    port map (
            O => \N__8867\,
            I => \CASn_c\
        );

    \I__2053\ : IoInMux
    port map (
            O => \N__8864\,
            I => \N__8861\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__8861\,
            I => \N__8858\
        );

    \I__2051\ : IoSpan4Mux
    port map (
            O => \N__8858\,
            I => \N__8855\
        );

    \I__2050\ : IoSpan4Mux
    port map (
            O => \N__8855\,
            I => \N__8852\
        );

    \I__2049\ : Sp12to4
    port map (
            O => \N__8852\,
            I => \N__8849\
        );

    \I__2048\ : Span12Mux_s9_v
    port map (
            O => \N__8849\,
            I => \N__8846\
        );

    \I__2047\ : Odrv12
    port map (
            O => \N__8846\,
            I => \WEn_c\
        );

    \I__2046\ : IoInMux
    port map (
            O => \N__8843\,
            I => \N__8840\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__8840\,
            I => \N__8837\
        );

    \I__2044\ : Span4Mux_s3_v
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__2043\ : Span4Mux_v
    port map (
            O => \N__8834\,
            I => \N__8831\
        );

    \I__2042\ : Span4Mux_h
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__8828\,
            I => \RASn_c\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__8825\,
            I => \N__8820\
        );

    \I__2039\ : InMux
    port map (
            O => \N__8824\,
            I => \N__8817\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__8823\,
            I => \N__8814\
        );

    \I__2037\ : InMux
    port map (
            O => \N__8820\,
            I => \N__8811\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__8817\,
            I => \N__8808\
        );

    \I__2035\ : InMux
    port map (
            O => \N__8814\,
            I => \N__8805\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__8811\,
            I => \N__8801\
        );

    \I__2033\ : Span4Mux_v
    port map (
            O => \N__8808\,
            I => \N__8798\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__8805\,
            I => \N__8794\
        );

    \I__2031\ : InMux
    port map (
            O => \N__8804\,
            I => \N__8791\
        );

    \I__2030\ : Span4Mux_v
    port map (
            O => \N__8801\,
            I => \N__8786\
        );

    \I__2029\ : Span4Mux_h
    port map (
            O => \N__8798\,
            I => \N__8786\
        );

    \I__2028\ : InMux
    port map (
            O => \N__8797\,
            I => \N__8783\
        );

    \I__2027\ : Span4Mux_h
    port map (
            O => \N__8794\,
            I => \N__8780\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__8791\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2025\ : Odrv4
    port map (
            O => \N__8786\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__8783\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__8780\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2022\ : IoInMux
    port map (
            O => \N__8771\,
            I => \N__8768\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__8768\,
            I => \N__8765\
        );

    \I__2020\ : Span4Mux_s2_v
    port map (
            O => \N__8765\,
            I => \N__8762\
        );

    \I__2019\ : Span4Mux_v
    port map (
            O => \N__8762\,
            I => \N__8759\
        );

    \I__2018\ : Span4Mux_v
    port map (
            O => \N__8759\,
            I => \N__8756\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__8756\,
            I => \CRCSn_c\
        );

    \I__2016\ : InMux
    port map (
            O => \N__8753\,
            I => \N__8750\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__8750\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__2014\ : InMux
    port map (
            O => \N__8747\,
            I => \N__8744\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__8744\,
            I => \N__8741\
        );

    \I__2012\ : Span4Mux_v
    port map (
            O => \N__8741\,
            I => \N__8738\
        );

    \I__2011\ : Sp12to4
    port map (
            O => \N__8738\,
            I => \N__8735\
        );

    \I__2010\ : Odrv12
    port map (
            O => \N__8735\,
            I => \RAS1n_c\
        );

    \I__2009\ : InMux
    port map (
            O => \N__8732\,
            I => \N__8728\
        );

    \I__2008\ : InMux
    port map (
            O => \N__8731\,
            I => \N__8725\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__8728\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__8725\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2005\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8717\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__8717\,
            I => \N__8714\
        );

    \I__2003\ : Span12Mux_v
    port map (
            O => \N__8714\,
            I => \N__8711\
        );

    \I__2002\ : Span12Mux_h
    port map (
            O => \N__8711\,
            I => \N__8708\
        );

    \I__2001\ : Odrv12
    port map (
            O => \N__8708\,
            I => \A_c_17\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__8705\,
            I => \N__8702\
        );

    \I__1999\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8699\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__8699\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1997\ : IoInMux
    port map (
            O => \N__8696\,
            I => \N__8693\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__8693\,
            I => \N__8690\
        );

    \I__1995\ : IoSpan4Mux
    port map (
            O => \N__8690\,
            I => \N__8687\
        );

    \I__1994\ : Span4Mux_s3_h
    port map (
            O => \N__8687\,
            I => \N__8684\
        );

    \I__1993\ : Span4Mux_v
    port map (
            O => \N__8684\,
            I => \N__8681\
        );

    \I__1992\ : Sp12to4
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__1991\ : Odrv12
    port map (
            O => \N__8678\,
            I => \CMA_c_8\
        );

    \I__1990\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__1988\ : Span12Mux_v
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__1987\ : Span12Mux_h
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__1986\ : Odrv12
    port map (
            O => \N__8663\,
            I => \A_c_19\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__8660\,
            I => \N__8656\
        );

    \I__1984\ : InMux
    port map (
            O => \N__8659\,
            I => \N__8653\
        );

    \I__1983\ : InMux
    port map (
            O => \N__8656\,
            I => \N__8650\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__8653\,
            I => \N__8645\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__8650\,
            I => \N__8645\
        );

    \I__1980\ : Span12Mux_v
    port map (
            O => \N__8645\,
            I => \N__8642\
        );

    \I__1979\ : Span12Mux_h
    port map (
            O => \N__8642\,
            I => \N__8639\
        );

    \I__1978\ : Odrv12
    port map (
            O => \N__8639\,
            I => \RAS0n_c\
        );

    \I__1977\ : CascadeMux
    port map (
            O => \N__8636\,
            I => \N__8626\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__8635\,
            I => \N__8622\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__8634\,
            I => \N__8619\
        );

    \I__1974\ : InMux
    port map (
            O => \N__8633\,
            I => \N__8610\
        );

    \I__1973\ : InMux
    port map (
            O => \N__8632\,
            I => \N__8610\
        );

    \I__1972\ : InMux
    port map (
            O => \N__8631\,
            I => \N__8607\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__8630\,
            I => \N__8602\
        );

    \I__1970\ : InMux
    port map (
            O => \N__8629\,
            I => \N__8599\
        );

    \I__1969\ : InMux
    port map (
            O => \N__8626\,
            I => \N__8587\
        );

    \I__1968\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8581\
        );

    \I__1967\ : InMux
    port map (
            O => \N__8622\,
            I => \N__8581\
        );

    \I__1966\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8578\
        );

    \I__1965\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8571\
        );

    \I__1964\ : InMux
    port map (
            O => \N__8617\,
            I => \N__8571\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8571\
        );

    \I__1962\ : InMux
    port map (
            O => \N__8615\,
            I => \N__8566\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__8610\,
            I => \N__8561\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__8607\,
            I => \N__8561\
        );

    \I__1959\ : InMux
    port map (
            O => \N__8606\,
            I => \N__8556\
        );

    \I__1958\ : InMux
    port map (
            O => \N__8605\,
            I => \N__8556\
        );

    \I__1957\ : InMux
    port map (
            O => \N__8602\,
            I => \N__8553\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__8599\,
            I => \N__8550\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8598\,
            I => \N__8541\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8597\,
            I => \N__8541\
        );

    \I__1953\ : InMux
    port map (
            O => \N__8596\,
            I => \N__8541\
        );

    \I__1952\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8541\
        );

    \I__1951\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8530\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8593\,
            I => \N__8530\
        );

    \I__1949\ : InMux
    port map (
            O => \N__8592\,
            I => \N__8530\
        );

    \I__1948\ : InMux
    port map (
            O => \N__8591\,
            I => \N__8530\
        );

    \I__1947\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8530\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__8587\,
            I => \N__8527\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8586\,
            I => \N__8524\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__8581\,
            I => \N__8519\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__8578\,
            I => \N__8516\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__8571\,
            I => \N__8513\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8510\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8507\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__8566\,
            I => \N__8502\
        );

    \I__1938\ : Span4Mux_h
    port map (
            O => \N__8561\,
            I => \N__8502\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__8556\,
            I => \N__8491\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8553\,
            I => \N__8491\
        );

    \I__1935\ : Span4Mux_h
    port map (
            O => \N__8550\,
            I => \N__8491\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__8541\,
            I => \N__8491\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__8530\,
            I => \N__8491\
        );

    \I__1932\ : Span4Mux_v
    port map (
            O => \N__8527\,
            I => \N__8486\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__8524\,
            I => \N__8486\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8523\,
            I => \N__8483\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8480\
        );

    \I__1928\ : Span4Mux_v
    port map (
            O => \N__8519\,
            I => \N__8475\
        );

    \I__1927\ : Span4Mux_h
    port map (
            O => \N__8516\,
            I => \N__8475\
        );

    \I__1926\ : Span12Mux_v
    port map (
            O => \N__8513\,
            I => \N__8468\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__8510\,
            I => \N__8468\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8507\,
            I => \N__8468\
        );

    \I__1923\ : Span4Mux_h
    port map (
            O => \N__8502\,
            I => \N__8465\
        );

    \I__1922\ : Span4Mux_h
    port map (
            O => \N__8491\,
            I => \N__8462\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__8486\,
            I => \CPU_CYCLEm\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__8483\,
            I => \CPU_CYCLEm\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__8480\,
            I => \CPU_CYCLEm\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__8475\,
            I => \CPU_CYCLEm\
        );

    \I__1917\ : Odrv12
    port map (
            O => \N__8468\,
            I => \CPU_CYCLEm\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__8465\,
            I => \CPU_CYCLEm\
        );

    \I__1915\ : Odrv4
    port map (
            O => \N__8462\,
            I => \CPU_CYCLEm\
        );

    \I__1914\ : IoInMux
    port map (
            O => \N__8447\,
            I => \N__8444\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__8444\,
            I => \N__8441\
        );

    \I__1912\ : Sp12to4
    port map (
            O => \N__8441\,
            I => \N__8438\
        );

    \I__1911\ : Span12Mux_h
    port map (
            O => \N__8438\,
            I => \N__8435\
        );

    \I__1910\ : Odrv12
    port map (
            O => \N__8435\,
            I => \CMA_c_9\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8432\,
            I => \N__8429\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8429\,
            I => \N__8395\
        );

    \I__1907\ : ClkMux
    port map (
            O => \N__8428\,
            I => \N__8297\
        );

    \I__1906\ : ClkMux
    port map (
            O => \N__8427\,
            I => \N__8297\
        );

    \I__1905\ : ClkMux
    port map (
            O => \N__8426\,
            I => \N__8297\
        );

    \I__1904\ : ClkMux
    port map (
            O => \N__8425\,
            I => \N__8297\
        );

    \I__1903\ : ClkMux
    port map (
            O => \N__8424\,
            I => \N__8297\
        );

    \I__1902\ : ClkMux
    port map (
            O => \N__8423\,
            I => \N__8297\
        );

    \I__1901\ : ClkMux
    port map (
            O => \N__8422\,
            I => \N__8297\
        );

    \I__1900\ : ClkMux
    port map (
            O => \N__8421\,
            I => \N__8297\
        );

    \I__1899\ : ClkMux
    port map (
            O => \N__8420\,
            I => \N__8297\
        );

    \I__1898\ : ClkMux
    port map (
            O => \N__8419\,
            I => \N__8297\
        );

    \I__1897\ : ClkMux
    port map (
            O => \N__8418\,
            I => \N__8297\
        );

    \I__1896\ : ClkMux
    port map (
            O => \N__8417\,
            I => \N__8297\
        );

    \I__1895\ : ClkMux
    port map (
            O => \N__8416\,
            I => \N__8297\
        );

    \I__1894\ : ClkMux
    port map (
            O => \N__8415\,
            I => \N__8297\
        );

    \I__1893\ : ClkMux
    port map (
            O => \N__8414\,
            I => \N__8297\
        );

    \I__1892\ : ClkMux
    port map (
            O => \N__8413\,
            I => \N__8297\
        );

    \I__1891\ : ClkMux
    port map (
            O => \N__8412\,
            I => \N__8297\
        );

    \I__1890\ : ClkMux
    port map (
            O => \N__8411\,
            I => \N__8297\
        );

    \I__1889\ : ClkMux
    port map (
            O => \N__8410\,
            I => \N__8297\
        );

    \I__1888\ : ClkMux
    port map (
            O => \N__8409\,
            I => \N__8297\
        );

    \I__1887\ : ClkMux
    port map (
            O => \N__8408\,
            I => \N__8297\
        );

    \I__1886\ : ClkMux
    port map (
            O => \N__8407\,
            I => \N__8297\
        );

    \I__1885\ : ClkMux
    port map (
            O => \N__8406\,
            I => \N__8297\
        );

    \I__1884\ : ClkMux
    port map (
            O => \N__8405\,
            I => \N__8297\
        );

    \I__1883\ : ClkMux
    port map (
            O => \N__8404\,
            I => \N__8297\
        );

    \I__1882\ : ClkMux
    port map (
            O => \N__8403\,
            I => \N__8297\
        );

    \I__1881\ : ClkMux
    port map (
            O => \N__8402\,
            I => \N__8297\
        );

    \I__1880\ : ClkMux
    port map (
            O => \N__8401\,
            I => \N__8297\
        );

    \I__1879\ : ClkMux
    port map (
            O => \N__8400\,
            I => \N__8297\
        );

    \I__1878\ : ClkMux
    port map (
            O => \N__8399\,
            I => \N__8297\
        );

    \I__1877\ : ClkMux
    port map (
            O => \N__8398\,
            I => \N__8297\
        );

    \I__1876\ : Glb2LocalMux
    port map (
            O => \N__8395\,
            I => \N__8297\
        );

    \I__1875\ : ClkMux
    port map (
            O => \N__8394\,
            I => \N__8297\
        );

    \I__1874\ : ClkMux
    port map (
            O => \N__8393\,
            I => \N__8297\
        );

    \I__1873\ : ClkMux
    port map (
            O => \N__8392\,
            I => \N__8297\
        );

    \I__1872\ : ClkMux
    port map (
            O => \N__8391\,
            I => \N__8297\
        );

    \I__1871\ : ClkMux
    port map (
            O => \N__8390\,
            I => \N__8297\
        );

    \I__1870\ : ClkMux
    port map (
            O => \N__8389\,
            I => \N__8297\
        );

    \I__1869\ : ClkMux
    port map (
            O => \N__8388\,
            I => \N__8297\
        );

    \I__1868\ : ClkMux
    port map (
            O => \N__8387\,
            I => \N__8297\
        );

    \I__1867\ : ClkMux
    port map (
            O => \N__8386\,
            I => \N__8297\
        );

    \I__1866\ : ClkMux
    port map (
            O => \N__8385\,
            I => \N__8297\
        );

    \I__1865\ : ClkMux
    port map (
            O => \N__8384\,
            I => \N__8297\
        );

    \I__1864\ : GlobalMux
    port map (
            O => \N__8297\,
            I => \CLK80_OUT\
        );

    \I__1863\ : CEMux
    port map (
            O => \N__8294\,
            I => \N__8288\
        );

    \I__1862\ : CEMux
    port map (
            O => \N__8293\,
            I => \N__8285\
        );

    \I__1861\ : CEMux
    port map (
            O => \N__8292\,
            I => \N__8282\
        );

    \I__1860\ : CEMux
    port map (
            O => \N__8291\,
            I => \N__8279\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__8288\,
            I => \N__8275\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__8285\,
            I => \N__8272\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__8282\,
            I => \N__8268\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8279\,
            I => \N__8265\
        );

    \I__1855\ : CEMux
    port map (
            O => \N__8278\,
            I => \N__8262\
        );

    \I__1854\ : Span4Mux_h
    port map (
            O => \N__8275\,
            I => \N__8257\
        );

    \I__1853\ : Span4Mux_v
    port map (
            O => \N__8272\,
            I => \N__8257\
        );

    \I__1852\ : CEMux
    port map (
            O => \N__8271\,
            I => \N__8254\
        );

    \I__1851\ : Span4Mux_h
    port map (
            O => \N__8268\,
            I => \N__8251\
        );

    \I__1850\ : Span4Mux_v
    port map (
            O => \N__8265\,
            I => \N__8248\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8262\,
            I => \N__8243\
        );

    \I__1848\ : Span4Mux_h
    port map (
            O => \N__8257\,
            I => \N__8243\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__8254\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__8251\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1845\ : Odrv4
    port map (
            O => \N__8248\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__8243\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8234\,
            I => \N__8231\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__8231\,
            I => \N__8228\
        );

    \I__1841\ : Span4Mux_h
    port map (
            O => \N__8228\,
            I => \N__8225\
        );

    \I__1840\ : Span4Mux_v
    port map (
            O => \N__8225\,
            I => \N__8222\
        );

    \I__1839\ : Span4Mux_h
    port map (
            O => \N__8222\,
            I => \N__8219\
        );

    \I__1838\ : Sp12to4
    port map (
            O => \N__8219\,
            I => \N__8216\
        );

    \I__1837\ : Odrv12
    port map (
            O => \N__8216\,
            I => \A_c_8\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__8213\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_6_cascade_\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8210\,
            I => \N__8207\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__8207\,
            I => \N__8204\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__8204\,
            I => \N__8201\
        );

    \I__1832\ : Span4Mux_v
    port map (
            O => \N__8201\,
            I => \N__8198\
        );

    \I__1831\ : Sp12to4
    port map (
            O => \N__8198\,
            I => \N__8195\
        );

    \I__1830\ : Span12Mux_h
    port map (
            O => \N__8195\,
            I => \N__8192\
        );

    \I__1829\ : Odrv12
    port map (
            O => \N__8192\,
            I => \A_c_15\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8189\,
            I => \N__8186\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8186\,
            I => \U712_CHIP_RAM.N_37\
        );

    \I__1826\ : InMux
    port map (
            O => \N__8183\,
            I => \N__8180\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__8180\,
            I => \N__8175\
        );

    \I__1824\ : InMux
    port map (
            O => \N__8179\,
            I => \N__8170\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8178\,
            I => \N__8170\
        );

    \I__1822\ : Span4Mux_v
    port map (
            O => \N__8175\,
            I => \N__8167\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8170\,
            I => \N__8164\
        );

    \I__1820\ : Sp12to4
    port map (
            O => \N__8167\,
            I => \N__8161\
        );

    \I__1819\ : Span12Mux_v
    port map (
            O => \N__8164\,
            I => \N__8158\
        );

    \I__1818\ : Span12Mux_h
    port map (
            O => \N__8161\,
            I => \N__8155\
        );

    \I__1817\ : Span12Mux_h
    port map (
            O => \N__8158\,
            I => \N__8152\
        );

    \I__1816\ : Span12Mux_v
    port map (
            O => \N__8155\,
            I => \N__8149\
        );

    \I__1815\ : Odrv12
    port map (
            O => \N__8152\,
            I => \CASLn_c\
        );

    \I__1814\ : Odrv12
    port map (
            O => \N__8149\,
            I => \CASLn_c\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8144\,
            I => \N__8140\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8143\,
            I => \N__8137\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8140\,
            I => \N__8133\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8137\,
            I => \N__8130\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8136\,
            I => \N__8127\
        );

    \I__1808\ : Span4Mux_h
    port map (
            O => \N__8133\,
            I => \N__8124\
        );

    \I__1807\ : Span4Mux_v
    port map (
            O => \N__8130\,
            I => \N__8119\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__8127\,
            I => \N__8119\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__8124\,
            I => \N__8116\
        );

    \I__1804\ : Sp12to4
    port map (
            O => \N__8119\,
            I => \N__8113\
        );

    \I__1803\ : Sp12to4
    port map (
            O => \N__8116\,
            I => \N__8110\
        );

    \I__1802\ : Span12Mux_h
    port map (
            O => \N__8113\,
            I => \N__8107\
        );

    \I__1801\ : Span12Mux_v
    port map (
            O => \N__8110\,
            I => \N__8104\
        );

    \I__1800\ : Span12Mux_v
    port map (
            O => \N__8107\,
            I => \N__8101\
        );

    \I__1799\ : Span12Mux_h
    port map (
            O => \N__8104\,
            I => \N__8098\
        );

    \I__1798\ : Odrv12
    port map (
            O => \N__8101\,
            I => \CASUn_c\
        );

    \I__1797\ : Odrv12
    port map (
            O => \N__8098\,
            I => \CASUn_c\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8093\,
            I => \N__8089\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8092\,
            I => \N__8086\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__8089\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8086\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8081\,
            I => \N__8078\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__8078\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1790\ : IoInMux
    port map (
            O => \N__8075\,
            I => \N__8072\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__8072\,
            I => \N__8069\
        );

    \I__1788\ : Sp12to4
    port map (
            O => \N__8069\,
            I => \N__8066\
        );

    \I__1787\ : Span12Mux_h
    port map (
            O => \N__8066\,
            I => \N__8063\
        );

    \I__1786\ : Odrv12
    port map (
            O => \N__8063\,
            I => \CMA_c_7\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8060\,
            I => \N__8057\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8057\,
            I => \N__8054\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__8054\,
            I => \N__8051\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__8051\,
            I => \N__8048\
        );

    \I__1781\ : Sp12to4
    port map (
            O => \N__8048\,
            I => \N__8045\
        );

    \I__1780\ : Span12Mux_h
    port map (
            O => \N__8045\,
            I => \N__8042\
        );

    \I__1779\ : Odrv12
    port map (
            O => \N__8042\,
            I => \A_c_18\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__8039\,
            I => \N__8036\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8036\,
            I => \N__8033\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__8033\,
            I => \N__8030\
        );

    \I__1775\ : Span4Mux_v
    port map (
            O => \N__8030\,
            I => \N__8027\
        );

    \I__1774\ : Span4Mux_v
    port map (
            O => \N__8027\,
            I => \N__8024\
        );

    \I__1773\ : Sp12to4
    port map (
            O => \N__8024\,
            I => \N__8021\
        );

    \I__1772\ : Span12Mux_h
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__1771\ : Odrv12
    port map (
            O => \N__8018\,
            I => \A_c_16\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__8012\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_7\
        );

    \I__1768\ : InMux
    port map (
            O => \N__8009\,
            I => \N__8006\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__8006\,
            I => \U712_CHIP_RAM.N_38\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8003\,
            I => \N__7999\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8002\,
            I => \N__7996\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__7999\,
            I => \N__7993\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__7996\,
            I => \N__7990\
        );

    \I__1762\ : Span4Mux_v
    port map (
            O => \N__7993\,
            I => \N__7987\
        );

    \I__1761\ : Sp12to4
    port map (
            O => \N__7990\,
            I => \N__7984\
        );

    \I__1760\ : Span4Mux_v
    port map (
            O => \N__7987\,
            I => \N__7981\
        );

    \I__1759\ : Span12Mux_v
    port map (
            O => \N__7984\,
            I => \N__7976\
        );

    \I__1758\ : Sp12to4
    port map (
            O => \N__7981\,
            I => \N__7976\
        );

    \I__1757\ : Span12Mux_h
    port map (
            O => \N__7976\,
            I => \N__7973\
        );

    \I__1756\ : Odrv12
    port map (
            O => \N__7973\,
            I => \DRA_c_6\
        );

    \I__1755\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7967\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__7967\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__1753\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7961\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__7961\,
            I => \N__7957\
        );

    \I__1751\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7954\
        );

    \I__1750\ : Span4Mux_h
    port map (
            O => \N__7957\,
            I => \N__7949\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__7954\,
            I => \N__7949\
        );

    \I__1748\ : Span4Mux_h
    port map (
            O => \N__7949\,
            I => \N__7946\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__7946\,
            I => \N__7943\
        );

    \I__1746\ : Sp12to4
    port map (
            O => \N__7943\,
            I => \N__7940\
        );

    \I__1745\ : Odrv12
    port map (
            O => \N__7940\,
            I => \DRA_c_7\
        );

    \I__1744\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7934\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__7934\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__1742\ : IoInMux
    port map (
            O => \N__7931\,
            I => \N__7928\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__1740\ : Span4Mux_s0_v
    port map (
            O => \N__7925\,
            I => \N__7922\
        );

    \I__1739\ : Sp12to4
    port map (
            O => \N__7922\,
            I => \N__7919\
        );

    \I__1738\ : Span12Mux_h
    port map (
            O => \N__7919\,
            I => \N__7916\
        );

    \I__1737\ : Span12Mux_v
    port map (
            O => \N__7916\,
            I => \N__7913\
        );

    \I__1736\ : Odrv12
    port map (
            O => \N__7913\,
            I => \CMA_c_10\
        );

    \I__1735\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7906\
        );

    \I__1734\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7903\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__7906\,
            I => \N__7900\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__7903\,
            I => \N__7897\
        );

    \I__1731\ : Span12Mux_h
    port map (
            O => \N__7900\,
            I => \N__7894\
        );

    \I__1730\ : Span12Mux_h
    port map (
            O => \N__7897\,
            I => \N__7891\
        );

    \I__1729\ : Span12Mux_v
    port map (
            O => \N__7894\,
            I => \N__7888\
        );

    \I__1728\ : Span12Mux_v
    port map (
            O => \N__7891\,
            I => \N__7885\
        );

    \I__1727\ : Odrv12
    port map (
            O => \N__7888\,
            I => \DRA_c_2\
        );

    \I__1726\ : Odrv12
    port map (
            O => \N__7885\,
            I => \DRA_c_2\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__7880\,
            I => \N__7877\
        );

    \I__1724\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7874\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__7874\,
            I => \N__7871\
        );

    \I__1722\ : Odrv12
    port map (
            O => \N__7871\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1721\ : InMux
    port map (
            O => \N__7868\,
            I => \N__7865\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__7865\,
            I => \N__7861\
        );

    \I__1719\ : InMux
    port map (
            O => \N__7864\,
            I => \N__7858\
        );

    \I__1718\ : Sp12to4
    port map (
            O => \N__7861\,
            I => \N__7853\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__7858\,
            I => \N__7853\
        );

    \I__1716\ : Span12Mux_v
    port map (
            O => \N__7853\,
            I => \N__7850\
        );

    \I__1715\ : Span12Mux_h
    port map (
            O => \N__7850\,
            I => \N__7847\
        );

    \I__1714\ : Odrv12
    port map (
            O => \N__7847\,
            I => \DRA_c_5\
        );

    \I__1713\ : InMux
    port map (
            O => \N__7844\,
            I => \N__7841\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__7841\,
            I => \N__7838\
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__7838\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1710\ : InMux
    port map (
            O => \N__7835\,
            I => \N__7831\
        );

    \I__1709\ : InMux
    port map (
            O => \N__7834\,
            I => \N__7828\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__7831\,
            I => \N__7825\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__7828\,
            I => \N__7822\
        );

    \I__1706\ : Span4Mux_h
    port map (
            O => \N__7825\,
            I => \N__7819\
        );

    \I__1705\ : Span4Mux_v
    port map (
            O => \N__7822\,
            I => \N__7816\
        );

    \I__1704\ : Sp12to4
    port map (
            O => \N__7819\,
            I => \N__7813\
        );

    \I__1703\ : Sp12to4
    port map (
            O => \N__7816\,
            I => \N__7810\
        );

    \I__1702\ : Span12Mux_v
    port map (
            O => \N__7813\,
            I => \N__7807\
        );

    \I__1701\ : Span12Mux_h
    port map (
            O => \N__7810\,
            I => \N__7804\
        );

    \I__1700\ : Span12Mux_h
    port map (
            O => \N__7807\,
            I => \N__7799\
        );

    \I__1699\ : Span12Mux_v
    port map (
            O => \N__7804\,
            I => \N__7799\
        );

    \I__1698\ : Odrv12
    port map (
            O => \N__7799\,
            I => \DRA_c_4\
        );

    \I__1697\ : InMux
    port map (
            O => \N__7796\,
            I => \N__7793\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__7793\,
            I => \N__7790\
        );

    \I__1695\ : Odrv12
    port map (
            O => \N__7790\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1694\ : InMux
    port map (
            O => \N__7787\,
            I => \N__7784\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__7784\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1692\ : CEMux
    port map (
            O => \N__7781\,
            I => \N__7777\
        );

    \I__1691\ : CEMux
    port map (
            O => \N__7780\,
            I => \N__7774\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__7777\,
            I => \N__7771\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__7774\,
            I => \N__7768\
        );

    \I__1688\ : Odrv4
    port map (
            O => \N__7771\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__7768\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__7763\,
            I => \N__7760\
        );

    \I__1685\ : InMux
    port map (
            O => \N__7760\,
            I => \N__7757\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__7757\,
            I => \N__7753\
        );

    \I__1683\ : InMux
    port map (
            O => \N__7756\,
            I => \N__7750\
        );

    \I__1682\ : Odrv12
    port map (
            O => \N__7753\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__7750\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4\
        );

    \I__1680\ : InMux
    port map (
            O => \N__7745\,
            I => \N__7742\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__7742\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1678\ : InMux
    port map (
            O => \N__7739\,
            I => \N__7736\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__7736\,
            I => \N__7733\
        );

    \I__1676\ : Odrv12
    port map (
            O => \N__7733\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1675\ : InMux
    port map (
            O => \N__7730\,
            I => \N__7727\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__7727\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1673\ : InMux
    port map (
            O => \N__7724\,
            I => \N__7721\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__7721\,
            I => \N__7718\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__7718\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__1670\ : InMux
    port map (
            O => \N__7715\,
            I => \N__7712\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__7712\,
            I => \N__7708\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7711\,
            I => \N__7705\
        );

    \I__1667\ : Span4Mux_h
    port map (
            O => \N__7708\,
            I => \N__7700\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__7705\,
            I => \N__7700\
        );

    \I__1665\ : Span4Mux_v
    port map (
            O => \N__7700\,
            I => \N__7697\
        );

    \I__1664\ : Sp12to4
    port map (
            O => \N__7697\,
            I => \N__7694\
        );

    \I__1663\ : Span12Mux_h
    port map (
            O => \N__7694\,
            I => \N__7691\
        );

    \I__1662\ : Span12Mux_v
    port map (
            O => \N__7691\,
            I => \N__7688\
        );

    \I__1661\ : Odrv12
    port map (
            O => \N__7688\,
            I => \DRA_c_1\
        );

    \I__1660\ : InMux
    port map (
            O => \N__7685\,
            I => \N__7682\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__7682\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1658\ : InMux
    port map (
            O => \N__7679\,
            I => \N__7676\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__7676\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1656\ : InMux
    port map (
            O => \N__7673\,
            I => \N__7670\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__7670\,
            I => \N__7666\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7669\,
            I => \N__7663\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__7666\,
            I => \N__7658\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__7663\,
            I => \N__7658\
        );

    \I__1651\ : Span4Mux_h
    port map (
            O => \N__7658\,
            I => \N__7655\
        );

    \I__1650\ : Span4Mux_v
    port map (
            O => \N__7655\,
            I => \N__7652\
        );

    \I__1649\ : Sp12to4
    port map (
            O => \N__7652\,
            I => \N__7649\
        );

    \I__1648\ : Span12Mux_h
    port map (
            O => \N__7649\,
            I => \N__7646\
        );

    \I__1647\ : Span12Mux_v
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__1646\ : Odrv12
    port map (
            O => \N__7643\,
            I => \DRA_c_0\
        );

    \I__1645\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7637\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7637\,
            I => \N__7634\
        );

    \I__1643\ : Odrv12
    port map (
            O => \N__7634\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1642\ : InMux
    port map (
            O => \N__7631\,
            I => \N__7628\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7628\,
            I => \N__7624\
        );

    \I__1640\ : InMux
    port map (
            O => \N__7627\,
            I => \N__7621\
        );

    \I__1639\ : Span4Mux_h
    port map (
            O => \N__7624\,
            I => \N__7616\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__7621\,
            I => \N__7616\
        );

    \I__1637\ : Sp12to4
    port map (
            O => \N__7616\,
            I => \N__7613\
        );

    \I__1636\ : Span12Mux_v
    port map (
            O => \N__7613\,
            I => \N__7610\
        );

    \I__1635\ : Span12Mux_h
    port map (
            O => \N__7610\,
            I => \N__7607\
        );

    \I__1634\ : Odrv12
    port map (
            O => \N__7607\,
            I => \DRA_c_3\
        );

    \I__1633\ : InMux
    port map (
            O => \N__7604\,
            I => \N__7601\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__7601\,
            I => \N__7598\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__7598\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1630\ : IoInMux
    port map (
            O => \N__7595\,
            I => \N__7592\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__7592\,
            I => \N__7589\
        );

    \I__1628\ : Span12Mux_s3_h
    port map (
            O => \N__7589\,
            I => \N__7586\
        );

    \I__1627\ : Span12Mux_h
    port map (
            O => \N__7586\,
            I => \N__7583\
        );

    \I__1626\ : Odrv12
    port map (
            O => \N__7583\,
            I => \CMA_c_6\
        );

    \I__1625\ : InMux
    port map (
            O => \N__7580\,
            I => \N__7577\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7577\,
            I => \N__7574\
        );

    \I__1623\ : Span4Mux_v
    port map (
            O => \N__7574\,
            I => \N__7571\
        );

    \I__1622\ : Span4Mux_v
    port map (
            O => \N__7571\,
            I => \N__7568\
        );

    \I__1621\ : Sp12to4
    port map (
            O => \N__7568\,
            I => \N__7565\
        );

    \I__1620\ : Span12Mux_h
    port map (
            O => \N__7565\,
            I => \N__7562\
        );

    \I__1619\ : Odrv12
    port map (
            O => \N__7562\,
            I => \A_c_14\
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__7559\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_5_cascade_\
        );

    \I__1617\ : InMux
    port map (
            O => \N__7556\,
            I => \N__7553\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__7553\,
            I => \N__7550\
        );

    \I__1615\ : Span12Mux_v
    port map (
            O => \N__7550\,
            I => \N__7547\
        );

    \I__1614\ : Span12Mux_h
    port map (
            O => \N__7547\,
            I => \N__7544\
        );

    \I__1613\ : Odrv12
    port map (
            O => \N__7544\,
            I => \A_c_7\
        );

    \I__1612\ : InMux
    port map (
            O => \N__7541\,
            I => \N__7538\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__7538\,
            I => \N__7535\
        );

    \I__1610\ : Odrv4
    port map (
            O => \N__7535\,
            I => \U712_CHIP_RAM.N_36\
        );

    \I__1609\ : InMux
    port map (
            O => \N__7532\,
            I => \N__7529\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__7529\,
            I => \N__7526\
        );

    \I__1607\ : Span4Mux_v
    port map (
            O => \N__7526\,
            I => \N__7523\
        );

    \I__1606\ : Sp12to4
    port map (
            O => \N__7523\,
            I => \N__7520\
        );

    \I__1605\ : Span12Mux_h
    port map (
            O => \N__7520\,
            I => \N__7517\
        );

    \I__1604\ : Span12Mux_v
    port map (
            O => \N__7517\,
            I => \N__7514\
        );

    \I__1603\ : Odrv12
    port map (
            O => \N__7514\,
            I => \A_c_4\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__7511\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7508\,
            I => \N__7505\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7505\,
            I => \N__7502\
        );

    \I__1599\ : Span12Mux_s11_v
    port map (
            O => \N__7502\,
            I => \N__7499\
        );

    \I__1598\ : Span12Mux_h
    port map (
            O => \N__7499\,
            I => \N__7496\
        );

    \I__1597\ : Odrv12
    port map (
            O => \N__7496\,
            I => \A_c_11\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7493\,
            I => \N__7490\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7490\,
            I => \U712_CHIP_RAM.N_33\
        );

    \I__1594\ : InMux
    port map (
            O => \N__7487\,
            I => \N__7484\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__7484\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_0\
        );

    \I__1592\ : InMux
    port map (
            O => \N__7481\,
            I => \N__7478\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__7478\,
            I => \N__7475\
        );

    \I__1590\ : Span4Mux_h
    port map (
            O => \N__7475\,
            I => \N__7469\
        );

    \I__1589\ : InMux
    port map (
            O => \N__7474\,
            I => \N__7466\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7473\,
            I => \N__7461\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7472\,
            I => \N__7461\
        );

    \I__1586\ : Odrv4
    port map (
            O => \N__7469\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7466\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7461\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__7454\,
            I => \N__7451\
        );

    \I__1582\ : InMux
    port map (
            O => \N__7451\,
            I => \N__7447\
        );

    \I__1581\ : CascadeMux
    port map (
            O => \N__7450\,
            I => \N__7444\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__7447\,
            I => \N__7436\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7444\,
            I => \N__7433\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__7443\,
            I => \N__7426\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__7442\,
            I => \N__7422\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__7441\,
            I => \N__7419\
        );

    \I__1575\ : InMux
    port map (
            O => \N__7440\,
            I => \N__7412\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7439\,
            I => \N__7412\
        );

    \I__1573\ : Span4Mux_h
    port map (
            O => \N__7436\,
            I => \N__7409\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__7433\,
            I => \N__7406\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7432\,
            I => \N__7399\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7431\,
            I => \N__7399\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7430\,
            I => \N__7399\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7429\,
            I => \N__7396\
        );

    \I__1567\ : InMux
    port map (
            O => \N__7426\,
            I => \N__7391\
        );

    \I__1566\ : InMux
    port map (
            O => \N__7425\,
            I => \N__7391\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7422\,
            I => \N__7388\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7385\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7418\,
            I => \N__7382\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7417\,
            I => \N__7379\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7412\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__7409\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__7406\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7399\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7396\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7391\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7388\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__7385\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__7382\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7379\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7358\,
            I => \N__7351\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7357\,
            I => \N__7344\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7356\,
            I => \N__7344\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7355\,
            I => \N__7344\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7354\,
            I => \N__7341\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__7351\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7344\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7341\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7334\,
            I => \N__7323\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7323\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7320\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__7331\,
            I => \N__7315\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__7330\,
            I => \N__7308\
        );

    \I__1538\ : InMux
    port map (
            O => \N__7329\,
            I => \N__7300\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7328\,
            I => \N__7300\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__7323\,
            I => \N__7288\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__7320\,
            I => \N__7288\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7285\
        );

    \I__1533\ : InMux
    port map (
            O => \N__7318\,
            I => \N__7280\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7315\,
            I => \N__7280\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7314\,
            I => \N__7274\
        );

    \I__1530\ : InMux
    port map (
            O => \N__7313\,
            I => \N__7274\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7312\,
            I => \N__7267\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7311\,
            I => \N__7267\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7308\,
            I => \N__7267\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7307\,
            I => \N__7262\
        );

    \I__1525\ : InMux
    port map (
            O => \N__7306\,
            I => \N__7262\
        );

    \I__1524\ : InMux
    port map (
            O => \N__7305\,
            I => \N__7257\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7300\,
            I => \N__7253\
        );

    \I__1522\ : InMux
    port map (
            O => \N__7299\,
            I => \N__7248\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7298\,
            I => \N__7248\
        );

    \I__1520\ : InMux
    port map (
            O => \N__7297\,
            I => \N__7241\
        );

    \I__1519\ : InMux
    port map (
            O => \N__7296\,
            I => \N__7241\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7295\,
            I => \N__7241\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7236\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7293\,
            I => \N__7236\
        );

    \I__1515\ : Span4Mux_v
    port map (
            O => \N__7288\,
            I => \N__7233\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__7285\,
            I => \N__7228\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7280\,
            I => \N__7228\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7279\,
            I => \N__7225\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7274\,
            I => \N__7222\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7267\,
            I => \N__7217\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__7262\,
            I => \N__7217\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7261\,
            I => \N__7214\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7260\,
            I => \N__7211\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7257\,
            I => \N__7208\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7256\,
            I => \N__7205\
        );

    \I__1504\ : Span4Mux_v
    port map (
            O => \N__7253\,
            I => \N__7200\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7248\,
            I => \N__7200\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7241\,
            I => \N__7195\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7236\,
            I => \N__7195\
        );

    \I__1500\ : Span4Mux_v
    port map (
            O => \N__7233\,
            I => \N__7188\
        );

    \I__1499\ : Span4Mux_v
    port map (
            O => \N__7228\,
            I => \N__7188\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7225\,
            I => \N__7188\
        );

    \I__1497\ : Span4Mux_h
    port map (
            O => \N__7222\,
            I => \N__7179\
        );

    \I__1496\ : Span4Mux_v
    port map (
            O => \N__7217\,
            I => \N__7179\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7214\,
            I => \N__7179\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7211\,
            I => \N__7179\
        );

    \I__1493\ : Span4Mux_v
    port map (
            O => \N__7208\,
            I => \N__7174\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7205\,
            I => \N__7174\
        );

    \I__1491\ : Span4Mux_v
    port map (
            O => \N__7200\,
            I => \N__7168\
        );

    \I__1490\ : Span4Mux_v
    port map (
            O => \N__7195\,
            I => \N__7168\
        );

    \I__1489\ : Span4Mux_h
    port map (
            O => \N__7188\,
            I => \N__7163\
        );

    \I__1488\ : Span4Mux_v
    port map (
            O => \N__7179\,
            I => \N__7163\
        );

    \I__1487\ : Sp12to4
    port map (
            O => \N__7174\,
            I => \N__7160\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7157\
        );

    \I__1485\ : Sp12to4
    port map (
            O => \N__7168\,
            I => \N__7154\
        );

    \I__1484\ : Sp12to4
    port map (
            O => \N__7163\,
            I => \N__7147\
        );

    \I__1483\ : Span12Mux_v
    port map (
            O => \N__7160\,
            I => \N__7147\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7157\,
            I => \N__7147\
        );

    \I__1481\ : Span12Mux_h
    port map (
            O => \N__7154\,
            I => \N__7144\
        );

    \I__1480\ : Span12Mux_h
    port map (
            O => \N__7147\,
            I => \N__7141\
        );

    \I__1479\ : Odrv12
    port map (
            O => \N__7144\,
            I => \RESETn_c\
        );

    \I__1478\ : Odrv12
    port map (
            O => \N__7141\,
            I => \RESETn_c\
        );

    \I__1477\ : IoInMux
    port map (
            O => \N__7136\,
            I => \N__7133\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7133\,
            I => \N__7130\
        );

    \I__1475\ : Span12Mux_s5_v
    port map (
            O => \N__7130\,
            I => \N__7127\
        );

    \I__1474\ : Odrv12
    port map (
            O => \N__7127\,
            I => \RESETn_c_i\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7124\,
            I => \N__7121\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__7121\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7115\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7115\,
            I => \N__7112\
        );

    \I__1469\ : Span4Mux_h
    port map (
            O => \N__7112\,
            I => \N__7109\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__7109\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7106\,
            I => \N__7103\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7103\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7095\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7099\,
            I => \N__7090\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7098\,
            I => \N__7090\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7095\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__7090\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__7085\,
            I => \N__7082\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7082\,
            I => \N__7079\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7079\,
            I => \N__7076\
        );

    \I__1457\ : Span12Mux_v
    port map (
            O => \N__7076\,
            I => \N__7071\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7075\,
            I => \N__7068\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7074\,
            I => \N__7065\
        );

    \I__1454\ : Odrv12
    port map (
            O => \N__7071\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7068\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__7065\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7058\,
            I => \N__7055\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7055\,
            I => \U712_REG_SM.N_159_0\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7052\,
            I => \N__7049\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7049\,
            I => \N__7045\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7048\,
            I => \N__7042\
        );

    \I__1446\ : Span4Mux_h
    port map (
            O => \N__7045\,
            I => \N__7039\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7042\,
            I => \N__7036\
        );

    \I__1444\ : Odrv4
    port map (
            O => \N__7039\,
            I => \REG_TACK\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__7036\,
            I => \REG_TACK\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__7031\,
            I => \N__7027\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7030\,
            I => \N__7024\
        );

    \I__1440\ : InMux
    port map (
            O => \N__7027\,
            I => \N__7021\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__7024\,
            I => \N__7018\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__7021\,
            I => \N__7015\
        );

    \I__1437\ : Span12Mux_v
    port map (
            O => \N__7018\,
            I => \N__7012\
        );

    \I__1436\ : Odrv12
    port map (
            O => \N__7015\,
            I => \CPU_TACKm\
        );

    \I__1435\ : Odrv12
    port map (
            O => \N__7012\,
            I => \CPU_TACKm\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7007\,
            I => \N__7000\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7006\,
            I => \N__7000\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7005\,
            I => \N__6997\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__7000\,
            I => \N__6994\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6997\,
            I => \N__6990\
        );

    \I__1429\ : Span4Mux_v
    port map (
            O => \N__6994\,
            I => \N__6987\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6993\,
            I => \N__6984\
        );

    \I__1427\ : Span4Mux_v
    port map (
            O => \N__6990\,
            I => \N__6981\
        );

    \I__1426\ : Span4Mux_v
    port map (
            O => \N__6987\,
            I => \N__6976\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__6984\,
            I => \N__6976\
        );

    \I__1424\ : Sp12to4
    port map (
            O => \N__6981\,
            I => \N__6973\
        );

    \I__1423\ : Span4Mux_h
    port map (
            O => \N__6976\,
            I => \N__6970\
        );

    \I__1422\ : Span12Mux_h
    port map (
            O => \N__6973\,
            I => \N__6965\
        );

    \I__1421\ : Sp12to4
    port map (
            O => \N__6970\,
            I => \N__6965\
        );

    \I__1420\ : Span12Mux_v
    port map (
            O => \N__6965\,
            I => \N__6962\
        );

    \I__1419\ : Odrv12
    port map (
            O => \N__6962\,
            I => \CLK40_OUT_i\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__6959\,
            I => \U712_CYCLE_TERM.N_49_cascade_\
        );

    \I__1417\ : InMux
    port map (
            O => \N__6956\,
            I => \N__6953\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__6953\,
            I => \N__6947\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6952\,
            I => \N__6942\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6951\,
            I => \N__6942\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6950\,
            I => \N__6939\
        );

    \I__1412\ : Span4Mux_v
    port map (
            O => \N__6947\,
            I => \N__6934\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6942\,
            I => \N__6934\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__6939\,
            I => \N__6931\
        );

    \I__1409\ : Odrv4
    port map (
            O => \N__6934\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1408\ : Odrv4
    port map (
            O => \N__6931\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1407\ : InMux
    port map (
            O => \N__6926\,
            I => \N__6923\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__6923\,
            I => \N__6918\
        );

    \I__1405\ : InMux
    port map (
            O => \N__6922\,
            I => \N__6913\
        );

    \I__1404\ : InMux
    port map (
            O => \N__6921\,
            I => \N__6913\
        );

    \I__1403\ : Span4Mux_v
    port map (
            O => \N__6918\,
            I => \N__6909\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__6913\,
            I => \N__6906\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6912\,
            I => \N__6903\
        );

    \I__1400\ : Odrv4
    port map (
            O => \N__6909\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1399\ : Odrv4
    port map (
            O => \N__6906\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6903\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1397\ : InMux
    port map (
            O => \N__6896\,
            I => \N__6891\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6895\,
            I => \N__6885\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6894\,
            I => \N__6885\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6891\,
            I => \N__6881\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6890\,
            I => \N__6878\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__6885\,
            I => \N__6875\
        );

    \I__1391\ : InMux
    port map (
            O => \N__6884\,
            I => \N__6872\
        );

    \I__1390\ : Span4Mux_h
    port map (
            O => \N__6881\,
            I => \N__6866\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__6878\,
            I => \N__6866\
        );

    \I__1388\ : Span4Mux_v
    port map (
            O => \N__6875\,
            I => \N__6861\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__6872\,
            I => \N__6861\
        );

    \I__1386\ : InMux
    port map (
            O => \N__6871\,
            I => \N__6858\
        );

    \I__1385\ : Span4Mux_v
    port map (
            O => \N__6866\,
            I => \N__6853\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__6861\,
            I => \N__6850\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__6858\,
            I => \N__6847\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6857\,
            I => \N__6844\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6856\,
            I => \N__6841\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__6853\,
            I => \DMA_CYCLEm\
        );

    \I__1379\ : Odrv4
    port map (
            O => \N__6850\,
            I => \DMA_CYCLEm\
        );

    \I__1378\ : Odrv4
    port map (
            O => \N__6847\,
            I => \DMA_CYCLEm\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__6844\,
            I => \DMA_CYCLEm\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__6841\,
            I => \DMA_CYCLEm\
        );

    \I__1375\ : CascadeMux
    port map (
            O => \N__6830\,
            I => \N__6826\
        );

    \I__1374\ : InMux
    port map (
            O => \N__6829\,
            I => \N__6823\
        );

    \I__1373\ : InMux
    port map (
            O => \N__6826\,
            I => \N__6820\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__6823\,
            I => \N__6816\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__6820\,
            I => \N__6813\
        );

    \I__1370\ : InMux
    port map (
            O => \N__6819\,
            I => \N__6810\
        );

    \I__1369\ : Span12Mux_v
    port map (
            O => \N__6816\,
            I => \N__6806\
        );

    \I__1368\ : Span4Mux_h
    port map (
            O => \N__6813\,
            I => \N__6801\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__6810\,
            I => \N__6801\
        );

    \I__1366\ : InMux
    port map (
            O => \N__6809\,
            I => \N__6798\
        );

    \I__1365\ : Odrv12
    port map (
            O => \N__6806\,
            I => \REG_CYCLEm\
        );

    \I__1364\ : Odrv4
    port map (
            O => \N__6801\,
            I => \REG_CYCLEm\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__6798\,
            I => \REG_CYCLEm\
        );

    \I__1362\ : IoInMux
    port map (
            O => \N__6791\,
            I => \N__6788\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6788\,
            I => \N__6785\
        );

    \I__1360\ : IoSpan4Mux
    port map (
            O => \N__6785\,
            I => \N__6782\
        );

    \I__1359\ : Sp12to4
    port map (
            O => \N__6782\,
            I => \N__6779\
        );

    \I__1358\ : Span12Mux_s7_h
    port map (
            O => \N__6779\,
            I => \N__6776\
        );

    \I__1357\ : Span12Mux_v
    port map (
            O => \N__6776\,
            I => \N__6773\
        );

    \I__1356\ : Odrv12
    port map (
            O => \N__6773\,
            I => \DRDENn_c\
        );

    \I__1355\ : IoInMux
    port map (
            O => \N__6770\,
            I => \N__6767\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6767\,
            I => \N__6764\
        );

    \I__1353\ : Span4Mux_s3_v
    port map (
            O => \N__6764\,
            I => \N__6761\
        );

    \I__1352\ : Span4Mux_h
    port map (
            O => \N__6761\,
            I => \N__6758\
        );

    \I__1351\ : Odrv4
    port map (
            O => \N__6758\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1350\ : IoInMux
    port map (
            O => \N__6755\,
            I => \N__6752\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6752\,
            I => \N__6749\
        );

    \I__1348\ : Span4Mux_s1_v
    port map (
            O => \N__6749\,
            I => \N__6746\
        );

    \I__1347\ : Span4Mux_v
    port map (
            O => \N__6746\,
            I => \N__6743\
        );

    \I__1346\ : Span4Mux_v
    port map (
            O => \N__6743\,
            I => \N__6740\
        );

    \I__1345\ : Odrv4
    port map (
            O => \N__6740\,
            I => \CMA_c_2\
        );

    \I__1344\ : IoInMux
    port map (
            O => \N__6737\,
            I => \N__6734\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__6734\,
            I => \N__6731\
        );

    \I__1342\ : IoSpan4Mux
    port map (
            O => \N__6731\,
            I => \N__6728\
        );

    \I__1341\ : IoSpan4Mux
    port map (
            O => \N__6728\,
            I => \N__6725\
        );

    \I__1340\ : Sp12to4
    port map (
            O => \N__6725\,
            I => \N__6722\
        );

    \I__1339\ : Span12Mux_s7_h
    port map (
            O => \N__6722\,
            I => \N__6719\
        );

    \I__1338\ : Odrv12
    port map (
            O => \N__6719\,
            I => \CMA_c_5\
        );

    \I__1337\ : InMux
    port map (
            O => \N__6716\,
            I => \N__6712\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6715\,
            I => \N__6709\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__6712\,
            I => \U712_CHIP_RAM.N_124\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__6709\,
            I => \U712_CHIP_RAM.N_124\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__6704\,
            I => \U712_CHIP_RAM.N_96_cascade_\
        );

    \I__1332\ : InMux
    port map (
            O => \N__6701\,
            I => \N__6696\
        );

    \I__1331\ : InMux
    port map (
            O => \N__6700\,
            I => \N__6690\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6699\,
            I => \N__6687\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6696\,
            I => \N__6684\
        );

    \I__1328\ : InMux
    port map (
            O => \N__6695\,
            I => \N__6681\
        );

    \I__1327\ : InMux
    port map (
            O => \N__6694\,
            I => \N__6676\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6693\,
            I => \N__6676\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__6690\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6687\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\
        );

    \I__1323\ : Odrv12
    port map (
            O => \N__6684\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6681\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6676\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__6665\,
            I => \N__6662\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6662\,
            I => \N__6656\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6656\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6656\,
            I => \U712_CHIP_RAM.N_72\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__6653\,
            I => \N__6649\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6652\,
            I => \N__6646\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6649\,
            I => \N__6642\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6646\,
            I => \N__6639\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6645\,
            I => \N__6636\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__6642\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1310\ : Odrv4
    port map (
            O => \N__6639\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6636\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1308\ : CascadeMux
    port map (
            O => \N__6629\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_0_cascade_\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__6626\,
            I => \N__6623\
        );

    \I__1306\ : InMux
    port map (
            O => \N__6623\,
            I => \N__6620\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6620\,
            I => \N__6616\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__6619\,
            I => \N__6613\
        );

    \I__1303\ : Span4Mux_v
    port map (
            O => \N__6616\,
            I => \N__6607\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6604\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6612\,
            I => \N__6601\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6611\,
            I => \N__6596\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6596\
        );

    \I__1298\ : Span4Mux_h
    port map (
            O => \N__6607\,
            I => \N__6582\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6604\,
            I => \N__6582\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__6601\,
            I => \N__6582\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__6596\,
            I => \N__6582\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6573\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6568\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6593\,
            I => \N__6568\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6592\,
            I => \N__6563\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6591\,
            I => \N__6563\
        );

    \I__1289\ : Span4Mux_v
    port map (
            O => \N__6582\,
            I => \N__6560\
        );

    \I__1288\ : InMux
    port map (
            O => \N__6581\,
            I => \N__6553\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6580\,
            I => \N__6553\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6579\,
            I => \N__6553\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6578\,
            I => \N__6546\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6546\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6546\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__6573\,
            I => \N__6543\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6568\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__6563\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1279\ : Odrv4
    port map (
            O => \N__6560\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__6553\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6546\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1276\ : Odrv4
    port map (
            O => \N__6543\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6530\,
            I => \N__6523\
        );

    \I__1274\ : CascadeMux
    port map (
            O => \N__6529\,
            I => \N__6520\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6528\,
            I => \N__6516\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__6527\,
            I => \N__6508\
        );

    \I__1271\ : InMux
    port map (
            O => \N__6526\,
            I => \N__6500\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__6523\,
            I => \N__6497\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6520\,
            I => \N__6494\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6491\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__6516\,
            I => \N__6488\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6515\,
            I => \N__6479\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6514\,
            I => \N__6479\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6513\,
            I => \N__6479\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6512\,
            I => \N__6479\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6511\,
            I => \N__6476\
        );

    \I__1261\ : InMux
    port map (
            O => \N__6508\,
            I => \N__6469\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6507\,
            I => \N__6469\
        );

    \I__1259\ : InMux
    port map (
            O => \N__6506\,
            I => \N__6469\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6505\,
            I => \N__6462\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6504\,
            I => \N__6462\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6462\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__6500\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__6497\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__6494\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__6491\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1251\ : Odrv12
    port map (
            O => \N__6488\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6479\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__6476\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6469\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6462\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__6443\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_3_cascade_\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__6440\,
            I => \N__6432\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6439\,
            I => \N__6429\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6438\,
            I => \N__6425\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6437\,
            I => \N__6422\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6436\,
            I => \N__6419\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6435\,
            I => \N__6416\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6432\,
            I => \N__6412\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6429\,
            I => \N__6409\
        );

    \I__1237\ : InMux
    port map (
            O => \N__6428\,
            I => \N__6406\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6425\,
            I => \N__6401\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6422\,
            I => \N__6401\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6419\,
            I => \N__6396\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6416\,
            I => \N__6396\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6415\,
            I => \N__6393\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__6412\,
            I => \U712_CHIP_RAM.N_65\
        );

    \I__1230\ : Odrv4
    port map (
            O => \N__6409\,
            I => \U712_CHIP_RAM.N_65\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__6406\,
            I => \U712_CHIP_RAM.N_65\
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__6401\,
            I => \U712_CHIP_RAM.N_65\
        );

    \I__1227\ : Odrv4
    port map (
            O => \N__6396\,
            I => \U712_CHIP_RAM.N_65\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6393\,
            I => \U712_CHIP_RAM.N_65\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__6380\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_cascade_\
        );

    \I__1224\ : CEMux
    port map (
            O => \N__6377\,
            I => \N__6374\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6374\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_1\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6367\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6370\,
            I => \N__6362\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6367\,
            I => \N__6359\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6366\,
            I => \N__6356\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6365\,
            I => \N__6353\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__6362\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__6359\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__6356\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6353\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__6344\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__6341\,
            I => \N__6336\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__6340\,
            I => \N__6333\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__6339\,
            I => \N__6330\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6324\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6333\,
            I => \N__6324\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6330\,
            I => \N__6321\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6329\,
            I => \N__6318\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6324\,
            I => \N__6313\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__6321\,
            I => \N__6313\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6318\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1202\ : Odrv4
    port map (
            O => \N__6313\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6308\,
            I => \N__6305\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6305\,
            I => \N__6301\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6304\,
            I => \N__6298\
        );

    \I__1198\ : Odrv4
    port map (
            O => \N__6301\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6298\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6286\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6292\,
            I => \N__6286\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6283\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6286\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6283\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6278\,
            I => \N__6275\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__6275\,
            I => \U712_CHIP_RAM.un6_CPU_CYCLE_START\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6272\,
            I => \N__6269\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6269\,
            I => \N__6266\
        );

    \I__1187\ : Span4Mux_h
    port map (
            O => \N__6266\,
            I => \N__6260\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6265\,
            I => \N__6257\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6264\,
            I => \N__6254\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6263\,
            I => \N__6251\
        );

    \I__1183\ : Odrv4
    port map (
            O => \N__6260\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6257\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6254\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6251\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6242\,
            I => \N__6236\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6233\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6240\,
            I => \N__6230\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6239\,
            I => \N__6227\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6236\,
            I => \U712_CHIP_RAM.N_52\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6233\,
            I => \U712_CHIP_RAM.N_52\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__6230\,
            I => \U712_CHIP_RAM.N_52\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6227\,
            I => \U712_CHIP_RAM.N_52\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6218\,
            I => \N__6215\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6215\,
            I => \N__6212\
        );

    \I__1169\ : Odrv4
    port map (
            O => \N__6212\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER35\
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__6209\,
            I => \U712_CHIP_RAM.N_46_cascade_\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__6206\,
            I => \N__6203\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6199\
        );

    \I__1165\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6196\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__6199\,
            I => \N__6192\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6196\,
            I => \N__6189\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6186\
        );

    \I__1161\ : Span4Mux_h
    port map (
            O => \N__6192\,
            I => \N__6183\
        );

    \I__1160\ : Odrv4
    port map (
            O => \N__6189\,
            I => \U712_CHIP_RAM.N_116\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6186\,
            I => \U712_CHIP_RAM.N_116\
        );

    \I__1158\ : Odrv4
    port map (
            O => \N__6183\,
            I => \U712_CHIP_RAM.N_116\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__6176\,
            I => \U712_CHIP_RAM.N_116_cascade_\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__6173\,
            I => \N__6168\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6172\,
            I => \N__6165\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6162\
        );

    \I__1153\ : InMux
    port map (
            O => \N__6168\,
            I => \N__6159\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6165\,
            I => \N__6156\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__6162\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER39\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6159\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER39\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__6156\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER39\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6149\,
            I => \N__6141\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6148\,
            I => \N__6141\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6147\,
            I => \N__6130\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6146\,
            I => \N__6130\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6141\,
            I => \N__6127\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6124\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6139\,
            I => \N__6121\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6138\,
            I => \N__6114\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6137\,
            I => \N__6114\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6136\,
            I => \N__6114\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6135\,
            I => \N__6111\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6130\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1136\ : Odrv4
    port map (
            O => \N__6127\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6124\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6121\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6114\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6111\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__6098\,
            I => \N__6093\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6090\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6096\,
            I => \N__6084\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6081\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__6090\,
            I => \N__6078\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6089\,
            I => \N__6073\
        );

    \I__1125\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6073\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6087\,
            I => \N__6070\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6084\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6081\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1121\ : Odrv4
    port map (
            O => \N__6078\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__6073\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6070\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__6059\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_1_1_cascade_\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6056\,
            I => \N__6051\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6055\,
            I => \N__6048\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6054\,
            I => \N__6045\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6051\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__6048\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6045\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6035\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6035\,
            I => \U712_CHIP_RAM.N_96\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__6032\,
            I => \N__6028\
        );

    \I__1108\ : InMux
    port map (
            O => \N__6031\,
            I => \N__6025\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6022\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6025\,
            I => \N__6017\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6022\,
            I => \N__6017\
        );

    \I__1104\ : Sp12to4
    port map (
            O => \N__6017\,
            I => \N__6013\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6016\,
            I => \N__6010\
        );

    \I__1102\ : Odrv12
    port map (
            O => \N__6013\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__6010\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__6005\,
            I => \N__6001\
        );

    \I__1099\ : InMux
    port map (
            O => \N__6004\,
            I => \N__5998\
        );

    \I__1098\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5995\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5998\,
            I => \N__5992\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5995\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1095\ : Odrv4
    port map (
            O => \N__5992\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5987\,
            I => \N__5983\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5986\,
            I => \N__5980\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__5983\,
            I => \U712_REG_SM.C1_SYNC_RNIPBP14Z0Z_2\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5980\,
            I => \U712_REG_SM.C1_SYNC_RNIPBP14Z0Z_2\
        );

    \I__1090\ : CEMux
    port map (
            O => \N__5975\,
            I => \N__5972\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5972\,
            I => \U712_REG_SM.N_180_0\
        );

    \I__1088\ : IoInMux
    port map (
            O => \N__5969\,
            I => \N__5966\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__5966\,
            I => \N__5963\
        );

    \I__1086\ : Span4Mux_s1_v
    port map (
            O => \N__5963\,
            I => \N__5960\
        );

    \I__1085\ : Span4Mux_v
    port map (
            O => \N__5960\,
            I => \N__5957\
        );

    \I__1084\ : Span4Mux_v
    port map (
            O => \N__5957\,
            I => \N__5954\
        );

    \I__1083\ : Span4Mux_h
    port map (
            O => \N__5954\,
            I => \N__5951\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__5951\,
            I => \CMA_c_0\
        );

    \I__1081\ : IoInMux
    port map (
            O => \N__5948\,
            I => \N__5945\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__5945\,
            I => \N__5942\
        );

    \I__1079\ : IoSpan4Mux
    port map (
            O => \N__5942\,
            I => \N__5939\
        );

    \I__1078\ : IoSpan4Mux
    port map (
            O => \N__5939\,
            I => \N__5936\
        );

    \I__1077\ : Sp12to4
    port map (
            O => \N__5936\,
            I => \N__5933\
        );

    \I__1076\ : Span12Mux_s7_h
    port map (
            O => \N__5933\,
            I => \N__5930\
        );

    \I__1075\ : Odrv12
    port map (
            O => \N__5930\,
            I => \CMA_c_4\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5924\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__5924\,
            I => \N__5921\
        );

    \I__1072\ : Sp12to4
    port map (
            O => \N__5921\,
            I => \N__5918\
        );

    \I__1071\ : Span12Mux_v
    port map (
            O => \N__5918\,
            I => \N__5915\
        );

    \I__1070\ : Span12Mux_h
    port map (
            O => \N__5915\,
            I => \N__5912\
        );

    \I__1069\ : Span12Mux_v
    port map (
            O => \N__5912\,
            I => \N__5909\
        );

    \I__1068\ : Odrv12
    port map (
            O => \N__5909\,
            I => \A_c_2\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__5906\,
            I => \N__5903\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5903\,
            I => \N__5900\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5900\,
            I => \N__5897\
        );

    \I__1064\ : Sp12to4
    port map (
            O => \N__5897\,
            I => \N__5894\
        );

    \I__1063\ : Span12Mux_v
    port map (
            O => \N__5894\,
            I => \N__5891\
        );

    \I__1062\ : Span12Mux_h
    port map (
            O => \N__5891\,
            I => \N__5888\
        );

    \I__1061\ : Odrv12
    port map (
            O => \N__5888\,
            I => \A_c_9\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5885\,
            I => \N__5882\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5882\,
            I => \U712_CHIP_RAM.N_31\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5879\,
            I => \N__5876\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__5876\,
            I => \N__5873\
        );

    \I__1056\ : Span12Mux_h
    port map (
            O => \N__5873\,
            I => \N__5870\
        );

    \I__1055\ : Odrv12
    port map (
            O => \N__5870\,
            I => \A_c_13\
        );

    \I__1054\ : CascadeMux
    port map (
            O => \N__5867\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_4_cascade_\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5864\,
            I => \N__5861\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5861\,
            I => \N__5858\
        );

    \I__1051\ : Span4Mux_v
    port map (
            O => \N__5858\,
            I => \N__5855\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__5855\,
            I => \N__5852\
        );

    \I__1049\ : Sp12to4
    port map (
            O => \N__5852\,
            I => \N__5849\
        );

    \I__1048\ : Span12Mux_h
    port map (
            O => \N__5849\,
            I => \N__5846\
        );

    \I__1047\ : Odrv12
    port map (
            O => \N__5846\,
            I => \A_c_6\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5843\,
            I => \N__5840\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5840\,
            I => \U712_CHIP_RAM.N_35\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5834\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5834\,
            I => \N__5830\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5833\,
            I => \N__5827\
        );

    \I__1041\ : Span4Mux_v
    port map (
            O => \N__5830\,
            I => \N__5824\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5827\,
            I => \N__5821\
        );

    \I__1039\ : Span4Mux_h
    port map (
            O => \N__5824\,
            I => \N__5816\
        );

    \I__1038\ : Span4Mux_v
    port map (
            O => \N__5821\,
            I => \N__5816\
        );

    \I__1037\ : Span4Mux_h
    port map (
            O => \N__5816\,
            I => \N__5813\
        );

    \I__1036\ : Sp12to4
    port map (
            O => \N__5813\,
            I => \N__5810\
        );

    \I__1035\ : Span12Mux_v
    port map (
            O => \N__5810\,
            I => \N__5807\
        );

    \I__1034\ : Odrv12
    port map (
            O => \N__5807\,
            I => \AWEn_c\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__5804\,
            I => \N__5801\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5797\
        );

    \I__1031\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5792\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5797\,
            I => \N__5789\
        );

    \I__1029\ : InMux
    port map (
            O => \N__5796\,
            I => \N__5785\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5795\,
            I => \N__5782\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5792\,
            I => \N__5779\
        );

    \I__1026\ : Span4Mux_h
    port map (
            O => \N__5789\,
            I => \N__5776\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5788\,
            I => \N__5773\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__5785\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__5782\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1022\ : Odrv4
    port map (
            O => \N__5779\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__5776\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5773\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5762\,
            I => \N__5756\
        );

    \I__1018\ : InMux
    port map (
            O => \N__5761\,
            I => \N__5753\
        );

    \I__1017\ : InMux
    port map (
            O => \N__5760\,
            I => \N__5750\
        );

    \I__1016\ : InMux
    port map (
            O => \N__5759\,
            I => \N__5747\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5756\,
            I => \N__5743\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5753\,
            I => \N__5740\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__5750\,
            I => \N__5735\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5747\,
            I => \N__5735\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5746\,
            I => \N__5732\
        );

    \I__1010\ : Span4Mux_v
    port map (
            O => \N__5743\,
            I => \N__5729\
        );

    \I__1009\ : Span4Mux_v
    port map (
            O => \N__5740\,
            I => \N__5726\
        );

    \I__1008\ : Span4Mux_v
    port map (
            O => \N__5735\,
            I => \N__5723\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__5732\,
            I => \N__5720\
        );

    \I__1006\ : Sp12to4
    port map (
            O => \N__5729\,
            I => \N__5713\
        );

    \I__1005\ : Sp12to4
    port map (
            O => \N__5726\,
            I => \N__5713\
        );

    \I__1004\ : Sp12to4
    port map (
            O => \N__5723\,
            I => \N__5713\
        );

    \I__1003\ : Span12Mux_v
    port map (
            O => \N__5720\,
            I => \N__5710\
        );

    \I__1002\ : Span12Mux_h
    port map (
            O => \N__5713\,
            I => \N__5707\
        );

    \I__1001\ : Span12Mux_h
    port map (
            O => \N__5710\,
            I => \N__5704\
        );

    \I__1000\ : Span12Mux_v
    port map (
            O => \N__5707\,
            I => \N__5701\
        );

    \I__999\ : Odrv12
    port map (
            O => \N__5704\,
            I => \RnW_c\
        );

    \I__998\ : Odrv12
    port map (
            O => \N__5701\,
            I => \RnW_c\
        );

    \I__997\ : InMux
    port map (
            O => \N__5696\,
            I => \N__5693\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5693\,
            I => \N__5690\
        );

    \I__995\ : Span4Mux_h
    port map (
            O => \N__5690\,
            I => \N__5687\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__5687\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_0\
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__5684\,
            I => \U712_CHIP_RAM.N_52_cascade_\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__5681\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0_cascade_\
        );

    \I__991\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5673\
        );

    \I__990\ : InMux
    port map (
            O => \N__5677\,
            I => \N__5670\
        );

    \I__989\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5667\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5673\,
            I => \N__5664\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__5670\,
            I => \N__5661\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5667\,
            I => \U712_CHIP_RAM.N_61\
        );

    \I__985\ : Odrv12
    port map (
            O => \N__5664\,
            I => \U712_CHIP_RAM.N_61\
        );

    \I__984\ : Odrv4
    port map (
            O => \N__5661\,
            I => \U712_CHIP_RAM.N_61\
        );

    \I__983\ : CascadeMux
    port map (
            O => \N__5654\,
            I => \U712_CHIP_RAM.N_90_cascade_\
        );

    \I__982\ : InMux
    port map (
            O => \N__5651\,
            I => \N__5648\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5648\,
            I => \U712_CHIP_RAM.N_69\
        );

    \I__980\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5640\
        );

    \I__979\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5635\
        );

    \I__978\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5635\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5640\,
            I => \U712_CHIP_RAM.N_57\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5635\,
            I => \U712_CHIP_RAM.N_57\
        );

    \I__975\ : IoInMux
    port map (
            O => \N__5630\,
            I => \N__5627\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__5627\,
            I => \N__5624\
        );

    \I__973\ : Span4Mux_s3_h
    port map (
            O => \N__5624\,
            I => \N__5621\
        );

    \I__972\ : Span4Mux_v
    port map (
            O => \N__5621\,
            I => \N__5618\
        );

    \I__971\ : Span4Mux_v
    port map (
            O => \N__5618\,
            I => \N__5615\
        );

    \I__970\ : Span4Mux_h
    port map (
            O => \N__5615\,
            I => \N__5612\
        );

    \I__969\ : Sp12to4
    port map (
            O => \N__5612\,
            I => \N__5608\
        );

    \I__968\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5605\
        );

    \I__967\ : Odrv12
    port map (
            O => \N__5608\,
            I => \CLK_EN_c\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5605\,
            I => \CLK_EN_c\
        );

    \I__965\ : InMux
    port map (
            O => \N__5600\,
            I => \N__5594\
        );

    \I__964\ : InMux
    port map (
            O => \N__5599\,
            I => \N__5594\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__5594\,
            I => \N__5591\
        );

    \I__962\ : Span4Mux_h
    port map (
            O => \N__5591\,
            I => \N__5588\
        );

    \I__961\ : Odrv4
    port map (
            O => \N__5588\,
            I => \U712_CHIP_RAM.DMA_CYCLE_7\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__5585\,
            I => \N__5582\
        );

    \I__959\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5577\
        );

    \I__958\ : InMux
    port map (
            O => \N__5581\,
            I => \N__5574\
        );

    \I__957\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5571\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__5577\,
            I => \U712_REG_SM.N_151_0\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5574\,
            I => \U712_REG_SM.N_151_0\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5571\,
            I => \U712_REG_SM.N_151_0\
        );

    \I__953\ : InMux
    port map (
            O => \N__5564\,
            I => \N__5560\
        );

    \I__952\ : InMux
    port map (
            O => \N__5563\,
            I => \N__5556\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__5560\,
            I => \N__5553\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__5559\,
            I => \N__5550\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5556\,
            I => \N__5547\
        );

    \I__948\ : Span4Mux_v
    port map (
            O => \N__5553\,
            I => \N__5544\
        );

    \I__947\ : InMux
    port map (
            O => \N__5550\,
            I => \N__5541\
        );

    \I__946\ : Odrv12
    port map (
            O => \N__5547\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__945\ : Odrv4
    port map (
            O => \N__5544\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5541\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__943\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5530\
        );

    \I__942\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5527\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5530\,
            I => \N__5524\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5527\,
            I => \N__5519\
        );

    \I__939\ : Span4Mux_v
    port map (
            O => \N__5524\,
            I => \N__5516\
        );

    \I__938\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5511\
        );

    \I__937\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5511\
        );

    \I__936\ : Odrv12
    port map (
            O => \N__5519\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__935\ : Odrv4
    port map (
            O => \N__5516\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5511\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__5504\,
            I => \U712_REG_SM.N_159_0_cascade_\
        );

    \I__932\ : InMux
    port map (
            O => \N__5501\,
            I => \N__5498\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5498\,
            I => \U712_REG_SM.N_165\
        );

    \I__930\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5492\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5492\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0\
        );

    \I__928\ : CascadeMux
    port map (
            O => \N__5489\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_0_cascade_\
        );

    \I__927\ : InMux
    port map (
            O => \N__5486\,
            I => \N__5481\
        );

    \I__926\ : InMux
    port map (
            O => \N__5485\,
            I => \N__5478\
        );

    \I__925\ : InMux
    port map (
            O => \N__5484\,
            I => \N__5475\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5481\,
            I => \U712_CHIP_RAM.N_68\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5478\,
            I => \U712_CHIP_RAM.N_68\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__5475\,
            I => \U712_CHIP_RAM.N_68\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__5468\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_1_1_cascade_\
        );

    \I__920\ : InMux
    port map (
            O => \N__5465\,
            I => \N__5462\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__5462\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_0_1\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__5459\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_cascade_\
        );

    \I__917\ : InMux
    port map (
            O => \N__5456\,
            I => \N__5450\
        );

    \I__916\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5450\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__5450\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__914\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5444\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5444\,
            I => \N__5441\
        );

    \I__912\ : Span4Mux_v
    port map (
            O => \N__5441\,
            I => \N__5438\
        );

    \I__911\ : Odrv4
    port map (
            O => \N__5438\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__5435\,
            I => \U712_CHIP_RAM.N_58_cascade_\
        );

    \I__909\ : CascadeMux
    port map (
            O => \N__5432\,
            I => \U712_CHIP_RAM.N_97_cascade_\
        );

    \I__908\ : InMux
    port map (
            O => \N__5429\,
            I => \N__5423\
        );

    \I__907\ : InMux
    port map (
            O => \N__5428\,
            I => \N__5420\
        );

    \I__906\ : InMux
    port map (
            O => \N__5427\,
            I => \N__5415\
        );

    \I__905\ : InMux
    port map (
            O => \N__5426\,
            I => \N__5415\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5423\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5420\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5415\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__901\ : InMux
    port map (
            O => \N__5408\,
            I => \N__5404\
        );

    \I__900\ : InMux
    port map (
            O => \N__5407\,
            I => \N__5401\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__5404\,
            I => \N__5398\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__5401\,
            I => \N__5395\
        );

    \I__897\ : Span4Mux_v
    port map (
            O => \N__5398\,
            I => \N__5391\
        );

    \I__896\ : Span4Mux_v
    port map (
            O => \N__5395\,
            I => \N__5388\
        );

    \I__895\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5385\
        );

    \I__894\ : Sp12to4
    port map (
            O => \N__5391\,
            I => \N__5378\
        );

    \I__893\ : Sp12to4
    port map (
            O => \N__5388\,
            I => \N__5378\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5385\,
            I => \N__5378\
        );

    \I__891\ : Span12Mux_h
    port map (
            O => \N__5378\,
            I => \N__5375\
        );

    \I__890\ : Span12Mux_v
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__889\ : Odrv12
    port map (
            O => \N__5372\,
            I => \TSn_c\
        );

    \I__888\ : InMux
    port map (
            O => \N__5369\,
            I => \N__5366\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__886\ : Span4Mux_v
    port map (
            O => \N__5363\,
            I => \N__5360\
        );

    \I__885\ : Span4Mux_h
    port map (
            O => \N__5360\,
            I => \N__5356\
        );

    \I__884\ : IoInMux
    port map (
            O => \N__5359\,
            I => \N__5353\
        );

    \I__883\ : Sp12to4
    port map (
            O => \N__5356\,
            I => \N__5350\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__5353\,
            I => \N__5347\
        );

    \I__881\ : Span12Mux_v
    port map (
            O => \N__5350\,
            I => \N__5344\
        );

    \I__880\ : IoSpan4Mux
    port map (
            O => \N__5347\,
            I => \N__5341\
        );

    \I__879\ : Odrv12
    port map (
            O => \N__5344\,
            I => \RAMENn_c\
        );

    \I__878\ : Odrv4
    port map (
            O => \N__5341\,
            I => \RAMENn_c\
        );

    \I__877\ : InMux
    port map (
            O => \N__5336\,
            I => \N__5333\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5333\,
            I => \U712_CHIP_RAM.N_421_tz\
        );

    \I__875\ : InMux
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5327\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1\
        );

    \I__873\ : InMux
    port map (
            O => \N__5324\,
            I => \N__5317\
        );

    \I__872\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5314\
        );

    \I__871\ : InMux
    port map (
            O => \N__5322\,
            I => \N__5309\
        );

    \I__870\ : InMux
    port map (
            O => \N__5321\,
            I => \N__5309\
        );

    \I__869\ : InMux
    port map (
            O => \N__5320\,
            I => \N__5306\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5317\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5314\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5309\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5306\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__864\ : InMux
    port map (
            O => \N__5297\,
            I => \N__5294\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5294\,
            I => \N__5290\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__5293\,
            I => \N__5287\
        );

    \I__861\ : Span4Mux_h
    port map (
            O => \N__5290\,
            I => \N__5282\
        );

    \I__860\ : InMux
    port map (
            O => \N__5287\,
            I => \N__5277\
        );

    \I__859\ : InMux
    port map (
            O => \N__5286\,
            I => \N__5277\
        );

    \I__858\ : InMux
    port map (
            O => \N__5285\,
            I => \N__5274\
        );

    \I__857\ : Odrv4
    port map (
            O => \N__5282\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__5277\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__5274\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__854\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5256\
        );

    \I__853\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5253\
        );

    \I__852\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5250\
        );

    \I__851\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5241\
        );

    \I__850\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5241\
        );

    \I__849\ : InMux
    port map (
            O => \N__5262\,
            I => \N__5241\
        );

    \I__848\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5241\
        );

    \I__847\ : InMux
    port map (
            O => \N__5260\,
            I => \N__5236\
        );

    \I__846\ : InMux
    port map (
            O => \N__5259\,
            I => \N__5236\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5256\,
            I => \N__5233\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5253\,
            I => \N__5230\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__5250\,
            I => \N__5225\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5241\,
            I => \N__5225\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5236\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__5233\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__839\ : Odrv4
    port map (
            O => \N__5230\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__5225\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__5216\,
            I => \N__5211\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__5215\,
            I => \N__5206\
        );

    \I__835\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5203\
        );

    \I__834\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5195\
        );

    \I__833\ : InMux
    port map (
            O => \N__5210\,
            I => \N__5195\
        );

    \I__832\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5195\
        );

    \I__831\ : InMux
    port map (
            O => \N__5206\,
            I => \N__5192\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5203\,
            I => \N__5189\
        );

    \I__829\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5185\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5195\,
            I => \N__5180\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5192\,
            I => \N__5180\
        );

    \I__826\ : Span4Mux_v
    port map (
            O => \N__5189\,
            I => \N__5177\
        );

    \I__825\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5174\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5185\,
            I => \N__5169\
        );

    \I__823\ : Span4Mux_h
    port map (
            O => \N__5180\,
            I => \N__5169\
        );

    \I__822\ : Odrv4
    port map (
            O => \N__5177\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5174\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__5169\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__819\ : InMux
    port map (
            O => \N__5162\,
            I => \N__5159\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5159\,
            I => \N__5155\
        );

    \I__817\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5152\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__5155\,
            I => \U712_REG_SM.N_187\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__5152\,
            I => \U712_REG_SM.N_187\
        );

    \I__814\ : IoInMux
    port map (
            O => \N__5147\,
            I => \N__5144\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5144\,
            I => \N__5140\
        );

    \I__812\ : IoInMux
    port map (
            O => \N__5143\,
            I => \N__5137\
        );

    \I__811\ : Span4Mux_s3_v
    port map (
            O => \N__5140\,
            I => \N__5134\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__5137\,
            I => \N__5131\
        );

    \I__809\ : Span4Mux_h
    port map (
            O => \N__5134\,
            I => \N__5128\
        );

    \I__808\ : Span4Mux_s3_v
    port map (
            O => \N__5131\,
            I => \N__5125\
        );

    \I__807\ : Span4Mux_h
    port map (
            O => \N__5128\,
            I => \N__5122\
        );

    \I__806\ : Span4Mux_h
    port map (
            O => \N__5125\,
            I => \N__5119\
        );

    \I__805\ : Sp12to4
    port map (
            O => \N__5122\,
            I => \N__5116\
        );

    \I__804\ : Sp12to4
    port map (
            O => \N__5119\,
            I => \N__5113\
        );

    \I__803\ : Span12Mux_v
    port map (
            O => \N__5116\,
            I => \N__5108\
        );

    \I__802\ : Span12Mux_v
    port map (
            O => \N__5113\,
            I => \N__5108\
        );

    \I__801\ : Odrv12
    port map (
            O => \N__5108\,
            I => \ASn_c\
        );

    \I__800\ : InMux
    port map (
            O => \N__5105\,
            I => \N__5101\
        );

    \I__799\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5098\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5101\,
            I => \N__5094\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5098\,
            I => \N__5091\
        );

    \I__796\ : InMux
    port map (
            O => \N__5097\,
            I => \N__5088\
        );

    \I__795\ : Odrv4
    port map (
            O => \N__5094\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__794\ : Odrv4
    port map (
            O => \N__5091\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5088\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__792\ : InMux
    port map (
            O => \N__5081\,
            I => \N__5078\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__5078\,
            I => \N__5075\
        );

    \I__790\ : Span4Mux_v
    port map (
            O => \N__5075\,
            I => \N__5071\
        );

    \I__789\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5068\
        );

    \I__788\ : Odrv4
    port map (
            O => \N__5071\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5068\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__786\ : IoInMux
    port map (
            O => \N__5063\,
            I => \N__5060\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5060\,
            I => \N__5057\
        );

    \I__784\ : Span4Mux_s3_v
    port map (
            O => \N__5057\,
            I => \N__5054\
        );

    \I__783\ : Sp12to4
    port map (
            O => \N__5054\,
            I => \N__5051\
        );

    \I__782\ : Span12Mux_h
    port map (
            O => \N__5051\,
            I => \N__5048\
        );

    \I__781\ : Odrv12
    port map (
            O => \N__5048\,
            I => \U712_REG_SM_un1_UDSn_i\
        );

    \I__780\ : IoInMux
    port map (
            O => \N__5045\,
            I => \N__5042\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5042\,
            I => \N__5039\
        );

    \I__778\ : IoSpan4Mux
    port map (
            O => \N__5039\,
            I => \N__5035\
        );

    \I__777\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5032\
        );

    \I__776\ : Span4Mux_s3_v
    port map (
            O => \N__5035\,
            I => \N__5029\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5032\,
            I => \N__5026\
        );

    \I__774\ : Span4Mux_v
    port map (
            O => \N__5029\,
            I => \N__5022\
        );

    \I__773\ : Span4Mux_v
    port map (
            O => \N__5026\,
            I => \N__5019\
        );

    \I__772\ : InMux
    port map (
            O => \N__5025\,
            I => \N__5016\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__5022\,
            I => \DBDIR_c\
        );

    \I__770\ : Odrv4
    port map (
            O => \N__5019\,
            I => \DBDIR_c\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5016\,
            I => \DBDIR_c\
        );

    \I__768\ : IoInMux
    port map (
            O => \N__5009\,
            I => \N__5006\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__5006\,
            I => \N__5003\
        );

    \I__766\ : IoSpan4Mux
    port map (
            O => \N__5003\,
            I => \N__5000\
        );

    \I__765\ : Span4Mux_s2_h
    port map (
            O => \N__5000\,
            I => \N__4997\
        );

    \I__764\ : Sp12to4
    port map (
            O => \N__4997\,
            I => \N__4994\
        );

    \I__763\ : Span12Mux_s9_h
    port map (
            O => \N__4994\,
            I => \N__4991\
        );

    \I__762\ : Span12Mux_v
    port map (
            O => \N__4991\,
            I => \N__4988\
        );

    \I__761\ : Odrv12
    port map (
            O => \N__4988\,
            I => \DRDDIR_0_i\
        );

    \I__760\ : InMux
    port map (
            O => \N__4985\,
            I => \N__4982\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4982\,
            I => \U712_CHIP_RAM.N_32\
        );

    \I__758\ : IoInMux
    port map (
            O => \N__4979\,
            I => \N__4976\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__4976\,
            I => \N__4973\
        );

    \I__756\ : IoSpan4Mux
    port map (
            O => \N__4973\,
            I => \N__4970\
        );

    \I__755\ : Sp12to4
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__754\ : Odrv12
    port map (
            O => \N__4967\,
            I => \CMA_c_1\
        );

    \I__753\ : InMux
    port map (
            O => \N__4964\,
            I => \N__4961\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__4961\,
            I => \U712_CHIP_RAM.N_34\
        );

    \I__751\ : IoInMux
    port map (
            O => \N__4958\,
            I => \N__4955\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__749\ : Span4Mux_s2_h
    port map (
            O => \N__4952\,
            I => \N__4949\
        );

    \I__748\ : Span4Mux_h
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__747\ : Sp12to4
    port map (
            O => \N__4946\,
            I => \N__4943\
        );

    \I__746\ : Span12Mux_s8_v
    port map (
            O => \N__4943\,
            I => \N__4940\
        );

    \I__745\ : Span12Mux_h
    port map (
            O => \N__4940\,
            I => \N__4937\
        );

    \I__744\ : Odrv12
    port map (
            O => \N__4937\,
            I => \CMA_c_3\
        );

    \I__743\ : CascadeMux
    port map (
            O => \N__4934\,
            I => \U712_REG_SM.N_147_0_cascade_\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__4931\,
            I => \N__4928\
        );

    \I__741\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4922\
        );

    \I__740\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4922\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4922\,
            I => \U712_REG_SM.N_161_0\
        );

    \I__738\ : InMux
    port map (
            O => \N__4919\,
            I => \N__4912\
        );

    \I__737\ : InMux
    port map (
            O => \N__4918\,
            I => \N__4912\
        );

    \I__736\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4909\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__4912\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__4909\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__4904\,
            I => \U712_REG_SM.N_161_0_cascade_\
        );

    \I__732\ : InMux
    port map (
            O => \N__4901\,
            I => \N__4897\
        );

    \I__731\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4894\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4897\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__4894\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__4889\,
            I => \U712_REG_SM.N_187_cascade_\
        );

    \I__727\ : InMux
    port map (
            O => \N__4886\,
            I => \N__4883\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4883\,
            I => \U712_REG_SM.N_183\
        );

    \I__725\ : InMux
    port map (
            O => \N__4880\,
            I => \N__4871\
        );

    \I__724\ : InMux
    port map (
            O => \N__4879\,
            I => \N__4871\
        );

    \I__723\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4871\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4871\,
            I => \U712_REG_SM.N_147_0\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__4868\,
            I => \N__4865\
        );

    \I__720\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4858\
        );

    \I__719\ : InMux
    port map (
            O => \N__4864\,
            I => \N__4855\
        );

    \I__718\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4848\
        );

    \I__717\ : InMux
    port map (
            O => \N__4862\,
            I => \N__4848\
        );

    \I__716\ : InMux
    port map (
            O => \N__4861\,
            I => \N__4848\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4858\,
            I => \U712_REG_SM.N_153_0\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__4855\,
            I => \U712_REG_SM.N_153_0\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__4848\,
            I => \U712_REG_SM.N_153_0\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__4841\,
            I => \N__4838\
        );

    \I__711\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4835\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4835\,
            I => \U712_REG_SM.N_174\
        );

    \I__709\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4828\
        );

    \I__708\ : InMux
    port map (
            O => \N__4831\,
            I => \N__4825\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__4828\,
            I => \N__4822\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4825\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__705\ : Odrv4
    port map (
            O => \N__4822\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__704\ : IoInMux
    port map (
            O => \N__4817\,
            I => \N__4814\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4814\,
            I => \N__4811\
        );

    \I__702\ : Span12Mux_s0_h
    port map (
            O => \N__4811\,
            I => \N__4808\
        );

    \I__701\ : Span12Mux_h
    port map (
            O => \N__4808\,
            I => \N__4804\
        );

    \I__700\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4801\
        );

    \I__699\ : Odrv12
    port map (
            O => \N__4804\,
            I => \TACK_OUTn\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__4801\,
            I => \TACK_OUTn\
        );

    \I__697\ : IoInMux
    port map (
            O => \N__4796\,
            I => \N__4793\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__4793\,
            I => \N__4790\
        );

    \I__695\ : Span12Mux_s4_h
    port map (
            O => \N__4790\,
            I => \N__4787\
        );

    \I__694\ : Odrv12
    port map (
            O => \N__4787\,
            I => \CLK40_OUT_i_i\
        );

    \I__693\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4781\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4781\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__4778\,
            I => \U712_CHIP_RAM.N_65_cascade_\
        );

    \I__690\ : InMux
    port map (
            O => \N__4775\,
            I => \N__4771\
        );

    \I__689\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4768\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__4771\,
            I => \U712_CHIP_RAM.N_114\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__4768\,
            I => \U712_CHIP_RAM.N_114\
        );

    \I__686\ : InMux
    port map (
            O => \N__4763\,
            I => \N__4756\
        );

    \I__685\ : InMux
    port map (
            O => \N__4762\,
            I => \N__4756\
        );

    \I__684\ : InMux
    port map (
            O => \N__4761\,
            I => \N__4753\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4756\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__4753\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__681\ : CascadeMux
    port map (
            O => \N__4748\,
            I => \N__4744\
        );

    \I__680\ : InMux
    port map (
            O => \N__4747\,
            I => \N__4739\
        );

    \I__679\ : InMux
    port map (
            O => \N__4744\,
            I => \N__4732\
        );

    \I__678\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4732\
        );

    \I__677\ : InMux
    port map (
            O => \N__4742\,
            I => \N__4732\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__4739\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__4732\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__674\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4724\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4724\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_0_sqmuxa\
        );

    \I__672\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4718\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4718\,
            I => \N__4714\
        );

    \I__670\ : InMux
    port map (
            O => \N__4717\,
            I => \N__4711\
        );

    \I__669\ : Odrv4
    port map (
            O => \N__4714\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4711\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__4706\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\
        );

    \I__666\ : InMux
    port map (
            O => \N__4703\,
            I => \N__4699\
        );

    \I__665\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4696\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4699\,
            I => \U712_REG_SM.N_148_0\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4696\,
            I => \U712_REG_SM.N_148_0\
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__4691\,
            I => \U712_REG_SM.N_151_0_cascade_\
        );

    \I__661\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4685\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4685\,
            I => \U712_REG_SM.N_160_0\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__4682\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_a2_0_1_0_cascade_\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__4679\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_cascade_\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__4676\,
            I => \U712_CHIP_RAM.N_68_cascade_\
        );

    \I__656\ : InMux
    port map (
            O => \N__4673\,
            I => \N__4670\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__4670\,
            I => \U712_CHIP_RAM.N_108\
        );

    \I__654\ : InMux
    port map (
            O => \N__4667\,
            I => \N__4663\
        );

    \I__653\ : InMux
    port map (
            O => \N__4666\,
            I => \N__4660\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__4663\,
            I => \U712_CHIP_RAM.N_109\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__4660\,
            I => \U712_CHIP_RAM.N_109\
        );

    \I__650\ : CascadeMux
    port map (
            O => \N__4655\,
            I => \U712_CHIP_RAM.N_108_cascade_\
        );

    \I__649\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4649\,
            I => \N__4646\
        );

    \I__647\ : Span4Mux_v
    port map (
            O => \N__4646\,
            I => \N__4643\
        );

    \I__646\ : Sp12to4
    port map (
            O => \N__4643\,
            I => \N__4640\
        );

    \I__645\ : Span12Mux_h
    port map (
            O => \N__4640\,
            I => \N__4637\
        );

    \I__644\ : Span12Mux_v
    port map (
            O => \N__4637\,
            I => \N__4634\
        );

    \I__643\ : Odrv12
    port map (
            O => \N__4634\,
            I => \A_c_3\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__4631\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\
        );

    \I__641\ : InMux
    port map (
            O => \N__4628\,
            I => \N__4625\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__639\ : Span4Mux_v
    port map (
            O => \N__4622\,
            I => \N__4619\
        );

    \I__638\ : Sp12to4
    port map (
            O => \N__4619\,
            I => \N__4616\
        );

    \I__637\ : Span12Mux_h
    port map (
            O => \N__4616\,
            I => \N__4613\
        );

    \I__636\ : Odrv12
    port map (
            O => \N__4613\,
            I => \A_c_10\
        );

    \I__635\ : InMux
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__4607\,
            I => \N__4604\
        );

    \I__633\ : Span4Mux_v
    port map (
            O => \N__4604\,
            I => \N__4601\
        );

    \I__632\ : Span4Mux_v
    port map (
            O => \N__4601\,
            I => \N__4598\
        );

    \I__631\ : Span4Mux_v
    port map (
            O => \N__4598\,
            I => \N__4595\
        );

    \I__630\ : Sp12to4
    port map (
            O => \N__4595\,
            I => \N__4592\
        );

    \I__629\ : Odrv12
    port map (
            O => \N__4592\,
            I => \A_c_5\
        );

    \I__628\ : CascadeMux
    port map (
            O => \N__4589\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_\
        );

    \I__627\ : InMux
    port map (
            O => \N__4586\,
            I => \N__4583\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__4583\,
            I => \N__4580\
        );

    \I__625\ : Span12Mux_h
    port map (
            O => \N__4580\,
            I => \N__4577\
        );

    \I__624\ : Odrv12
    port map (
            O => \N__4577\,
            I => \A_c_12\
        );

    \I__623\ : InMux
    port map (
            O => \N__4574\,
            I => \N__4571\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__4571\,
            I => \N__4568\
        );

    \I__621\ : Span4Mux_v
    port map (
            O => \N__4568\,
            I => \N__4565\
        );

    \I__620\ : Sp12to4
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__619\ : Span12Mux_h
    port map (
            O => \N__4562\,
            I => \N__4559\
        );

    \I__618\ : Span12Mux_v
    port map (
            O => \N__4559\,
            I => \N__4556\
        );

    \I__617\ : Odrv12
    port map (
            O => \N__4556\,
            I => \DBRn_c\
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__4553\,
            I => \U712_CHIP_RAM.N_61_cascade_\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__4550\,
            I => \U712_CHIP_RAM.N_101_cascade_\
        );

    \I__614\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4541\
        );

    \I__613\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4541\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4541\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__611\ : InMux
    port map (
            O => \N__4538\,
            I => \N__4533\
        );

    \I__610\ : InMux
    port map (
            O => \N__4537\,
            I => \N__4528\
        );

    \I__609\ : InMux
    port map (
            O => \N__4536\,
            I => \N__4528\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__4533\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__4528\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__606\ : InMux
    port map (
            O => \N__4523\,
            I => \N__4520\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4520\,
            I => \U712_REG_SM.N_181\
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__4517\,
            I => \U712_REG_SM.DS_EN_7_0_cascade_\
        );

    \I__603\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4511\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4511\,
            I => \N__4507\
        );

    \I__601\ : IoInMux
    port map (
            O => \N__4510\,
            I => \N__4504\
        );

    \I__600\ : Span4Mux_v
    port map (
            O => \N__4507\,
            I => \N__4501\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4504\,
            I => \N__4498\
        );

    \I__598\ : Sp12to4
    port map (
            O => \N__4501\,
            I => \N__4495\
        );

    \I__597\ : Span4Mux_s3_h
    port map (
            O => \N__4498\,
            I => \N__4492\
        );

    \I__596\ : Span12Mux_h
    port map (
            O => \N__4495\,
            I => \N__4487\
        );

    \I__595\ : Sp12to4
    port map (
            O => \N__4492\,
            I => \N__4487\
        );

    \I__594\ : Span12Mux_v
    port map (
            O => \N__4487\,
            I => \N__4484\
        );

    \I__593\ : Odrv12
    port map (
            O => \N__4484\,
            I => \C1_c\
        );

    \I__592\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4478\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4478\,
            I => \N__4475\
        );

    \I__590\ : Span12Mux_h
    port map (
            O => \N__4475\,
            I => \N__4472\
        );

    \I__589\ : Span12Mux_v
    port map (
            O => \N__4472\,
            I => \N__4469\
        );

    \I__588\ : Odrv12
    port map (
            O => \N__4469\,
            I => \C3_c\
        );

    \I__587\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4463\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4463\,
            I => \N__4460\
        );

    \I__585\ : Span4Mux_v
    port map (
            O => \N__4460\,
            I => \N__4456\
        );

    \I__584\ : InMux
    port map (
            O => \N__4459\,
            I => \N__4453\
        );

    \I__583\ : Odrv4
    port map (
            O => \N__4456\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__4453\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__581\ : IoInMux
    port map (
            O => \N__4448\,
            I => \N__4445\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4445\,
            I => \N__4442\
        );

    \I__579\ : Span4Mux_s3_v
    port map (
            O => \N__4442\,
            I => \N__4439\
        );

    \I__578\ : Span4Mux_h
    port map (
            O => \N__4439\,
            I => \N__4436\
        );

    \I__577\ : Sp12to4
    port map (
            O => \N__4436\,
            I => \N__4433\
        );

    \I__576\ : Span12Mux_v
    port map (
            O => \N__4433\,
            I => \N__4430\
        );

    \I__575\ : Span12Mux_h
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__574\ : Odrv12
    port map (
            O => \N__4427\,
            I => \U712_REG_SM_un1_LDSn_i\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__572\ : InMux
    port map (
            O => \N__4421\,
            I => \N__4418\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__570\ : Odrv4
    port map (
            O => \N__4415\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__569\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4409\,
            I => \U712_REG_SM.N_175\
        );

    \I__567\ : InMux
    port map (
            O => \N__4406\,
            I => \N__4401\
        );

    \I__566\ : InMux
    port map (
            O => \N__4405\,
            I => \N__4396\
        );

    \I__565\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4396\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4401\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4396\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__562\ : InMux
    port map (
            O => \N__4391\,
            I => \N__4387\
        );

    \I__561\ : InMux
    port map (
            O => \N__4390\,
            I => \N__4384\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4387\,
            I => \U712_REG_SM.N_156_0\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4384\,
            I => \U712_REG_SM.N_156_0\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__4379\,
            I => \U712_REG_SM.N_156_0_cascade_\
        );

    \I__557\ : InMux
    port map (
            O => \N__4376\,
            I => \N__4373\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4373\,
            I => \U712_REG_SM.N_166_0\
        );

    \I__555\ : InMux
    port map (
            O => \N__4370\,
            I => \N__4363\
        );

    \I__554\ : InMux
    port map (
            O => \N__4369\,
            I => \N__4363\
        );

    \I__553\ : InMux
    port map (
            O => \N__4368\,
            I => \N__4360\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__4363\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__4360\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__4355\,
            I => \U712_REG_SM.N_148_0_cascade_\
        );

    \I__549\ : InMux
    port map (
            O => \N__4352\,
            I => \N__4347\
        );

    \I__548\ : InMux
    port map (
            O => \N__4351\,
            I => \N__4342\
        );

    \I__547\ : InMux
    port map (
            O => \N__4350\,
            I => \N__4342\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__4347\,
            I => \U712_REG_SM.N_164_0\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__4342\,
            I => \U712_REG_SM.N_164_0\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__4337\,
            I => \N__4333\
        );

    \I__543\ : InMux
    port map (
            O => \N__4336\,
            I => \N__4330\
        );

    \I__542\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4327\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__4330\,
            I => \N__4322\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4327\,
            I => \N__4322\
        );

    \I__539\ : Span4Mux_v
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__538\ : Sp12to4
    port map (
            O => \N__4319\,
            I => \N__4316\
        );

    \I__537\ : Span12Mux_h
    port map (
            O => \N__4316\,
            I => \N__4313\
        );

    \I__536\ : Odrv12
    port map (
            O => \N__4313\,
            I => \REGSPACEn_c\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__4310\,
            I => \N__4306\
        );

    \I__534\ : InMux
    port map (
            O => \N__4309\,
            I => \N__4303\
        );

    \I__533\ : InMux
    port map (
            O => \N__4306\,
            I => \N__4300\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__4303\,
            I => \N__4296\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__4300\,
            I => \N__4293\
        );

    \I__530\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4290\
        );

    \I__529\ : Span4Mux_v
    port map (
            O => \N__4296\,
            I => \N__4285\
        );

    \I__528\ : Span4Mux_v
    port map (
            O => \N__4293\,
            I => \N__4285\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4290\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__526\ : Odrv4
    port map (
            O => \N__4285\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__525\ : CascadeMux
    port map (
            O => \N__4280\,
            I => \N__4276\
        );

    \I__524\ : InMux
    port map (
            O => \N__4279\,
            I => \N__4271\
        );

    \I__523\ : InMux
    port map (
            O => \N__4276\,
            I => \N__4271\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4271\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0\
        );

    \I__521\ : CascadeMux
    port map (
            O => \N__4268\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_cascade_\
        );

    \I__520\ : CascadeMux
    port map (
            O => \N__4265\,
            I => \U712_REG_SM.N_175_cascade_\
        );

    \I__519\ : CEMux
    port map (
            O => \N__4262\,
            I => \N__4259\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4259\,
            I => \N__4256\
        );

    \I__517\ : Odrv4
    port map (
            O => \N__4256\,
            I => \U712_REG_SM.N_175_0_0\
        );

    \I__516\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4250\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa_1\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__4247\,
            I => \U712_REG_SM.N_178_cascade_\
        );

    \I__513\ : InMux
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__4241\,
            I => \U712_REG_SM.N_163_0\
        );

    \I__511\ : InMux
    port map (
            O => \N__4238\,
            I => \N__4234\
        );

    \I__510\ : InMux
    port map (
            O => \N__4237\,
            I => \N__4231\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4234\,
            I => \N__4228\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4231\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__507\ : Odrv4
    port map (
            O => \N__4228\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__506\ : InMux
    port map (
            O => \N__4223\,
            I => \N__4220\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4220\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__504\ : InMux
    port map (
            O => \N__4217\,
            I => \N__4214\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4214\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__502\ : CascadeMux
    port map (
            O => \N__4211\,
            I => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__4208\,
            I => \U712_CYCLE_TERM.N_45_0_0_en_cascade_\
        );

    \I__500\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4202\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4202\,
            I => \TACK_EN_i_ess\
        );

    \I__498\ : CEMux
    port map (
            O => \N__4199\,
            I => \N__4196\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4196\,
            I => \N__4193\
        );

    \I__496\ : Span4Mux_v
    port map (
            O => \N__4193\,
            I => \N__4190\
        );

    \I__495\ : Span4Mux_h
    port map (
            O => \N__4190\,
            I => \N__4187\
        );

    \I__494\ : Odrv4
    port map (
            O => \N__4187\,
            I => \U712_CYCLE_TERM.N_45_0_0_en_0\
        );

    \I__493\ : InMux
    port map (
            O => \N__4184\,
            I => \N__4180\
        );

    \I__492\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4177\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4180\,
            I => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4177\,
            I => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1\
        );

    \I__489\ : InMux
    port map (
            O => \N__4172\,
            I => \N__4169\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4169\,
            I => \U712_BYTE_ENABLE.LMBE_0\
        );

    \I__487\ : IoInMux
    port map (
            O => \N__4166\,
            I => \N__4163\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__485\ : IoSpan4Mux
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__484\ : Sp12to4
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__483\ : Span12Mux_s9_h
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__482\ : Span12Mux_h
    port map (
            O => \N__4151\,
            I => \N__4148\
        );

    \I__481\ : Span12Mux_v
    port map (
            O => \N__4148\,
            I => \N__4145\
        );

    \I__480\ : Odrv12
    port map (
            O => \N__4145\,
            I => \CLMBEn_c\
        );

    \I__479\ : IoInMux
    port map (
            O => \N__4142\,
            I => \N__4139\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4139\,
            I => \N__4136\
        );

    \I__477\ : Span12Mux_s4_v
    port map (
            O => \N__4136\,
            I => \N__4133\
        );

    \I__476\ : Odrv12
    port map (
            O => \N__4133\,
            I => \VBENn_c\
        );

    \I__475\ : InMux
    port map (
            O => \N__4130\,
            I => \N__4122\
        );

    \I__474\ : InMux
    port map (
            O => \N__4129\,
            I => \N__4122\
        );

    \I__473\ : CascadeMux
    port map (
            O => \N__4128\,
            I => \N__4119\
        );

    \I__472\ : IoInMux
    port map (
            O => \N__4127\,
            I => \N__4116\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4122\,
            I => \N__4113\
        );

    \I__470\ : InMux
    port map (
            O => \N__4119\,
            I => \N__4110\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4116\,
            I => \N__4107\
        );

    \I__468\ : Span4Mux_v
    port map (
            O => \N__4113\,
            I => \N__4102\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4110\,
            I => \N__4102\
        );

    \I__466\ : Span12Mux_s11_v
    port map (
            O => \N__4107\,
            I => \N__4098\
        );

    \I__465\ : Span4Mux_v
    port map (
            O => \N__4102\,
            I => \N__4095\
        );

    \I__464\ : InMux
    port map (
            O => \N__4101\,
            I => \N__4092\
        );

    \I__463\ : Odrv12
    port map (
            O => \N__4098\,
            I => \DBENn_c\
        );

    \I__462\ : Odrv4
    port map (
            O => \N__4095\,
            I => \DBENn_c\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4092\,
            I => \DBENn_c\
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__4085\,
            I => \U712_BYTE_ENABLE.LLBE_0_cascade_\
        );

    \I__459\ : IoInMux
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__457\ : IoSpan4Mux
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__456\ : Span4Mux_s3_v
    port map (
            O => \N__4073\,
            I => \N__4070\
        );

    \I__455\ : Sp12to4
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__454\ : Span12Mux_s8_v
    port map (
            O => \N__4067\,
            I => \N__4064\
        );

    \I__453\ : Odrv12
    port map (
            O => \N__4064\,
            I => \CLLBEn_c\
        );

    \I__452\ : InMux
    port map (
            O => \N__4061\,
            I => \N__4054\
        );

    \I__451\ : InMux
    port map (
            O => \N__4060\,
            I => \N__4047\
        );

    \I__450\ : InMux
    port map (
            O => \N__4059\,
            I => \N__4047\
        );

    \I__449\ : InMux
    port map (
            O => \N__4058\,
            I => \N__4047\
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__4057\,
            I => \N__4043\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__4054\,
            I => \N__4038\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__4047\,
            I => \N__4038\
        );

    \I__445\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4033\
        );

    \I__444\ : InMux
    port map (
            O => \N__4043\,
            I => \N__4033\
        );

    \I__443\ : Span4Mux_v
    port map (
            O => \N__4038\,
            I => \N__4028\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4033\,
            I => \N__4028\
        );

    \I__441\ : Span4Mux_h
    port map (
            O => \N__4028\,
            I => \N__4025\
        );

    \I__440\ : Span4Mux_v
    port map (
            O => \N__4025\,
            I => \N__4022\
        );

    \I__439\ : Sp12to4
    port map (
            O => \N__4022\,
            I => \N__4019\
        );

    \I__438\ : Odrv12
    port map (
            O => \N__4019\,
            I => \A_c_0\
        );

    \I__437\ : InMux
    port map (
            O => \N__4016\,
            I => \N__4009\
        );

    \I__436\ : InMux
    port map (
            O => \N__4015\,
            I => \N__4009\
        );

    \I__435\ : CascadeMux
    port map (
            O => \N__4014\,
            I => \N__4006\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__4009\,
            I => \N__4002\
        );

    \I__433\ : InMux
    port map (
            O => \N__4006\,
            I => \N__3997\
        );

    \I__432\ : InMux
    port map (
            O => \N__4005\,
            I => \N__3997\
        );

    \I__431\ : Span4Mux_h
    port map (
            O => \N__4002\,
            I => \N__3992\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3997\,
            I => \N__3992\
        );

    \I__429\ : Span4Mux_v
    port map (
            O => \N__3992\,
            I => \N__3989\
        );

    \I__428\ : Span4Mux_v
    port map (
            O => \N__3989\,
            I => \N__3986\
        );

    \I__427\ : Sp12to4
    port map (
            O => \N__3986\,
            I => \N__3983\
        );

    \I__426\ : Odrv12
    port map (
            O => \N__3983\,
            I => \A_c_1\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__3980\,
            I => \U712_BYTE_ENABLE.N_79_cascade_\
        );

    \I__424\ : CascadeMux
    port map (
            O => \N__3977\,
            I => \N__3973\
        );

    \I__423\ : CascadeMux
    port map (
            O => \N__3976\,
            I => \N__3968\
        );

    \I__422\ : InMux
    port map (
            O => \N__3973\,
            I => \N__3963\
        );

    \I__421\ : InMux
    port map (
            O => \N__3972\,
            I => \N__3963\
        );

    \I__420\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3958\
        );

    \I__419\ : InMux
    port map (
            O => \N__3968\,
            I => \N__3958\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3963\,
            I => \N__3953\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3958\,
            I => \N__3953\
        );

    \I__416\ : Span4Mux_v
    port map (
            O => \N__3953\,
            I => \N__3947\
        );

    \I__415\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3944\
        );

    \I__414\ : InMux
    port map (
            O => \N__3951\,
            I => \N__3939\
        );

    \I__413\ : InMux
    port map (
            O => \N__3950\,
            I => \N__3939\
        );

    \I__412\ : Sp12to4
    port map (
            O => \N__3947\,
            I => \N__3932\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__3944\,
            I => \N__3932\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3939\,
            I => \N__3932\
        );

    \I__409\ : Span12Mux_s11_h
    port map (
            O => \N__3932\,
            I => \N__3929\
        );

    \I__408\ : Span12Mux_v
    port map (
            O => \N__3929\,
            I => \N__3926\
        );

    \I__407\ : Odrv12
    port map (
            O => \N__3926\,
            I => \SIZ_c_0\
        );

    \I__406\ : InMux
    port map (
            O => \N__3923\,
            I => \N__3915\
        );

    \I__405\ : InMux
    port map (
            O => \N__3922\,
            I => \N__3915\
        );

    \I__404\ : InMux
    port map (
            O => \N__3921\,
            I => \N__3910\
        );

    \I__403\ : InMux
    port map (
            O => \N__3920\,
            I => \N__3910\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3915\,
            I => \N__3907\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__3910\,
            I => \N__3904\
        );

    \I__400\ : Sp12to4
    port map (
            O => \N__3907\,
            I => \N__3901\
        );

    \I__399\ : Span12Mux_h
    port map (
            O => \N__3904\,
            I => \N__3898\
        );

    \I__398\ : Span12Mux_v
    port map (
            O => \N__3901\,
            I => \N__3895\
        );

    \I__397\ : Span12Mux_v
    port map (
            O => \N__3898\,
            I => \N__3892\
        );

    \I__396\ : Odrv12
    port map (
            O => \N__3895\,
            I => \SIZ_c_1\
        );

    \I__395\ : Odrv12
    port map (
            O => \N__3892\,
            I => \SIZ_c_1\
        );

    \I__394\ : CascadeMux
    port map (
            O => \N__3887\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_iZ0Z_0_cascade_\
        );

    \I__393\ : IoInMux
    port map (
            O => \N__3884\,
            I => \N__3881\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__3881\,
            I => \N__3878\
        );

    \I__391\ : IoSpan4Mux
    port map (
            O => \N__3878\,
            I => \N__3875\
        );

    \I__390\ : Span4Mux_s3_h
    port map (
            O => \N__3875\,
            I => \N__3872\
        );

    \I__389\ : Span4Mux_v
    port map (
            O => \N__3872\,
            I => \N__3869\
        );

    \I__388\ : Span4Mux_v
    port map (
            O => \N__3869\,
            I => \N__3866\
        );

    \I__387\ : Sp12to4
    port map (
            O => \N__3866\,
            I => \N__3863\
        );

    \I__386\ : Span12Mux_s10_h
    port map (
            O => \N__3863\,
            I => \N__3860\
        );

    \I__385\ : Span12Mux_h
    port map (
            O => \N__3860\,
            I => \N__3857\
        );

    \I__384\ : Odrv12
    port map (
            O => \N__3857\,
            I => \N_54_i\
        );

    \I__383\ : SRMux
    port map (
            O => \N__3854\,
            I => \N__3851\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3851\,
            I => \N__3848\
        );

    \I__381\ : Span4Mux_h
    port map (
            O => \N__3848\,
            I => \N__3845\
        );

    \I__380\ : Odrv4
    port map (
            O => \N__3845\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__379\ : CascadeMux
    port map (
            O => \N__3842\,
            I => \U712_REG_SM.N_163_0_cascade_\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__3839\,
            I => \N_71_cascade_\
        );

    \I__377\ : IoInMux
    port map (
            O => \N__3836\,
            I => \N__3833\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__3833\,
            I => \N__3830\
        );

    \I__375\ : Span4Mux_s1_h
    port map (
            O => \N__3830\,
            I => \N__3827\
        );

    \I__374\ : Span4Mux_h
    port map (
            O => \N__3827\,
            I => \N__3824\
        );

    \I__373\ : Sp12to4
    port map (
            O => \N__3824\,
            I => \N__3821\
        );

    \I__372\ : Span12Mux_v
    port map (
            O => \N__3821\,
            I => \N__3818\
        );

    \I__371\ : Odrv12
    port map (
            O => \N__3818\,
            I => \N_736_i\
        );

    \I__370\ : InMux
    port map (
            O => \N__3815\,
            I => \N__3812\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__3812\,
            I => \U712_REG_SM.UDS_OUT_2_0_a2_0\
        );

    \I__368\ : InMux
    port map (
            O => \N__3809\,
            I => \N__3806\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__3806\,
            I => \U712_BYTE_ENABLE.N_82\
        );

    \I__366\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3800\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__3800\,
            I => \U712_BYTE_ENABLE.un1_CUUBEn_iZ0Z_0\
        );

    \I__364\ : IoInMux
    port map (
            O => \N__3797\,
            I => \N__3794\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3794\,
            I => \N__3791\
        );

    \I__362\ : Span4Mux_s1_h
    port map (
            O => \N__3791\,
            I => \N__3788\
        );

    \I__361\ : Sp12to4
    port map (
            O => \N__3788\,
            I => \N__3785\
        );

    \I__360\ : Span12Mux_v
    port map (
            O => \N__3785\,
            I => \N__3782\
        );

    \I__359\ : Span12Mux_h
    port map (
            O => \N__3782\,
            I => \N__3779\
        );

    \I__358\ : Odrv12
    port map (
            O => \N__3779\,
            I => \N_55_i\
        );

    \I__357\ : InMux
    port map (
            O => \N__3776\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__356\ : InMux
    port map (
            O => \N__3773\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__355\ : InMux
    port map (
            O => \N__3770\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__354\ : InMux
    port map (
            O => \N__3767\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__353\ : InMux
    port map (
            O => \N__3764\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__352\ : ClkMux
    port map (
            O => \N__3761\,
            I => \N__3758\
        );

    \I__351\ : GlobalMux
    port map (
            O => \N__3758\,
            I => \N__3755\
        );

    \I__350\ : gio2CtrlBuf
    port map (
            O => \N__3755\,
            I => \C1_c_g\
        );

    \I__349\ : InMux
    port map (
            O => \N__3752\,
            I => \N__3748\
        );

    \I__348\ : InMux
    port map (
            O => \N__3751\,
            I => \N__3745\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__3748\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__3745\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__345\ : InMux
    port map (
            O => \N__3740\,
            I => \N__3736\
        );

    \I__344\ : InMux
    port map (
            O => \N__3739\,
            I => \N__3733\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3736\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3733\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__341\ : InMux
    port map (
            O => \N__3728\,
            I => \N__3724\
        );

    \I__340\ : InMux
    port map (
            O => \N__3727\,
            I => \N__3721\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__3724\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__3721\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__337\ : InMux
    port map (
            O => \N__3716\,
            I => \N__3712\
        );

    \I__336\ : InMux
    port map (
            O => \N__3715\,
            I => \N__3709\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__3712\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__3709\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__333\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3700\
        );

    \I__332\ : InMux
    port map (
            O => \N__3703\,
            I => \N__3697\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__3700\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__3697\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__329\ : CascadeMux
    port map (
            O => \N__3692\,
            I => \N__3688\
        );

    \I__328\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3685\
        );

    \I__327\ : InMux
    port map (
            O => \N__3688\,
            I => \N__3682\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__3685\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__3682\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__324\ : InMux
    port map (
            O => \N__3677\,
            I => \N__3673\
        );

    \I__323\ : InMux
    port map (
            O => \N__3676\,
            I => \N__3670\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__3673\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__3670\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__320\ : IoInMux
    port map (
            O => \N__3665\,
            I => \N__3662\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__3662\,
            I => \N__3659\
        );

    \I__318\ : Span12Mux_s6_v
    port map (
            O => \N__3659\,
            I => \N__3656\
        );

    \I__317\ : Odrv12
    port map (
            O => \N__3656\,
            I => \CLK80_OUT_i_i\
        );

    \I__316\ : InMux
    port map (
            O => \N__3653\,
            I => \bfn_6_8_0_\
        );

    \I__315\ : InMux
    port map (
            O => \N__3650\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__314\ : InMux
    port map (
            O => \N__3647\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__313\ : IoInMux
    port map (
            O => \N__3644\,
            I => \N__3641\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__3641\,
            I => \N__3638\
        );

    \I__311\ : Span4Mux_s0_v
    port map (
            O => \N__3638\,
            I => \N__3635\
        );

    \I__310\ : Span4Mux_v
    port map (
            O => \N__3635\,
            I => \N__3632\
        );

    \I__309\ : Sp12to4
    port map (
            O => \N__3632\,
            I => \N__3629\
        );

    \I__308\ : Span12Mux_h
    port map (
            O => \N__3629\,
            I => \N__3626\
        );

    \I__307\ : Span12Mux_v
    port map (
            O => \N__3626\,
            I => \N__3623\
        );

    \I__306\ : Odrv12
    port map (
            O => \N__3623\,
            I => \CLK40_IN_c\
        );

    \IN_MUX_bfv_6_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_8_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7136\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4510\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8432\,
            lcout => \CLK80_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3704\,
            in2 => \_gnd_net_\,
            in3 => \N__3653\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_6_8_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__3761\,
            ce => 'H',
            sr => \N__3854\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3677\,
            in2 => \_gnd_net_\,
            in3 => \N__3650\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__3761\,
            ce => 'H',
            sr => \N__3854\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3716\,
            in2 => \_gnd_net_\,
            in3 => \N__3647\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__3761\,
            ce => 'H',
            sr => \N__3854\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4237\,
            in2 => \_gnd_net_\,
            in3 => \N__3776\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__3761\,
            ce => 'H',
            sr => \N__3854\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3691\,
            in2 => \_gnd_net_\,
            in3 => \N__3773\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__3761\,
            ce => 'H',
            sr => \N__3854\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3728\,
            in2 => \_gnd_net_\,
            in3 => \N__3770\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__3761\,
            ce => 'H',
            sr => \N__3854\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3740\,
            in2 => \_gnd_net_\,
            in3 => \N__3767\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__3761\,
            ce => 'H',
            sr => \N__3854\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3752\,
            in2 => \_gnd_net_\,
            in3 => \N__3764\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3761\,
            ce => 'H',
            sr => \N__3854\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__3751\,
            in1 => \N__3739\,
            in2 => \_gnd_net_\,
            in3 => \N__3727\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__3715\,
            in1 => \N__3703\,
            in2 => \N__3692\,
            in3 => \N__3676\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__8143\,
            in1 => \N__3809\,
            in2 => \N__4128\,
            in3 => \N__6884\,
            lcout => \U712_BYTE_ENABLE.un1_CUUBEn_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_o2_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__4061\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3972\,
            lcout => OPEN,
            ltout => \N_71_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDS_OUT_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__5760\,
            in1 => \N__4459\,
            in2 => \N__3839\,
            in3 => \N__4351\,
            lcout => \U712_REG_SM.LDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8427\,
            ce => 'H',
            sr => \N__9385\
        );

    \U712_REG_SM.UDS_OUT_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111111001100"
        )
    port map (
            in0 => \N__3815\,
            in1 => \N__5074\,
            in2 => \N__3977\,
            in3 => \N__4350\,
            lcout => \U712_REG_SM.UDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8427\,
            ce => 'H',
            sr => \N__9385\
        );

    \TACKn_obuft_RNO_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4205\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_736_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_RNO_0_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4060\,
            in2 => \_gnd_net_\,
            in3 => \N__5759\,
            lcout => \U712_REG_SM.UDS_OUT_2_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4059\,
            in1 => \N__4016\,
            in2 => \_gnd_net_\,
            in3 => \N__8625\,
            lcout => \U712_BYTE_ENABLE.N_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LMBE_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110110000"
        )
    port map (
            in0 => \N__4058\,
            in1 => \N__4015\,
            in2 => \N__3976\,
            in3 => \N__3922\,
            lcout => \U712_BYTE_ENABLE.LMBE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_55_i_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100100011"
        )
    port map (
            in0 => \N__3923\,
            in1 => \N__3803\,
            in2 => \N__8635\,
            in3 => \N__3971\,
            lcout => \N_55_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un3_CLLBEn_1_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6895\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4130\,
            lcout => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101000100"
        )
    port map (
            in0 => \N__4005\,
            in1 => \N__3920\,
            in2 => \N__4057\,
            in3 => \N__3950\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.LLBE_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100110001"
        )
    port map (
            in0 => \N__8617\,
            in1 => \N__4183\,
            in2 => \N__4085\,
            in3 => \N__8178\,
            lcout => \CLLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100000000"
        )
    port map (
            in0 => \N__4046\,
            in1 => \N__3951\,
            in2 => \N__4014\,
            in3 => \N__8618\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_79_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__4129\,
            in1 => \N__8179\,
            in2 => \N__3980\,
            in3 => \N__6894\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.un1_CUMBEn_iZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_54_i_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000001111"
        )
    port map (
            in0 => \N__3952\,
            in1 => \N__3921\,
            in2 => \N__3887\,
            in3 => \N__8616\,
            lcout => \N_54_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9134\,
            in1 => \N__8971\,
            in2 => \N__8823\,
            in3 => \N__9249\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_esr_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4406\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8419\,
            ce => \N__4262\,
            sr => \N__9393\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4390\,
            in2 => \_gnd_net_\,
            in3 => \N__4703\,
            lcout => \U712_REG_SM.N_163_0\,
            ltout => \U712_REG_SM.N_163_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3842\,
            in3 => \N__4369\,
            lcout => \U712_REG_SM.N_164_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000101"
        )
    port map (
            in0 => \N__4370\,
            in1 => \N__5394\,
            in2 => \N__4310\,
            in3 => \N__4336\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_178_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001100"
        )
    port map (
            in0 => \N__4309\,
            in1 => \N__7319\,
            in2 => \N__4247\,
            in3 => \N__4244\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8422\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010110000"
        )
    port map (
            in0 => \N__4238\,
            in1 => \N__4223\,
            in2 => \N__7331\,
            in3 => \N__4217\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7048\,
            in2 => \_gnd_net_\,
            in3 => \N__7030\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010101010"
        )
    port map (
            in0 => \N__6004\,
            in1 => \N__6950\,
            in2 => \N__4211\,
            in3 => \N__7318\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_45_0_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9457\,
            in1 => \_gnd_net_\,
            in2 => \N__4208\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.N_45_0_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__7279\,
            in1 => \N__4831\,
            in2 => \_gnd_net_\,
            in3 => \N__6956\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8428\,
            ce => \N__4199\,
            sr => \N__9365\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000101"
        )
    port map (
            in0 => \N__4184\,
            in1 => \N__4172\,
            in2 => \N__8636\,
            in3 => \N__8136\,
            lcout => \CLMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6829\,
            in2 => \_gnd_net_\,
            in3 => \N__8586\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111111101110000"
        )
    port map (
            in0 => \N__5600\,
            in1 => \N__7640\,
            in2 => \N__4280\,
            in3 => \N__4101\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8407\,
            ce => 'H',
            sr => \N__9402\
        );

    \U712_CHIP_RAM.DMA_CYCLE_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6856\,
            in1 => \N__5599\,
            in2 => \_gnd_net_\,
            in3 => \N__4279\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8407\,
            ce => 'H',
            sr => \N__9402\
        );

    \U712_CHIP_RAM.DBDIR_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__4721\,
            in1 => \N__5833\,
            in2 => \_gnd_net_\,
            in3 => \N__5025\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8407\,
            ce => 'H',
            sr => \N__9402\
        );

    \U712_REG_SM.C1_SYNC_2_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5297\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8413\,
            ce => 'H',
            sr => \N__9394\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__5407\,
            in1 => \N__4299\,
            in2 => \N__4337\,
            in3 => \N__4253\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8413\,
            ce => 'H',
            sr => \N__9394\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_2_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__6202\,
            in1 => \N__4775\,
            in2 => \_gnd_net_\,
            in3 => \N__4717\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__8522\,
            in1 => \N__6530\,
            in2 => \N__4268\,
            in3 => \N__5796\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8413\,
            ce => 'H',
            sr => \N__9394\
        );

    \U712_REG_SM.STATE_COUNT_RNIFFKI2_4_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__7074\,
            in1 => \N__4404\,
            in2 => \_gnd_net_\,
            in3 => \N__5580\,
            lcout => \U712_REG_SM.N_175\,
            ltout => \U712_REG_SM.N_175_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_esr_RNO_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__9459\,
            in1 => \_gnd_net_\,
            in2 => \N__4265\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.N_175_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI20MC2_2_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__5188\,
            in1 => \N__5267\,
            in2 => \_gnd_net_\,
            in3 => \N__5158\,
            lcout => \U712_REG_SM.DS_EN_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__7295\,
            in1 => \N__6871\,
            in2 => \N__4424\,
            in3 => \N__8523\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8417\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__4412\,
            in1 => \N__7297\,
            in2 => \N__4868\,
            in3 => \N__4391\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8417\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010001000"
        )
    port map (
            in0 => \N__7296\,
            in1 => \N__4688\,
            in2 => \N__5585\,
            in3 => \N__4405\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8417\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__7299\,
            in1 => \N__4376\,
            in2 => \N__4841\,
            in3 => \N__4901\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8420\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_1_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5202\,
            in1 => \N__5322\,
            in2 => \N__5293\,
            in3 => \N__5266\,
            lcout => \U712_REG_SM.N_156_0\,
            ltout => \U712_REG_SM.N_156_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7075\,
            in2 => \N__4379\,
            in3 => \N__4864\,
            lcout => \U712_REG_SM.N_166_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4546\,
            in2 => \_gnd_net_\,
            in3 => \N__4536\,
            lcout => \U712_REG_SM.N_148_0\,
            ltout => \U712_REG_SM.N_148_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNINB3L1_1_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5321\,
            in1 => \N__4368\,
            in2 => \N__4355\,
            in3 => \N__5286\,
            lcout => \U712_REG_SM.N_183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__4919\,
            in1 => \N__7298\,
            in2 => \N__4931\,
            in3 => \N__4352\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8420\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4918\,
            in2 => \_gnd_net_\,
            in3 => \N__4927\,
            lcout => \U712_REG_SM.N_181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI90BP_0_2_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4547\,
            in2 => \_gnd_net_\,
            in3 => \N__4537\,
            lcout => \U712_REG_SM.N_153_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_2_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4538\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8423\,
            ce => 'H',
            sr => \N__9366\
        );

    \U712_REG_SM.C3_SYNC_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5260\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8423\,
            ce => 'H',
            sr => \N__9366\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__5259\,
            in1 => \N__5762\,
            in2 => \_gnd_net_\,
            in3 => \N__5323\,
            lcout => OPEN,
            ltout => \U712_REG_SM.DS_EN_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111101001110"
        )
    port map (
            in0 => \N__4523\,
            in1 => \N__5097\,
            in2 => \N__4517\,
            in3 => \N__5987\,
            lcout => \U712_REG_SM.DS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8423\,
            ce => 'H',
            sr => \N__9366\
        );

    \U712_REG_SM.C1_SYNC_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4514\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8423\,
            ce => 'H',
            sr => \N__9366\
        );

    \U712_REG_SM.C3_SYNC_0_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4481\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8426\,
            ce => 'H',
            sr => \N__9360\
        );

    \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__4466\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5104\,
            lcout => \U712_REG_SM_un1_LDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__7118\,
            in1 => \N__8596\,
            in2 => \N__7880\,
            in3 => \N__9098\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__8598\,
            in1 => \N__4652\,
            in2 => \N__4631\,
            in3 => \N__4628\,
            lcout => \U712_CHIP_RAM.N_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__7739\,
            in1 => \N__8595\,
            in2 => \N__9132\,
            in3 => \N__7796\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__8597\,
            in1 => \N__4610\,
            in2 => \N__4589\,
            in3 => \N__4586\,
            lcout => \U712_CHIP_RAM.N_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBR_SYNC_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4574\,
            lcout => \U712_REG_SM_DBR_SYNC_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8402\,
            ce => 'H',
            sr => \N__9395\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5523\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM_DBR_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8402\,
            ce => 'H',
            sr => \N__9395\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__5522\,
            in1 => \N__5788\,
            in2 => \N__5559\,
            in3 => \N__6291\,
            lcout => \U712_CHIP_RAM.N_61\,
            ltout => \U712_CHIP_RAM.N_61_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRB433_2_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001001"
        )
    port map (
            in0 => \N__6139\,
            in1 => \N__6595\,
            in2 => \N__4553\,
            in3 => \N__6511\,
            lcout => \U712_CHIP_RAM.N_421_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKLSF6_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__7328\,
            in1 => \N__4667\,
            in2 => \N__6206\,
            in3 => \N__4673\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_101_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHPUTC_3_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__5330\,
            in1 => \N__6437\,
            in2 => \N__4550\,
            in3 => \N__7329\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOO5O1_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6576\,
            in1 => \N__6136\,
            in2 => \N__7441\,
            in3 => \N__6088\,
            lcout => \U712_CHIP_RAM.N_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6138\,
            in1 => \N__6263\,
            in2 => \N__7443\,
            in3 => \N__6578\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_a2_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000000"
        )
    port map (
            in0 => \N__6438\,
            in1 => \N__7314\,
            in2 => \N__4682\,
            in3 => \N__6716\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__5428\,
            in1 => \_gnd_net_\,
            in2 => \N__4679\,
            in3 => \N__8970\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__6857\,
            in1 => \N__5795\,
            in2 => \N__7763\,
            in3 => \N__7313\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__6089\,
            in1 => \N__4747\,
            in2 => \_gnd_net_\,
            in3 => \N__4761\,
            lcout => \U712_CHIP_RAM.N_68\,
            ltout => \U712_CHIP_RAM.N_68_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_0_2_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__6577\,
            in1 => \N__7425\,
            in2 => \N__4676\,
            in3 => \N__6137\,
            lcout => \U712_CHIP_RAM.N_108\,
            ltout => \U712_CHIP_RAM.N_108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMMGI5_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4666\,
            in2 => \N__4655\,
            in3 => \N__4774\,
            lcout => \U712_CHIP_RAM.N_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__4784\,
            in1 => \N__7293\,
            in2 => \N__4748\,
            in3 => \N__4727\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__6526\,
            in1 => \N__6581\,
            in2 => \_gnd_net_\,
            in3 => \N__5645\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100001"
        )
    port map (
            in0 => \N__6580\,
            in1 => \N__5485\,
            in2 => \N__6529\,
            in3 => \N__6241\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__6087\,
            in1 => \N__4762\,
            in2 => \_gnd_net_\,
            in3 => \N__4742\,
            lcout => \U712_CHIP_RAM.N_65\,
            ltout => \U712_CHIP_RAM.N_65_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__6579\,
            in1 => \N__7418\,
            in2 => \N__4778\,
            in3 => \N__6140\,
            lcout => \U712_CHIP_RAM.N_114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__6694\,
            in1 => \N__4763\,
            in2 => \_gnd_net_\,
            in3 => \N__4743\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLE_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI7Q5U5_0_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6415\,
            in1 => \N__5678\,
            in2 => \_gnd_net_\,
            in3 => \N__6693\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101000100000"
        )
    port map (
            in0 => \N__7294\,
            in1 => \N__5696\,
            in2 => \N__4706\,
            in3 => \N__6264\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5261\,
            in1 => \N__4702\,
            in2 => \N__5215\,
            in3 => \N__4878\,
            lcout => \U712_REG_SM.N_151_0\,
            ltout => \U712_REG_SM.N_151_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_4_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7098\,
            in1 => \N__5563\,
            in2 => \N__4691\,
            in3 => \N__5533\,
            lcout => \U712_REG_SM.N_160_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5285\,
            in2 => \_gnd_net_\,
            in3 => \N__5320\,
            lcout => \U712_REG_SM.N_147_0\,
            ltout => \U712_REG_SM.N_147_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_0_2_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5209\,
            in1 => \N__5262\,
            in2 => \N__4934\,
            in3 => \N__4862\,
            lcout => \U712_REG_SM.N_161_0\,
            ltout => \U712_REG_SM.N_161_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4917\,
            in2 => \N__4904\,
            in3 => \N__7099\,
            lcout => \U712_REG_SM.N_165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4879\,
            in1 => \N__4900\,
            in2 => \_gnd_net_\,
            in3 => \N__4861\,
            lcout => \U712_REG_SM.N_187\,
            ltout => \U712_REG_SM.N_187_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIPBP14_2_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__5263\,
            in1 => \N__5210\,
            in2 => \N__4889\,
            in3 => \N__4886\,
            lcout => \U712_REG_SM.C1_SYNC_RNIPBP14Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_1_6_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__4880\,
            in1 => \N__5264\,
            in2 => \N__5216\,
            in3 => \N__4863\,
            lcout => \U712_REG_SM.N_174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010001010000"
        )
    port map (
            in0 => \N__6921\,
            in1 => \N__4832\,
            in2 => \N__6005\,
            in3 => \N__5447\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8421\,
            ce => 'H',
            sr => \N__9361\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111100011111100"
        )
    port map (
            in0 => \N__7006\,
            in1 => \N__4807\,
            in2 => \N__6032\,
            in3 => \N__6922\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8421\,
            ce => 'H',
            sr => \N__9361\
        );

    \CLK40C_obuf_RNO_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7007\,
            lcout => \CLK40_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5324\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8421\,
            ce => 'H',
            sr => \N__9361\
        );

    \U712_REG_SM.REGENn_1_ess_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__5265\,
            in1 => \N__5214\,
            in2 => \_gnd_net_\,
            in3 => \N__5162\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8424\,
            ce => \N__5975\,
            sr => \N__9355\
        );

    \U712_REG_SM.UDS_OUT_RNIUP9B_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5105\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5081\,
            lcout => \U712_REG_SM_un1_UDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_0_i_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__6890\,
            in1 => \N__5038\,
            in2 => \N__6830\,
            in3 => \N__5761\,
            lcout => \DRDDIR_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100000001"
        )
    port map (
            in0 => \N__9243\,
            in1 => \N__9133\,
            in2 => \N__9020\,
            in3 => \N__4985\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8386\,
            ce => \N__8271\,
            sr => \N__9403\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__4964\,
            in1 => \N__9244\,
            in2 => \_gnd_net_\,
            in3 => \N__9011\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8386\,
            ce => \N__8271\,
            sr => \N__9403\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7334\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5456\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6993\,
            in1 => \N__7333\,
            in2 => \_gnd_net_\,
            in3 => \N__6926\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000010011"
        )
    port map (
            in0 => \N__9207\,
            in1 => \N__8797\,
            in2 => \N__9125\,
            in3 => \N__8972\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA31_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9460\,
            in1 => \_gnd_net_\,
            in2 => \N__5459\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6016\,
            in2 => \_gnd_net_\,
            in3 => \N__5455\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000000"
        )
    port map (
            in0 => \N__6439\,
            in1 => \N__7332\,
            in2 => \N__6619\,
            in3 => \N__6661\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5426\,
            in2 => \N__5435\,
            in3 => \N__8804\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6701\,
            in1 => \N__5484\,
            in2 => \_gnd_net_\,
            in3 => \N__7312\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_97_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110100000001"
        )
    port map (
            in0 => \N__5465\,
            in1 => \N__5429\,
            in2 => \N__5432\,
            in3 => \N__9102\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111011"
        )
    port map (
            in0 => \N__9221\,
            in1 => \N__5427\,
            in2 => \N__6665\,
            in3 => \N__7311\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000010000"
        )
    port map (
            in0 => \N__5408\,
            in1 => \N__5369\,
            in2 => \N__7330\,
            in3 => \N__6278\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5JPD5_3_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5336\,
            in1 => \N__7429\,
            in2 => \_gnd_net_\,
            in3 => \N__6056\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000001"
        )
    port map (
            in0 => \N__5676\,
            in1 => \N__6514\,
            in2 => \N__6440\,
            in3 => \N__6700\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__9455\,
            in1 => \_gnd_net_\,
            in2 => \N__5489\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5643\,
            in1 => \N__7474\,
            in2 => \_gnd_net_\,
            in3 => \N__7440\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__6515\,
            in1 => \N__6147\,
            in2 => \N__6626\,
            in3 => \N__5644\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__7307\,
            in1 => \N__7439\,
            in2 => \N__6173\,
            in3 => \N__6096\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6513\,
            in1 => \N__7306\,
            in2 => \_gnd_net_\,
            in3 => \N__6594\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__5486\,
            in1 => \N__6242\,
            in2 => \N__5468\,
            in3 => \N__6038\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6512\,
            in1 => \N__6593\,
            in2 => \_gnd_net_\,
            in3 => \N__6146\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7417\,
            in1 => \N__6135\,
            in2 => \_gnd_net_\,
            in3 => \N__6054\,
            lcout => \U712_CHIP_RAM.N_52\,
            ltout => \U712_CHIP_RAM.N_52_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111110"
        )
    port map (
            in0 => \N__6506\,
            in1 => \N__6591\,
            in2 => \N__5684\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI7Q5U5_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6436\,
            in2 => \N__5681\,
            in3 => \N__5677\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_90_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQU7BE_0_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__9454\,
            in1 => \N__6195\,
            in2 => \N__5654\,
            in3 => \N__5651\,
            lcout => \U712_CHIP_RAM.N_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111111001100"
        )
    port map (
            in0 => \N__6265\,
            in1 => \N__5611\,
            in2 => \N__6527\,
            in3 => \N__5495\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8409\,
            ce => 'H',
            sr => \N__9367\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000011"
        )
    port map (
            in0 => \N__6592\,
            in1 => \N__6507\,
            in2 => \N__6098\,
            in3 => \N__6239\,
            lcout => \U712_CHIP_RAM.N_124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5800\,
            in2 => \_gnd_net_\,
            in3 => \N__6528\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5581\,
            in1 => \N__5564\,
            in2 => \_gnd_net_\,
            in3 => \N__5534\,
            lcout => \U712_REG_SM.N_159_0\,
            ltout => \U712_REG_SM.N_159_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__7261\,
            in1 => \_gnd_net_\,
            in2 => \N__5504\,
            in3 => \N__5501\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8415\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000110011"
        )
    port map (
            in0 => \N__6172\,
            in1 => \N__6428\,
            in2 => \N__7450\,
            in3 => \N__6699\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7260\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6031\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8418\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_1_ess_RNO_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9450\,
            in2 => \_gnd_net_\,
            in3 => \N__5986\,
            lcout => \U712_REG_SM.N_180_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__5885\,
            in1 => \_gnd_net_\,
            in2 => \N__9265\,
            in3 => \N__9008\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8385\,
            ce => \N__8278\,
            sr => \N__9396\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__9007\,
            in1 => \N__9245\,
            in2 => \_gnd_net_\,
            in3 => \N__5843\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8385\,
            ce => \N__8278\,
            sr => \N__9396\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__8605\,
            in1 => \N__5927\,
            in2 => \N__5906\,
            in3 => \N__7487\,
            lcout => \U712_CHIP_RAM.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__7844\,
            in1 => \N__9097\,
            in2 => \N__8630\,
            in3 => \N__7724\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8606\,
            in1 => \N__5879\,
            in2 => \N__5867\,
            in3 => \N__5864\,
            lcout => \U712_CHIP_RAM.N_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000101"
        )
    port map (
            in0 => \N__6293\,
            in1 => \N__5837\,
            in2 => \N__5804\,
            in3 => \N__5746\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8615\,
            in2 => \_gnd_net_\,
            in3 => \N__6292\,
            lcout => \U712_CHIP_RAM.un6_CPU_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__6308\,
            in1 => \N__9456\,
            in2 => \N__6653\,
            in3 => \N__6371\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__6218\,
            in1 => \N__6272\,
            in2 => \N__8634\,
            in3 => \N__6171\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8399\,
            ce => \N__6377\,
            sr => \N__9368\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6505\,
            in2 => \_gnd_net_\,
            in3 => \N__6240\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6365\,
            in1 => \N__7354\,
            in2 => \N__6339\,
            in3 => \N__6645\,
            lcout => \U712_CHIP_RAM.N_46\,
            ltout => \U712_CHIP_RAM.N_46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6209\,
            in3 => \N__6503\,
            lcout => \U712_CHIP_RAM.N_116\,
            ltout => \U712_CHIP_RAM.N_116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_2_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6610\,
            in2 => \N__6176\,
            in3 => \N__6148\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIGB4P1_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__6149\,
            in1 => \N__7305\,
            in2 => \N__7442\,
            in3 => \N__6097\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6504\,
            in1 => \N__6611\,
            in2 => \N__6059\,
            in3 => \N__6055\,
            lcout => \U712_CHIP_RAM.N_96\,
            ltout => \U712_CHIP_RAM.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOF0DC_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6715\,
            in2 => \N__6704\,
            in3 => \N__6695\,
            lcout => \U712_CHIP_RAM.N_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6652\,
            in2 => \_gnd_net_\,
            in3 => \N__6366\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7430\,
            in1 => \N__6329\,
            in2 => \N__6629\,
            in3 => \N__7355\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__6612\,
            in1 => \N__6519\,
            in2 => \N__6443\,
            in3 => \N__6435\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9451\,
            in1 => \_gnd_net_\,
            in2 => \N__6380\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__6370\,
            in1 => \N__6304\,
            in2 => \_gnd_net_\,
            in3 => \N__9453\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__7432\,
            in1 => \N__7357\,
            in2 => \N__6341\,
            in3 => \N__7472\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6344\,
            in3 => \N__9452\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7431\,
            in1 => \N__7356\,
            in2 => \N__6340\,
            in3 => \N__7473\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010101100"
        )
    port map (
            in0 => \N__7100\,
            in1 => \N__6809\,
            in2 => \N__7085\,
            in3 => \N__7058\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8410\,
            ce => 'H',
            sr => \N__9356\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010111"
        )
    port map (
            in0 => \N__6951\,
            in1 => \N__7052\,
            in2 => \N__7031\,
            in3 => \N__6912\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__7256\,
            in1 => \N__7005\,
            in2 => \N__6959\,
            in3 => \N__6952\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8416\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6896\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6819\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__7493\,
            in1 => \N__9259\,
            in2 => \_gnd_net_\,
            in3 => \N__9010\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8384\,
            ce => \N__8292\,
            sr => \N__9384\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100011001101"
        )
    port map (
            in0 => \N__9009\,
            in1 => \N__7541\,
            in2 => \N__9269\,
            in3 => \N__9144\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8384\,
            ce => \N__8292\,
            sr => \N__9384\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7679\,
            in1 => \N__8591\,
            in2 => \N__9157\,
            in3 => \N__7730\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8593\,
            in1 => \N__7580\,
            in2 => \N__7559\,
            in3 => \N__7556\,
            lcout => \U712_CHIP_RAM.N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7604\,
            in1 => \N__8592\,
            in2 => \N__9158\,
            in3 => \N__7106\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__8594\,
            in1 => \N__7532\,
            in2 => \N__7511\,
            in3 => \N__7508\,
            lcout => \U712_CHIP_RAM.N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7685\,
            in1 => \N__8590\,
            in2 => \N__9156\,
            in3 => \N__7124\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__7481\,
            in1 => \N__9449\,
            in2 => \N__7454\,
            in3 => \N__7358\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7173\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7673\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8387\,
            ce => \N__8891\,
            sr => \N__9386\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7715\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8387\,
            ce => \N__8891\,
            sr => \N__9386\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7910\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8387\,
            ce => \N__8891\,
            sr => \N__9386\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7631\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8387\,
            ce => \N__8891\,
            sr => \N__9386\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7868\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8387\,
            ce => \N__8891\,
            sr => \N__9386\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7835\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8387\,
            ce => \N__8891\,
            sr => \N__9386\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7964\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8390\,
            ce => \N__7780\,
            sr => \N__9374\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7711\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8390\,
            ce => \N__7780\,
            sr => \N__9374\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8002\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8390\,
            ce => \N__7780\,
            sr => \N__9374\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7669\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8390\,
            ce => \N__7780\,
            sr => \N__9374\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7627\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8390\,
            ce => \N__7780\,
            sr => \N__9374\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__9264\,
            in1 => \N__8189\,
            in2 => \_gnd_net_\,
            in3 => \N__9017\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8400\,
            ce => \N__8291\,
            sr => \N__9369\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9263\,
            in1 => \N__9155\,
            in2 => \N__8825\,
            in3 => \N__9016\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8400\,
            ce => \N__8291\,
            sr => \N__9369\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8918\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8391\,
            ce => \N__7781\,
            sr => \N__9397\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7909\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8391\,
            ce => \N__7781\,
            sr => \N__9397\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7864\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8391\,
            ce => \N__7781\,
            sr => \N__9397\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7834\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8391\,
            ce => \N__7781\,
            sr => \N__9397\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7787\,
            in1 => \N__8631\,
            in2 => \N__9151\,
            in3 => \N__7937\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9458\,
            in2 => \_gnd_net_\,
            in3 => \N__7756\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNILUVG_1_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8092\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8081\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7745\,
            in1 => \N__8569\,
            in2 => \N__9161\,
            in3 => \N__7970\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__8234\,
            in1 => \N__8570\,
            in2 => \N__8213\,
            in3 => \N__8210\,
            lcout => \U712_CHIP_RAM.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8183\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8144\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8411\,
            ce => 'H',
            sr => \N__9370\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8093\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8411\,
            ce => 'H',
            sr => \N__9370\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__8009\,
            in1 => \N__9267\,
            in2 => \_gnd_net_\,
            in3 => \N__9018\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8392\,
            ce => \N__8293\,
            sr => \N__9408\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__8060\,
            in1 => \N__8629\,
            in2 => \N__8039\,
            in3 => \N__8015\,
            lcout => \U712_CHIP_RAM.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__9461\,
            in1 => \N__8753\,
            in2 => \_gnd_net_\,
            in3 => \N__8731\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8003\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8405\,
            ce => \N__8887\,
            sr => \N__9398\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7960\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8405\,
            ce => \N__8887\,
            sr => \N__9398\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8914\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8405\,
            ce => \N__8887\,
            sr => \N__9398\
        );

    \U712_CHIP_RAM.CASn_LC_16_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9160\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8393\,
            ce => 'H',
            sr => \N__9411\
        );

    \U712_CHIP_RAM.WEn_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9019\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8401\,
            ce => 'H',
            sr => \N__9410\
        );

    \U712_CHIP_RAM.RASn_LC_16_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9268\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8401\,
            ce => 'H',
            sr => \N__9410\
        );

    \U712_CHIP_RAM.CRCSn_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8824\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8406\,
            ce => 'H',
            sr => \N__9409\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8732\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8406\,
            ce => 'H',
            sr => \N__9409\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8659\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8747\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8406\,
            ce => 'H',
            sr => \N__9409\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__8720\,
            in1 => \N__8926\,
            in2 => \N__8705\,
            in3 => \N__8632\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8412\,
            ce => \N__8294\,
            sr => \N__9404\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__8675\,
            in1 => \N__8927\,
            in2 => \N__8660\,
            in3 => \N__8633\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8412\,
            ce => \N__8294\,
            sr => \N__9404\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__9266\,
            in1 => \N__9159\,
            in2 => \_gnd_net_\,
            in3 => \N__9015\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Sep 11 2025 19:59:55

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U111_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U111_TOP
entity U111_TOP is
port (
    D_LM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UM_AMIGA : inout std_logic_vector(7 downto 0);
    D_LL_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_AMIGA : inout std_logic_vector(7 downto 0);
    D_LL_040 : inout std_logic_vector(7 downto 0);
    D_UU_040 : inout std_logic_vector(7 downto 0);
    D_LM_040 : inout std_logic_vector(7 downto 0);
    D_UM_040 : inout std_logic_vector(7 downto 0);
    A_AMIGA : out std_logic_vector(1 downto 0);
    A_040 : in std_logic_vector(1 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    TBIn : in std_logic;
    TEAn : in std_logic;
    TSn : out std_logic;
    RESETn : in std_logic;
    CLKRAMA : out std_logic;
    PORTSIZE : in std_logic;
    DMAAn : out std_logic;
    TEA_CPUn : out std_logic;
    LBENn : in std_logic;
    CLK40B : out std_logic;
    TBI_CPUn : out std_logic;
    TAn : inout std_logic;
    CPUBGn : out std_logic;
    BUFENn : out std_logic;
    RnW : in std_logic;
    CLK80_CPU : out std_logic;
    BUFDIR : out std_logic;
    TCI_CPUn : out std_logic;
    TS_CPUn : inout std_logic;
    CLKRAMB : out std_logic;
    CLK40A : out std_logic;
    TCIn : in std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    BBn : in std_logic;
    TACKn : inout std_logic;
    BGn : in std_logic);
end U111_TOP;

-- Architecture of U111_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U111_TOP is

signal \N__9524\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2655\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \TAn_in\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U111_CYCLE_SM_A_AMIGA_0_i_1\ : std_logic;
signal \A_040_c_0\ : std_logic;
signal \A_AMIGA_c_0\ : std_logic;
signal \D_UM_040_in_2\ : std_logic;
signal \D_LL_040_in_2\ : std_logic;
signal \un1_D_UM_040_2\ : std_logic;
signal \D_UU_040_in_4\ : std_logic;
signal \D_LM_040_in_4\ : std_logic;
signal \un1_D_UU_040_4\ : std_logic;
signal \D_UM_040_in_4\ : std_logic;
signal \D_LL_040_in_4\ : std_logic;
signal \un1_D_UM_040_4\ : std_logic;
signal \D_LL_AMIGA_in_1\ : std_logic;
signal \un2_D_LL_AMIGA_1\ : std_logic;
signal \CPUBGn_c_i_0\ : std_logic;
signal \D_LL_AMIGA_in_5\ : std_logic;
signal \un2_D_LL_AMIGA_5\ : std_logic;
signal \D_LL_AMIGA_in_7\ : std_logic;
signal \un2_D_LL_AMIGA_7\ : std_logic;
signal \A_040_c_1\ : std_logic;
signal \D_LM_AMIGA_in_5\ : std_logic;
signal \N_108\ : std_logic;
signal \D_LM_AMIGA_in_3\ : std_logic;
signal \N_110\ : std_logic;
signal \D_LM_AMIGA_in_2\ : std_logic;
signal \N_111\ : std_logic;
signal \D_UM_040_in_6\ : std_logic;
signal \D_LL_040_in_6\ : std_logic;
signal \un1_D_UM_040_6\ : std_logic;
signal \D_UU_040_in_0\ : std_logic;
signal \D_LM_040_in_0\ : std_logic;
signal \un1_D_UU_040_0\ : std_logic;
signal \D_UU_040_in_6\ : std_logic;
signal \D_LM_040_in_6\ : std_logic;
signal \un1_D_UU_040_6\ : std_logic;
signal \D_LL_AMIGA_in_4\ : std_logic;
signal \un2_D_LL_AMIGA_4\ : std_logic;
signal \D_LL_AMIGA_in_2\ : std_logic;
signal \un2_D_LL_AMIGA_2\ : std_logic;
signal \D_LL_040_in_0\ : std_logic;
signal \D_UM_040_in_0\ : std_logic;
signal \un1_D_UM_040_0\ : std_logic;
signal \D_LM_AMIGA_in_1\ : std_logic;
signal \N_112\ : std_logic;
signal \N_96\ : std_logic;
signal \N_94_i\ : std_logic;
signal \BBn_c\ : std_logic;
signal \BUFDIR_c\ : std_logic;
signal \GB_BUFFER_CLK40_THRU_CO\ : std_logic;
signal \U111_CYCLE_SM.N_141\ : std_logic;
signal \U111_CYCLE_SM.TS_ENZ0\ : std_logic;
signal \INVU111_CYCLE_SM.TS_OUTC_net\ : std_logic;
signal \D_LM_AMIGA_in_7\ : std_logic;
signal \N_106\ : std_logic;
signal \D_LM_AMIGA_in_6\ : std_logic;
signal \N_107\ : std_logic;
signal \D_UM_040_in_3\ : std_logic;
signal \D_LL_040_in_3\ : std_logic;
signal \un1_D_UM_040_3\ : std_logic;
signal \D_LL_AMIGA_in_3\ : std_logic;
signal \un2_D_LL_AMIGA_3\ : std_logic;
signal \LBENn_c_i\ : std_logic;
signal \D_LM_AMIGA_in_0\ : std_logic;
signal \un2_D_LM_AMIGA_0\ : std_logic;
signal \U111_CYCLE_SM.A2_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.N_179\ : std_logic;
signal \U111_CYCLE_SM.N_179_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_101_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_98\ : std_logic;
signal \U111_CYCLE_SM.N_10\ : std_logic;
signal \U111_CYCLE_SM.N_101\ : std_logic;
signal \U111_CYCLE_SM.N_12_i_1_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_55\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNTZ0Z_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNTZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.LW_TRANSZ0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\ : std_logic;
signal \PORTSIZE_c\ : std_logic;
signal \TS_CPUn_in\ : std_logic;
signal \D_LM_AMIGA_in_4\ : std_logic;
signal \N_109\ : std_logic;
signal \D_UU_040_in_2\ : std_logic;
signal \D_LM_040_in_2\ : std_logic;
signal \un1_D_UU_040_2\ : std_logic;
signal \D_UU_AMIGA_in_2\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\ : std_logic;
signal \N_118\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\ : std_logic;
signal \D_UU_AMIGA_in_4\ : std_logic;
signal \N_116\ : std_logic;
signal \D_UU_AMIGA_in_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\ : std_logic;
signal \N_113\ : std_logic;
signal \D_LM_040_in_3\ : std_logic;
signal \D_UU_040_in_3\ : std_logic;
signal \un1_D_UU_040_3\ : std_logic;
signal \D_UU_AMIGA_in_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\ : std_logic;
signal \N_115\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_i_i_o2_0_5_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\ : std_logic;
signal \U111_CYCLE_SM.PORT_MISMATCHZ0\ : std_logic;
signal \U111_CYCLE_SM.BURSTZ0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_a3_2_0_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_133\ : std_logic;
signal \U111_CYCLE_SM.N_131\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_2_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.TS_DELAYZ0\ : std_logic;
signal \U111_CYCLE_SM.un4_TS_OUT_i_0_cascade_\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\ : std_logic;
signal \U111_CYCLE_SM.N_99_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\ : std_logic;
signal \U111_CYCLE_SM.N_51\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\ : std_logic;
signal \D_LM_040_in_1\ : std_logic;
signal \D_UU_040_in_1\ : std_logic;
signal \un1_D_UU_040_1\ : std_logic;
signal \TS_OUT\ : std_logic;
signal \TSnz\ : std_logic;
signal \D_LM_040_in_7\ : std_logic;
signal \D_UU_040_in_7\ : std_logic;
signal \un1_D_UU_040_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\ : std_logic;
signal \D_UU_AMIGA_in_6\ : std_logic;
signal \N_114\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \BGn_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0\ : std_logic;
signal \U111_CYCLE_SM_OFFBOARD_EN_0\ : std_logic;
signal \U111_CYCLE_SM.un4_TS_OUT_i_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U111_CYCLE_SM.N_99\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_99_i\ : std_logic;
signal \D_UM_040_in_1\ : std_logic;
signal \D_LL_040_in_1\ : std_logic;
signal \un1_D_UM_040_1\ : std_logic;
signal \D_UU_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\ : std_logic;
signal \N_119\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\ : std_logic;
signal \D_UM_AMIGA_in_4\ : std_logic;
signal \un1_D_UM_AMIGA_4\ : std_logic;
signal \CLK80\ : std_logic;
signal \GB_BUFFER_CLK80_THRU_CO\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\ : std_logic;
signal \D_UU_AMIGA_in_0\ : std_logic;
signal \un1_D_UU_AMIGA_0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\ : std_logic;
signal \D_UU_AMIGA_in_3\ : std_logic;
signal \N_117\ : std_logic;
signal \D_LL_AMIGA_in_0\ : std_logic;
signal \un2_D_LL_AMIGA_0\ : std_logic;
signal \TBIn_c\ : std_logic;
signal \U111_CYCLE_SM_TBI_CPUn_0_i\ : std_logic;
signal \D_LL_AMIGA_in_6\ : std_logic;
signal \un2_D_LL_AMIGA_6\ : std_logic;
signal \un1_D_UM_AMIGA_2\ : std_logic;
signal \un1_D_UM_AMIGA_0\ : std_logic;
signal \TEAn_c\ : std_logic;
signal \U111_CYCLE_SM_TEA_CPUn_0_i\ : std_logic;
signal \D_UM_AMIGA_in_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\ : std_logic;
signal \D_UM_AMIGA_in_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\ : std_logic;
signal \CLK40\ : std_logic;
signal \U111_CYCLE_SM.N_99_i_0\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\ : std_logic;
signal \D_UM_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\ : std_logic;
signal \un1_D_UM_AMIGA_1\ : std_logic;
signal \U111_CYCLE_SM.TA_DISZ0\ : std_logic;
signal \N_64\ : std_logic;
signal \TCIn_c\ : std_logic;
signal \LBENn_c\ : std_logic;
signal \U111_CYCLE_SM_TCI_CPUn_0_i\ : std_logic;
signal \D_UM_AMIGA_in_3\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\ : std_logic;
signal \un1_D_UM_AMIGA_3\ : std_logic;
signal \D_LL_040_in_7\ : std_logic;
signal \D_UM_040_in_7\ : std_logic;
signal \un1_D_UM_040_7\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\ : std_logic;
signal \D_UM_AMIGA_in_7\ : std_logic;
signal \un1_D_UM_AMIGA_7\ : std_logic;
signal \D_LM_040_in_5\ : std_logic;
signal \D_UU_040_in_5\ : std_logic;
signal \un1_D_UU_040_5\ : std_logic;
signal \D_UM_040_in_5\ : std_logic;
signal \D_LL_040_in_5\ : std_logic;
signal \U111_CYCLE_SM.FLIP_WORDZ0\ : std_logic;
signal \un1_D_UM_040_5\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\ : std_logic;
signal \D_UM_AMIGA_in_5\ : std_logic;
signal \un1_D_UM_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\ : std_logic;
signal \CPUBGn_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \N_60_i\ : std_logic;
signal \U111_CYCLE_SM.LATCH_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\ : std_logic;
signal \D_UM_AMIGA_in_6\ : std_logic;
signal \un1_D_UM_AMIGA_6\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \LBENn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \CPUBGn_wire\ : std_logic;
signal \TEA_CPUn_wire\ : std_logic;
signal \A_040_wire\ : std_logic_vector(1 downto 0);
signal \A_AMIGA_wire\ : std_logic_vector(1 downto 0);
signal \CLK40B_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \BUFDIR_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \CLKRAMB_wire\ : std_logic;
signal \TEAn_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \CLK80_CPU_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \BGn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \TBI_CPUn_wire\ : std_logic;
signal \CLK40A_wire\ : std_logic;
signal \CLKRAMA_wire\ : std_logic;
signal \TCI_CPUn_wire\ : std_logic;
signal \BBn_wire\ : std_logic;
signal \DMAAn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \pll_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \LBENn_wire\ <= LBENn;
    TSn <= \TSn_wire\;
    CPUBGn <= \CPUBGn_wire\;
    TEA_CPUn <= \TEA_CPUn_wire\;
    \A_040_wire\ <= A_040;
    A_AMIGA <= \A_AMIGA_wire\;
    CLK40B <= \CLK40B_wire\;
    \TBIn_wire\ <= TBIn;
    BUFDIR <= \BUFDIR_wire\;
    \SIZ_wire\ <= SIZ;
    CLKRAMB <= \CLKRAMB_wire\;
    \TEAn_wire\ <= TEAn;
    BUFENn <= \BUFENn_wire\;
    CLK80_CPU <= \CLK80_CPU_wire\;
    \PORTSIZE_wire\ <= PORTSIZE;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    \BGn_wire\ <= BGn;
    \TCIn_wire\ <= TCIn;
    TBI_CPUn <= \TBI_CPUn_wire\;
    CLK40A <= \CLK40A_wire\;
    CLKRAMA <= \CLKRAMA_wire\;
    TCI_CPUn <= \TCI_CPUn_wire\;
    \BBn_wire\ <= BBn;
    DMAAn <= \DMAAn_wire\;
    \RnW_wire\ <= RnW;
    \pll_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_pll\ : PLL40_2F
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            SCLK => '0',
            PLLOUTGLOBALA => \CLK80\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALB => \CLK40\,
            SDI => '0',
            PLLOUTCOREA => OPEN,
            BYPASS => '0',
            RESETB => \N__5553\,
            PLLOUTCOREB => OPEN,
            LOCK => OPEN,
            SDO => OPEN,
            EXTFEEDBACK => '0',
            DYNAMICDELAY => \pll_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__9524\
        );

    \pll_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__9524\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \LBENn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9508\,
            DIN => \N__9507\,
            DOUT => \N__9506\,
            PACKAGEPIN => \LBENn_wire\
        );

    \LBENn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9508\,
            PADOUT => \N__9507\,
            PADIN => \N__9506\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \LBENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9499\,
            DIN => \N__9498\,
            DOUT => \N__9497\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9499\,
            PADOUT => \N__9498\,
            PADIN => \N__9497\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2763\,
            DIN0 => OPEN,
            DOUT0 => \N__5760\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9490\,
            DIN => \N__9489\,
            DOUT => \N__9488\,
            PACKAGEPIN => D_UM_040(3)
        );

    \D_UM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9490\,
            PADOUT => \N__9489\,
            PADIN => \N__9488\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7637\,
            DIN0 => \D_UM_040_in_3\,
            DOUT0 => \N__8556\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9481\,
            DIN => \N__9480\,
            DOUT => \N__9479\,
            PACKAGEPIN => TAn
        );

    \TAn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9481\,
            PADOUT => \N__9480\,
            PADIN => \N__9479\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6918\,
            DIN0 => \TAn_in\,
            DOUT0 => \N__5205\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9472\,
            DIN => \N__9471\,
            DOUT => \N__9470\,
            PACKAGEPIN => D_LL_AMIGA(1)
        );

    \D_LL_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9472\,
            PADOUT => \N__9471\,
            PADIN => \N__9470\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5435\,
            DIN0 => \D_LL_AMIGA_in_1\,
            DOUT0 => \N__6099\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9463\,
            DIN => \N__9462\,
            DOUT => \N__9461\,
            PACKAGEPIN => D_UU_AMIGA(5)
        );

    \D_UU_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9463\,
            PADOUT => \N__9462\,
            PADIN => \N__9461\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5475\,
            DIN0 => \D_UU_AMIGA_in_5\,
            DOUT0 => \N__8304\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9454\,
            DIN => \N__9453\,
            DOUT => \N__9452\,
            PACKAGEPIN => D_UU_040(6)
        );

    \D_UU_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9454\,
            PADOUT => \N__9453\,
            PADIN => \N__9452\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7646\,
            DIN0 => \D_UU_040_in_6\,
            DOUT0 => \N__5574\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUBGn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9445\,
            DIN => \N__9444\,
            DOUT => \N__9443\,
            PACKAGEPIN => \CPUBGn_wire\
        );

    \CPUBGn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9445\,
            PADOUT => \N__9444\,
            PADIN => \N__9443\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7824\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9436\,
            DIN => \N__9435\,
            DOUT => \N__9434\,
            PACKAGEPIN => D_LL_040(7)
        );

    \D_LL_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9436\,
            PADOUT => \N__9435\,
            PADIN => \N__9434\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7528\,
            DIN0 => \D_LL_040_in_7\,
            DOUT0 => \N__2706\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9427\,
            DIN => \N__9426\,
            DOUT => \N__9425\,
            PACKAGEPIN => D_LL_AMIGA(4)
        );

    \D_LL_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9427\,
            PADOUT => \N__9426\,
            PADIN => \N__9425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5434\,
            DIN0 => \D_LL_AMIGA_in_4\,
            DOUT0 => \N__2865\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9418\,
            DIN => \N__9417\,
            DOUT => \N__9416\,
            PACKAGEPIN => D_UM_AMIGA(3)
        );

    \D_UM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9418\,
            PADOUT => \N__9417\,
            PADIN => \N__9416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5431\,
            DIN0 => \D_UM_AMIGA_in_3\,
            DOUT0 => \N__3921\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9409\,
            DIN => \N__9408\,
            DOUT => \N__9407\,
            PACKAGEPIN => D_UU_040(3)
        );

    \D_UU_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9409\,
            PADOUT => \N__9408\,
            PADIN => \N__9407\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7480\,
            DIN0 => \D_UU_040_in_3\,
            DOUT0 => \N__6678\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEA_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9400\,
            DIN => \N__9399\,
            DOUT => \N__9398\,
            PACKAGEPIN => \TEA_CPUn_wire\
        );

    \TEA_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9400\,
            PADOUT => \N__9399\,
            PADIN => \N__9398\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6432\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9391\,
            DIN => \N__9390\,
            DOUT => \N__9389\,
            PACKAGEPIN => \A_040_wire\(1)
        );

    \A_040_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9391\,
            PADOUT => \N__9390\,
            PADIN => \N__9389\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9382\,
            DIN => \N__9381\,
            DOUT => \N__9380\,
            PACKAGEPIN => D_LM_AMIGA(3)
        );

    \D_LM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9382\,
            PADOUT => \N__9381\,
            PADIN => \N__9380\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5266\,
            DIN0 => \D_LM_AMIGA_in_3\,
            DOUT0 => \N__4413\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9373\,
            DIN => \N__9372\,
            DOUT => \N__9371\,
            PACKAGEPIN => D_LM_040(0)
        );

    \D_LM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9373\,
            PADOUT => \N__9372\,
            PADIN => \N__9371\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7529\,
            DIN0 => \D_LM_040_in_0\,
            DOUT0 => \N__3834\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9364\,
            DIN => \N__9363\,
            DOUT => \N__9362\,
            PACKAGEPIN => D_UM_AMIGA(6)
        );

    \D_UM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9364\,
            PADOUT => \N__9363\,
            PADIN => \N__9362\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5457\,
            DIN0 => \D_UM_AMIGA_in_6\,
            DOUT0 => \N__3294\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9355\,
            DIN => \N__9354\,
            DOUT => \N__9353\,
            PACKAGEPIN => D_LM_AMIGA(4)
        );

    \D_LM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9355\,
            PADOUT => \N__9354\,
            PADIN => \N__9353\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5326\,
            DIN0 => \D_LM_AMIGA_in_4\,
            DOUT0 => \N__2940\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9346\,
            DIN => \N__9345\,
            DOUT => \N__9344\,
            PACKAGEPIN => \A_AMIGA_wire\(1)
        );

    \A_AMIGA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9346\,
            PADOUT => \N__9345\,
            PADIN => \N__9344\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3078\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9337\,
            DIN => \N__9336\,
            DOUT => \N__9335\,
            PACKAGEPIN => D_LM_040(7)
        );

    \D_LM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9337\,
            PADOUT => \N__9336\,
            PADIN => \N__9335\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7600\,
            DIN0 => \D_LM_040_in_7\,
            DOUT0 => \N__4035\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9328\,
            DIN => \N__9327\,
            DOUT => \N__9326\,
            PACKAGEPIN => D_UM_040(4)
        );

    \D_UM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9328\,
            PADOUT => \N__9327\,
            PADIN => \N__9326\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7481\,
            DIN0 => \D_UM_040_in_4\,
            DOUT0 => \N__5892\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9319\,
            DIN => \N__9318\,
            DOUT => \N__9317\,
            PACKAGEPIN => \CLK40B_wire\
        );

    \CLK40B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9319\,
            PADOUT => \N__9318\,
            PADIN => \N__9317\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3552\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9310\,
            DIN => \N__9309\,
            DOUT => \N__9308\,
            PACKAGEPIN => D_UU_AMIGA(0)
        );

    \D_UU_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9310\,
            PADOUT => \N__9309\,
            PADIN => \N__9308\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5465\,
            DIN0 => \D_UU_AMIGA_in_0\,
            DOUT0 => \N__3210\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9301\,
            DIN => \N__9300\,
            DOUT => \N__9299\,
            PACKAGEPIN => D_UM_040(1)
        );

    \D_UM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9301\,
            PADOUT => \N__9300\,
            PADIN => \N__9299\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7479\,
            DIN0 => \D_UM_040_in_1\,
            DOUT0 => \N__6966\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9292\,
            DIN => \N__9291\,
            DOUT => \N__9290\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9292\,
            PADOUT => \N__9291\,
            PADIN => \N__9290\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TBIn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9283\,
            DIN => \N__9282\,
            DOUT => \N__9281\,
            PACKAGEPIN => D_LL_040(4)
        );

    \D_LL_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9283\,
            PADOUT => \N__9282\,
            PADIN => \N__9281\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7633\,
            DIN0 => \D_LL_040_in_4\,
            DOUT0 => \N__3099\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9274\,
            DIN => \N__9273\,
            DOUT => \N__9272\,
            PACKAGEPIN => D_LL_AMIGA(7)
        );

    \D_LL_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9274\,
            PADOUT => \N__9273\,
            PADIN => \N__9272\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5395\,
            DIN0 => \D_LL_AMIGA_in_7\,
            DOUT0 => \N__8535\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9265\,
            DIN => \N__9264\,
            DOUT => \N__9263\,
            PACKAGEPIN => D_UU_AMIGA(7)
        );

    \D_UU_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9265\,
            PADOUT => \N__9264\,
            PADIN => \N__9263\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5467\,
            DIN0 => \D_UU_AMIGA_in_7\,
            DOUT0 => \N__5646\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9256\,
            DIN => \N__9255\,
            DOUT => \N__9254\,
            PACKAGEPIN => \BUFDIR_wire\
        );

    \BUFDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9256\,
            PADOUT => \N__9255\,
            PADIN => \N__9254\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3582\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9247\,
            DIN => \N__9246\,
            DOUT => \N__9245\,
            PACKAGEPIN => D_UU_040(4)
        );

    \D_UU_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9247\,
            PADOUT => \N__9246\,
            PADIN => \N__9245\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7614\,
            DIN0 => \D_UU_040_in_4\,
            DOUT0 => \N__4515\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9238\,
            DIN => \N__9237\,
            DOUT => \N__9236\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9238\,
            PADOUT => \N__9237\,
            PADIN => \N__9236\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9229\,
            DIN => \N__9228\,
            DOUT => \N__9227\,
            PACKAGEPIN => D_LL_040(1)
        );

    \D_LL_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9229\,
            PADOUT => \N__9228\,
            PADIN => \N__9227\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7632\,
            DIN0 => \D_LL_040_in_1\,
            DOUT0 => \N__2787\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9220\,
            DIN => \N__9219\,
            DOUT => \N__9218\,
            PACKAGEPIN => D_UM_AMIGA(5)
        );

    \D_UM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9220\,
            PADOUT => \N__9219\,
            PADIN => \N__9218\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5466\,
            DIN0 => \D_UM_AMIGA_in_5\,
            DOUT0 => \N__7980\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9211\,
            DIN => \N__9210\,
            DOUT => \N__9209\,
            PACKAGEPIN => D_UU_040(1)
        );

    \D_UU_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9211\,
            PADOUT => \N__9210\,
            PADIN => \N__9209\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7653\,
            DIN0 => \D_UU_040_in_1\,
            DOUT0 => \N__5976\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9202\,
            DIN => \N__9201\,
            DOUT => \N__9200\,
            PACKAGEPIN => D_LM_AMIGA(1)
        );

    \D_LM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9202\,
            PADOUT => \N__9201\,
            PADIN => \N__9200\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5323\,
            DIN0 => \D_LM_AMIGA_in_1\,
            DOUT0 => \N__5019\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9193\,
            DIN => \N__9192\,
            DOUT => \N__9191\,
            PACKAGEPIN => D_LM_040(2)
        );

    \D_LM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9193\,
            PADOUT => \N__9192\,
            PADIN => \N__9191\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7495\,
            DIN0 => \D_LM_040_in_2\,
            DOUT0 => \N__3375\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9184\,
            DIN => \N__9183\,
            DOUT => \N__9182\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9184\,
            PADOUT => \N__9183\,
            PADIN => \N__9182\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3861\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__2685\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9175\,
            DIN => \N__9174\,
            DOUT => \N__9173\,
            PACKAGEPIN => D_UM_040(2)
        );

    \D_UM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9175\,
            PADOUT => \N__9174\,
            PADIN => \N__9173\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7558\,
            DIN0 => \D_UM_040_in_2\,
            DOUT0 => \N__6537\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9166\,
            DIN => \N__9165\,
            DOUT => \N__9164\,
            PACKAGEPIN => \CLKRAMB_wire\
        );

    \CLKRAMB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9166\,
            PADOUT => \N__9165\,
            PADIN => \N__9164\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5856\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9157\,
            DIN => \N__9156\,
            DOUT => \N__9155\,
            PACKAGEPIN => D_LL_AMIGA(2)
        );

    \D_LL_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9157\,
            PADOUT => \N__9156\,
            PADIN => \N__9155\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5285\,
            DIN0 => \D_LL_AMIGA_in_2\,
            DOUT0 => \N__3027\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9148\,
            DIN => \N__9147\,
            DOUT => \N__9146\,
            PACKAGEPIN => D_UU_AMIGA(2)
        );

    \D_UU_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9148\,
            PADOUT => \N__9147\,
            PADIN => \N__9146\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5464\,
            DIN0 => \D_UU_AMIGA_in_2\,
            DOUT0 => \N__4677\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEAn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9139\,
            DIN => \N__9138\,
            DOUT => \N__9137\,
            PACKAGEPIN => \TEAn_wire\
        );

    \TEAn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9139\,
            PADOUT => \N__9138\,
            PADIN => \N__9137\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TEAn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9130\,
            DIN => \N__9129\,
            DOUT => \N__9128\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9130\,
            PADOUT => \N__9129\,
            PADIN => \N__9128\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3624\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9121\,
            DIN => \N__9120\,
            DOUT => \N__9119\,
            PACKAGEPIN => D_LL_040(6)
        );

    \D_LL_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9121\,
            PADOUT => \N__9120\,
            PADIN => \N__9119\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7630\,
            DIN0 => \D_LL_040_in_6\,
            DOUT0 => \N__6558\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9112\,
            DIN => \N__9111\,
            DOUT => \N__9110\,
            PACKAGEPIN => D_LL_AMIGA(5)
        );

    \D_LL_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9112\,
            PADOUT => \N__9111\,
            PADIN => \N__9110\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5398\,
            DIN0 => \D_LL_AMIGA_in_5\,
            DOUT0 => \N__8268\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9103\,
            DIN => \N__9102\,
            DOUT => \N__9101\,
            PACKAGEPIN => D_UM_AMIGA(0)
        );

    \D_UM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9103\,
            PADOUT => \N__9102\,
            PADIN => \N__9101\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5325\,
            DIN0 => \D_UM_AMIGA_in_0\,
            DOUT0 => \N__3693\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9094\,
            DIN => \N__9093\,
            DOUT => \N__9092\,
            PACKAGEPIN => D_UU_040(2)
        );

    \D_UU_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9094\,
            PADOUT => \N__9093\,
            PADIN => \N__9092\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7527\,
            DIN0 => \D_UU_040_in_2\,
            DOUT0 => \N__4590\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9085\,
            DIN => \N__9084\,
            DOUT => \N__9083\,
            PACKAGEPIN => D_LM_AMIGA(2)
        );

    \D_LM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9085\,
            PADOUT => \N__9084\,
            PADIN => \N__9083\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5324\,
            DIN0 => \D_LM_AMIGA_in_2\,
            DOUT0 => \N__4725\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TS_CPUn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9076\,
            DIN => \N__9075\,
            DOUT => \N__9074\,
            PACKAGEPIN => TS_CPUn
        );

    \TS_CPUn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9076\,
            PADOUT => \N__9075\,
            PADIN => \N__9074\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7820\,
            DIN0 => \TS_CPUn_in\,
            DOUT0 => \N__5724\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK80_CPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9067\,
            DIN => \N__9066\,
            DOUT => \N__9065\,
            PACKAGEPIN => \CLK80_CPU_wire\
        );

    \CLK80_CPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9067\,
            PADOUT => \N__9066\,
            PADIN => \N__9065\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5855\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9058\,
            DIN => \N__9057\,
            DOUT => \N__9056\,
            PACKAGEPIN => D_LL_040(3)
        );

    \D_LL_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9058\,
            PADOUT => \N__9057\,
            PADIN => \N__9056\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7634\,
            DIN0 => \D_LL_040_in_3\,
            DOUT0 => \N__3885\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9049\,
            DIN => \N__9048\,
            DOUT => \N__9047\,
            PACKAGEPIN => D_LM_040(1)
        );

    \D_LM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9049\,
            PADOUT => \N__9048\,
            PADIN => \N__9047\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7494\,
            DIN0 => \D_LM_040_in_1\,
            DOUT0 => \N__3663\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9040\,
            DIN => \N__9039\,
            DOUT => \N__9038\,
            PACKAGEPIN => D_UM_AMIGA(7)
        );

    \D_UM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9040\,
            PADOUT => \N__9039\,
            PADIN => \N__9038\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5432\,
            DIN0 => \D_UM_AMIGA_in_7\,
            DOUT0 => \N__8463\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9031\,
            DIN => \N__9030\,
            DOUT => \N__9029\,
            PACKAGEPIN => D_LM_AMIGA(7)
        );

    \D_LM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9031\,
            PADOUT => \N__9030\,
            PADIN => \N__9029\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5372\,
            DIN0 => \D_LM_AMIGA_in_7\,
            DOUT0 => \N__5706\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9022\,
            DIN => \N__9021\,
            DOUT => \N__9020\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9022\,
            PADOUT => \N__9021\,
            PADIN => \N__9020\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PORTSIZE_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9013\,
            DIN => \N__9012\,
            DOUT => \N__9011\,
            PACKAGEPIN => \A_AMIGA_wire\(0)
        );

    \A_AMIGA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9013\,
            PADOUT => \N__9012\,
            PADIN => \N__9011\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3054\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9004\,
            DIN => \N__9003\,
            DOUT => \N__9002\,
            PACKAGEPIN => D_LM_040(4)
        );

    \D_LM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9004\,
            PADOUT => \N__9003\,
            PADIN => \N__9002\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7610\,
            DIN0 => \D_LM_040_in_4\,
            DOUT0 => \N__4764\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8995\,
            DIN => \N__8994\,
            DOUT => \N__8993\,
            PACKAGEPIN => D_UM_040(7)
        );

    \D_UM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8995\,
            PADOUT => \N__8994\,
            PADIN => \N__8993\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7636\,
            DIN0 => \D_UM_040_in_7\,
            DOUT0 => \N__8382\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8986\,
            DIN => \N__8985\,
            DOUT => \N__8984\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8986\,
            PADOUT => \N__8985\,
            PADIN => \N__8984\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8977\,
            DIN => \N__8976\,
            DOUT => \N__8975\,
            PACKAGEPIN => D_UU_AMIGA(1)
        );

    \D_UU_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8977\,
            PADOUT => \N__8976\,
            PADIN => \N__8975\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5430\,
            DIN0 => \D_UU_AMIGA_in_1\,
            DOUT0 => \N__4968\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8968\,
            DIN => \N__8967\,
            DOUT => \N__8966\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8968\,
            PADOUT => \N__8967\,
            PADIN => \N__8966\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3556\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8959\,
            DIN => \N__8958\,
            DOUT => \N__8957\,
            PACKAGEPIN => D_UM_040(0)
        );

    \D_UM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8959\,
            PADOUT => \N__8958\,
            PADIN => \N__8957\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7559\,
            DIN0 => \D_UM_040_in_0\,
            DOUT0 => \N__6525\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8950\,
            DIN => \N__8949\,
            DOUT => \N__8948\,
            PACKAGEPIN => D_LL_AMIGA(0)
        );

    \D_LL_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8950\,
            PADOUT => \N__8949\,
            PADIN => \N__8948\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5462\,
            DIN0 => \D_LL_AMIGA_in_0\,
            DOUT0 => \N__3753\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8941\,
            DIN => \N__8940\,
            DOUT => \N__8939\,
            PACKAGEPIN => D_UU_AMIGA(4)
        );

    \D_UU_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8941\,
            PADOUT => \N__8940\,
            PADIN => \N__8939\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5463\,
            DIN0 => \D_UU_AMIGA_in_4\,
            DOUT0 => \N__2901\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8932\,
            DIN => \N__8931\,
            DOUT => \N__8930\,
            PACKAGEPIN => D_UU_040(7)
        );

    \D_UU_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8932\,
            PADOUT => \N__8931\,
            PADIN => \N__8930\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7645\,
            DIN0 => \D_UU_040_in_7\,
            DOUT0 => \N__4434\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8923\,
            DIN => \N__8922\,
            DOUT => \N__8921\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8923\,
            PADOUT => \N__8922\,
            PADIN => \N__8921\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BGn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8914\,
            DIN => \N__8913\,
            DOUT => \N__8912\,
            PACKAGEPIN => \BGn_wire\
        );

    \BGn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8914\,
            PADOUT => \N__8913\,
            PADIN => \N__8912\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BGn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8905\,
            DIN => \N__8904\,
            DOUT => \N__8903\,
            PACKAGEPIN => D_LL_040(0)
        );

    \D_LL_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8905\,
            PADOUT => \N__8904\,
            PADIN => \N__8903\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7635\,
            DIN0 => \D_LL_040_in_0\,
            DOUT0 => \N__6639\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8896\,
            DIN => \N__8895\,
            DOUT => \N__8894\,
            PACKAGEPIN => D_UM_AMIGA(2)
        );

    \D_UM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8896\,
            PADOUT => \N__8895\,
            PADIN => \N__8894\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5327\,
            DIN0 => \D_UM_AMIGA_in_2\,
            DOUT0 => \N__2982\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8887\,
            DIN => \N__8886\,
            DOUT => \N__8885\,
            PACKAGEPIN => D_UU_040(0)
        );

    \D_UU_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8887\,
            PADOUT => \N__8886\,
            PADIN => \N__8885\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7644\,
            DIN0 => \D_UU_040_in_0\,
            DOUT0 => \N__6768\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8878\,
            DIN => \N__8877\,
            DOUT => \N__8876\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8878\,
            PADOUT => \N__8877\,
            PADIN => \N__8876\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TCIn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8869\,
            DIN => \N__8868\,
            DOUT => \N__8867\,
            PACKAGEPIN => \A_040_wire\(0)
        );

    \A_040_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8869\,
            PADOUT => \N__8868\,
            PADIN => \N__8867\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8860\,
            DIN => \N__8859\,
            DOUT => \N__8858\,
            PACKAGEPIN => D_LM_AMIGA(0)
        );

    \D_LM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8860\,
            PADOUT => \N__8859\,
            PADIN => \N__8858\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5396\,
            DIN0 => \D_LM_AMIGA_in_0\,
            DOUT0 => \N__3258\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8851\,
            DIN => \N__8850\,
            DOUT => \N__8849\,
            PACKAGEPIN => \TBI_CPUn_wire\
        );

    \TBI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8851\,
            PADOUT => \N__8850\,
            PADIN => \N__8849\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6588\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8842\,
            DIN => \N__8841\,
            DOUT => \N__8840\,
            PACKAGEPIN => \CLK40A_wire\
        );

    \CLK40A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8842\,
            PADOUT => \N__8841\,
            PADIN => \N__8840\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3563\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8833\,
            DIN => \N__8832\,
            DOUT => \N__8831\,
            PACKAGEPIN => D_LM_040(3)
        );

    \D_LM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8833\,
            PADOUT => \N__8832\,
            PADIN => \N__8831\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7654\,
            DIN0 => \D_LM_040_in_3\,
            DOUT0 => \N__3411\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8824\,
            DIN => \N__8823\,
            DOUT => \N__8822\,
            PACKAGEPIN => D_LM_AMIGA(5)
        );

    \D_LM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8824\,
            PADOUT => \N__8823\,
            PADIN => \N__8822\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5370\,
            DIN0 => \D_LM_AMIGA_in_5\,
            DOUT0 => \N__8361\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8815\,
            DIN => \N__8814\,
            DOUT => \N__8813\,
            PACKAGEPIN => D_LM_040(6)
        );

    \D_LM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8815\,
            PADOUT => \N__8814\,
            PADIN => \N__8813\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7547\,
            DIN0 => \D_LM_040_in_6\,
            DOUT0 => \N__3999\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8806\,
            DIN => \N__8805\,
            DOUT => \N__8804\,
            PACKAGEPIN => D_UM_040(5)
        );

    \D_UM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8806\,
            PADOUT => \N__8805\,
            PADIN => \N__8804\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7655\,
            DIN0 => \D_UM_040_in_5\,
            DOUT0 => \N__7902\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8797\,
            DIN => \N__8796\,
            DOUT => \N__8795\,
            PACKAGEPIN => D_LL_AMIGA(3)
        );

    \D_LL_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8797\,
            PADOUT => \N__8796\,
            PADIN => \N__8795\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5284\,
            DIN0 => \D_LL_AMIGA_in_3\,
            DOUT0 => \N__3965\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8788\,
            DIN => \N__8787\,
            DOUT => \N__8786\,
            PACKAGEPIN => D_UU_AMIGA(3)
        );

    \D_UU_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8788\,
            PADOUT => \N__8787\,
            PADIN => \N__8786\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5461\,
            DIN0 => \D_UU_AMIGA_in_3\,
            DOUT0 => \N__4344\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8779\,
            DIN => \N__8778\,
            DOUT => \N__8777\,
            PACKAGEPIN => D_LL_040(5)
        );

    \D_LL_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8779\,
            PADOUT => \N__8778\,
            PADIN => \N__8777\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7629\,
            DIN0 => \D_LL_040_in_5\,
            DOUT0 => \N__2733\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8770\,
            DIN => \N__8769\,
            DOUT => \N__8768\,
            PACKAGEPIN => D_LL_AMIGA(6)
        );

    \D_LL_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8770\,
            PADOUT => \N__8769\,
            PADIN => \N__8768\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5397\,
            DIN0 => \D_LL_AMIGA_in_6\,
            DOUT0 => \N__3339\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8761\,
            DIN => \N__8760\,
            DOUT => \N__8759\,
            PACKAGEPIN => D_UU_AMIGA(6)
        );

    \D_UU_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8761\,
            PADOUT => \N__8760\,
            PADIN => \N__8759\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5468\,
            DIN0 => \D_UU_AMIGA_in_6\,
            DOUT0 => \N__3132\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8752\,
            DIN => \N__8751\,
            DOUT => \N__8750\,
            PACKAGEPIN => D_UM_AMIGA(1)
        );

    \D_UM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8752\,
            PADOUT => \N__8751\,
            PADIN => \N__8750\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5371\,
            DIN0 => \D_UM_AMIGA_in_1\,
            DOUT0 => \N__6054\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8743\,
            DIN => \N__8742\,
            DOUT => \N__8741\,
            PACKAGEPIN => D_UU_040(5)
        );

    \D_UU_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8743\,
            PADOUT => \N__8742\,
            PADIN => \N__8741\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7656\,
            DIN0 => \D_UU_040_in_5\,
            DOUT0 => \N__4926\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8734\,
            DIN => \N__8733\,
            DOUT => \N__8732\,
            PACKAGEPIN => \CLKRAMA_wire\
        );

    \CLKRAMA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8734\,
            PADOUT => \N__8733\,
            PADIN => \N__8732\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3564\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8725\,
            DIN => \N__8724\,
            DOUT => \N__8723\,
            PACKAGEPIN => D_LL_040(2)
        );

    \D_LL_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8725\,
            PADOUT => \N__8724\,
            PADIN => \N__8723\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7631\,
            DIN0 => \D_LL_040_in_2\,
            DOUT0 => \N__3768\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8716\,
            DIN => \N__8715\,
            DOUT => \N__8714\,
            PACKAGEPIN => \TCI_CPUn_wire\
        );

    \TCI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8716\,
            PADOUT => \N__8715\,
            PADIN => \N__8714\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6789\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BBn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8707\,
            DIN => \N__8706\,
            DOUT => \N__8705\,
            PACKAGEPIN => \BBn_wire\
        );

    \BBn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8707\,
            PADOUT => \N__8706\,
            PADIN => \N__8705\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BBn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMAAn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8698\,
            DIN => \N__8697\,
            DOUT => \N__8696\,
            PACKAGEPIN => \DMAAn_wire\
        );

    \DMAAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8698\,
            PADOUT => \N__8697\,
            PADIN => \N__8696\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3642\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8689\,
            DIN => \N__8688\,
            DOUT => \N__8687\,
            PACKAGEPIN => D_UM_AMIGA(4)
        );

    \D_UM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8689\,
            PADOUT => \N__8688\,
            PADIN => \N__8687\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5433\,
            DIN0 => \D_UM_AMIGA_in_4\,
            DOUT0 => \N__2823\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8680\,
            DIN => \N__8679\,
            DOUT => \N__8678\,
            PACKAGEPIN => D_LM_AMIGA(6)
        );

    \D_LM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8680\,
            PADOUT => \N__8679\,
            PADIN => \N__8678\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5373\,
            DIN0 => \D_LM_AMIGA_in_6\,
            DOUT0 => \N__3171\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8671\,
            DIN => \N__8670\,
            DOUT => \N__8669\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8671\,
            PADOUT => \N__8670\,
            PADIN => \N__8669\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8662\,
            DIN => \N__8661\,
            DOUT => \N__8660\,
            PACKAGEPIN => D_LM_040(5)
        );

    \D_LM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8662\,
            PADOUT => \N__8661\,
            PADIN => \N__8660\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7560\,
            DIN0 => \D_LM_040_in_5\,
            DOUT0 => \N__3438\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8653\,
            DIN => \N__8652\,
            DOUT => \N__8651\,
            PACKAGEPIN => D_UM_040(6)
        );

    \D_UM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8653\,
            PADOUT => \N__8652\,
            PADIN => \N__8651\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7546\,
            DIN0 => \D_UM_040_in_6\,
            DOUT0 => \N__8634\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2218\ : IoInMux
    port map (
            O => \N__8634\,
            I => \N__8631\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__8631\,
            I => \N__8628\
        );

    \I__2216\ : Span4Mux_s2_h
    port map (
            O => \N__8628\,
            I => \N__8625\
        );

    \I__2215\ : Sp12to4
    port map (
            O => \N__8625\,
            I => \N__8622\
        );

    \I__2214\ : Span12Mux_v
    port map (
            O => \N__8622\,
            I => \N__8619\
        );

    \I__2213\ : Odrv12
    port map (
            O => \N__8619\,
            I => \un1_D_UM_AMIGA_6\
        );

    \I__2212\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8612\
        );

    \I__2211\ : InMux
    port map (
            O => \N__8615\,
            I => \N__8609\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__8612\,
            I => \N__8605\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__8609\,
            I => \N__8602\
        );

    \I__2208\ : InMux
    port map (
            O => \N__8608\,
            I => \N__8599\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__8605\,
            I => \N__8596\
        );

    \I__2206\ : Span4Mux_v
    port map (
            O => \N__8602\,
            I => \N__8591\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__8599\,
            I => \N__8591\
        );

    \I__2204\ : Sp12to4
    port map (
            O => \N__8596\,
            I => \N__8588\
        );

    \I__2203\ : Span4Mux_v
    port map (
            O => \N__8591\,
            I => \N__8585\
        );

    \I__2202\ : Span12Mux_h
    port map (
            O => \N__8588\,
            I => \N__8582\
        );

    \I__2201\ : Span4Mux_v
    port map (
            O => \N__8585\,
            I => \N__8579\
        );

    \I__2200\ : Span12Mux_v
    port map (
            O => \N__8582\,
            I => \N__8576\
        );

    \I__2199\ : Sp12to4
    port map (
            O => \N__8579\,
            I => \N__8573\
        );

    \I__2198\ : Span12Mux_v
    port map (
            O => \N__8576\,
            I => \N__8568\
        );

    \I__2197\ : Span12Mux_h
    port map (
            O => \N__8573\,
            I => \N__8568\
        );

    \I__2196\ : Odrv12
    port map (
            O => \N__8568\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__2195\ : InMux
    port map (
            O => \N__8565\,
            I => \N__8562\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__8559\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\
        );

    \I__2192\ : IoInMux
    port map (
            O => \N__8556\,
            I => \N__8553\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__8553\,
            I => \N__8550\
        );

    \I__2190\ : IoSpan4Mux
    port map (
            O => \N__8550\,
            I => \N__8547\
        );

    \I__2189\ : Span4Mux_s0_h
    port map (
            O => \N__8547\,
            I => \N__8544\
        );

    \I__2188\ : Sp12to4
    port map (
            O => \N__8544\,
            I => \N__8541\
        );

    \I__2187\ : Span12Mux_h
    port map (
            O => \N__8541\,
            I => \N__8538\
        );

    \I__2186\ : Odrv12
    port map (
            O => \N__8538\,
            I => \un1_D_UM_AMIGA_3\
        );

    \I__2185\ : IoInMux
    port map (
            O => \N__8535\,
            I => \N__8532\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__8532\,
            I => \N__8528\
        );

    \I__2183\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8525\
        );

    \I__2182\ : IoSpan4Mux
    port map (
            O => \N__8528\,
            I => \N__8522\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__8525\,
            I => \N__8519\
        );

    \I__2180\ : Span4Mux_s3_h
    port map (
            O => \N__8522\,
            I => \N__8516\
        );

    \I__2179\ : Span4Mux_h
    port map (
            O => \N__8519\,
            I => \N__8513\
        );

    \I__2178\ : Sp12to4
    port map (
            O => \N__8516\,
            I => \N__8510\
        );

    \I__2177\ : Sp12to4
    port map (
            O => \N__8513\,
            I => \N__8507\
        );

    \I__2176\ : Span12Mux_v
    port map (
            O => \N__8510\,
            I => \N__8504\
        );

    \I__2175\ : Span12Mux_v
    port map (
            O => \N__8507\,
            I => \N__8501\
        );

    \I__2174\ : Span12Mux_h
    port map (
            O => \N__8504\,
            I => \N__8498\
        );

    \I__2173\ : Span12Mux_v
    port map (
            O => \N__8501\,
            I => \N__8495\
        );

    \I__2172\ : Span12Mux_h
    port map (
            O => \N__8498\,
            I => \N__8492\
        );

    \I__2171\ : Span12Mux_h
    port map (
            O => \N__8495\,
            I => \N__8489\
        );

    \I__2170\ : Odrv12
    port map (
            O => \N__8492\,
            I => \D_LL_040_in_7\
        );

    \I__2169\ : Odrv12
    port map (
            O => \N__8489\,
            I => \D_LL_040_in_7\
        );

    \I__2168\ : InMux
    port map (
            O => \N__8484\,
            I => \N__8481\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__8481\,
            I => \N__8478\
        );

    \I__2166\ : Span4Mux_v
    port map (
            O => \N__8478\,
            I => \N__8475\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__8475\,
            I => \N__8472\
        );

    \I__2164\ : Sp12to4
    port map (
            O => \N__8472\,
            I => \N__8469\
        );

    \I__2163\ : Span12Mux_h
    port map (
            O => \N__8469\,
            I => \N__8466\
        );

    \I__2162\ : Odrv12
    port map (
            O => \N__8466\,
            I => \D_UM_040_in_7\
        );

    \I__2161\ : IoInMux
    port map (
            O => \N__8463\,
            I => \N__8460\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__8460\,
            I => \N__8457\
        );

    \I__2159\ : IoSpan4Mux
    port map (
            O => \N__8457\,
            I => \N__8454\
        );

    \I__2158\ : Span4Mux_s0_h
    port map (
            O => \N__8454\,
            I => \N__8451\
        );

    \I__2157\ : Sp12to4
    port map (
            O => \N__8451\,
            I => \N__8448\
        );

    \I__2156\ : Span12Mux_s11_h
    port map (
            O => \N__8448\,
            I => \N__8445\
        );

    \I__2155\ : Odrv12
    port map (
            O => \N__8445\,
            I => \un1_D_UM_040_7\
        );

    \I__2154\ : InMux
    port map (
            O => \N__8442\,
            I => \N__8439\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__8439\,
            I => \N__8436\
        );

    \I__2152\ : Span12Mux_s9_v
    port map (
            O => \N__8436\,
            I => \N__8433\
        );

    \I__2151\ : Odrv12
    port map (
            O => \N__8433\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\
        );

    \I__2150\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8427\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__8427\,
            I => \N__8423\
        );

    \I__2148\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8419\
        );

    \I__2147\ : Span4Mux_v
    port map (
            O => \N__8423\,
            I => \N__8416\
        );

    \I__2146\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8413\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__8419\,
            I => \N__8410\
        );

    \I__2144\ : Span4Mux_v
    port map (
            O => \N__8416\,
            I => \N__8405\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__8413\,
            I => \N__8405\
        );

    \I__2142\ : Span4Mux_v
    port map (
            O => \N__8410\,
            I => \N__8402\
        );

    \I__2141\ : Span4Mux_v
    port map (
            O => \N__8405\,
            I => \N__8399\
        );

    \I__2140\ : Sp12to4
    port map (
            O => \N__8402\,
            I => \N__8396\
        );

    \I__2139\ : Sp12to4
    port map (
            O => \N__8399\,
            I => \N__8393\
        );

    \I__2138\ : Span12Mux_v
    port map (
            O => \N__8396\,
            I => \N__8390\
        );

    \I__2137\ : Span12Mux_h
    port map (
            O => \N__8393\,
            I => \N__8387\
        );

    \I__2136\ : Odrv12
    port map (
            O => \N__8390\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__2135\ : Odrv12
    port map (
            O => \N__8387\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__2134\ : IoInMux
    port map (
            O => \N__8382\,
            I => \N__8379\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__8379\,
            I => \N__8376\
        );

    \I__2132\ : IoSpan4Mux
    port map (
            O => \N__8376\,
            I => \N__8373\
        );

    \I__2131\ : IoSpan4Mux
    port map (
            O => \N__8373\,
            I => \N__8370\
        );

    \I__2130\ : Span4Mux_s3_h
    port map (
            O => \N__8370\,
            I => \N__8367\
        );

    \I__2129\ : Sp12to4
    port map (
            O => \N__8367\,
            I => \N__8364\
        );

    \I__2128\ : Odrv12
    port map (
            O => \N__8364\,
            I => \un1_D_UM_AMIGA_7\
        );

    \I__2127\ : IoInMux
    port map (
            O => \N__8361\,
            I => \N__8358\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__8358\,
            I => \N__8355\
        );

    \I__2125\ : IoSpan4Mux
    port map (
            O => \N__8355\,
            I => \N__8352\
        );

    \I__2124\ : IoSpan4Mux
    port map (
            O => \N__8352\,
            I => \N__8349\
        );

    \I__2123\ : Span4Mux_s2_h
    port map (
            O => \N__8349\,
            I => \N__8345\
        );

    \I__2122\ : InMux
    port map (
            O => \N__8348\,
            I => \N__8342\
        );

    \I__2121\ : Sp12to4
    port map (
            O => \N__8345\,
            I => \N__8339\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__8342\,
            I => \N__8336\
        );

    \I__2119\ : Span12Mux_h
    port map (
            O => \N__8339\,
            I => \N__8333\
        );

    \I__2118\ : Span12Mux_v
    port map (
            O => \N__8336\,
            I => \N__8330\
        );

    \I__2117\ : Span12Mux_h
    port map (
            O => \N__8333\,
            I => \N__8327\
        );

    \I__2116\ : Span12Mux_h
    port map (
            O => \N__8330\,
            I => \N__8324\
        );

    \I__2115\ : Odrv12
    port map (
            O => \N__8327\,
            I => \D_LM_040_in_5\
        );

    \I__2114\ : Odrv12
    port map (
            O => \N__8324\,
            I => \D_LM_040_in_5\
        );

    \I__2113\ : InMux
    port map (
            O => \N__8319\,
            I => \N__8316\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__8316\,
            I => \N__8313\
        );

    \I__2111\ : Span12Mux_v
    port map (
            O => \N__8313\,
            I => \N__8310\
        );

    \I__2110\ : Span12Mux_h
    port map (
            O => \N__8310\,
            I => \N__8307\
        );

    \I__2109\ : Odrv12
    port map (
            O => \N__8307\,
            I => \D_UU_040_in_5\
        );

    \I__2108\ : IoInMux
    port map (
            O => \N__8304\,
            I => \N__8301\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__8301\,
            I => \N__8298\
        );

    \I__2106\ : Span4Mux_s2_h
    port map (
            O => \N__8298\,
            I => \N__8295\
        );

    \I__2105\ : Span4Mux_v
    port map (
            O => \N__8295\,
            I => \N__8292\
        );

    \I__2104\ : Sp12to4
    port map (
            O => \N__8292\,
            I => \N__8289\
        );

    \I__2103\ : Span12Mux_s10_h
    port map (
            O => \N__8289\,
            I => \N__8286\
        );

    \I__2102\ : Odrv12
    port map (
            O => \N__8286\,
            I => \un1_D_UU_040_5\
        );

    \I__2101\ : InMux
    port map (
            O => \N__8283\,
            I => \N__8280\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__8280\,
            I => \N__8277\
        );

    \I__2099\ : Span12Mux_s7_v
    port map (
            O => \N__8277\,
            I => \N__8274\
        );

    \I__2098\ : Span12Mux_h
    port map (
            O => \N__8274\,
            I => \N__8271\
        );

    \I__2097\ : Odrv12
    port map (
            O => \N__8271\,
            I => \D_UM_040_in_5\
        );

    \I__2096\ : IoInMux
    port map (
            O => \N__8268\,
            I => \N__8265\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__8265\,
            I => \N__8261\
        );

    \I__2094\ : InMux
    port map (
            O => \N__8264\,
            I => \N__8258\
        );

    \I__2093\ : IoSpan4Mux
    port map (
            O => \N__8261\,
            I => \N__8255\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__8258\,
            I => \N__8252\
        );

    \I__2091\ : Span4Mux_s3_h
    port map (
            O => \N__8255\,
            I => \N__8249\
        );

    \I__2090\ : Span4Mux_h
    port map (
            O => \N__8252\,
            I => \N__8246\
        );

    \I__2089\ : Sp12to4
    port map (
            O => \N__8249\,
            I => \N__8243\
        );

    \I__2088\ : Sp12to4
    port map (
            O => \N__8246\,
            I => \N__8240\
        );

    \I__2087\ : Span12Mux_v
    port map (
            O => \N__8243\,
            I => \N__8237\
        );

    \I__2086\ : Span12Mux_v
    port map (
            O => \N__8240\,
            I => \N__8234\
        );

    \I__2085\ : Span12Mux_h
    port map (
            O => \N__8237\,
            I => \N__8231\
        );

    \I__2084\ : Span12Mux_v
    port map (
            O => \N__8234\,
            I => \N__8228\
        );

    \I__2083\ : Span12Mux_h
    port map (
            O => \N__8231\,
            I => \N__8225\
        );

    \I__2082\ : Span12Mux_h
    port map (
            O => \N__8228\,
            I => \N__8222\
        );

    \I__2081\ : Odrv12
    port map (
            O => \N__8225\,
            I => \D_LL_040_in_5\
        );

    \I__2080\ : Odrv12
    port map (
            O => \N__8222\,
            I => \D_LL_040_in_5\
        );

    \I__2079\ : InMux
    port map (
            O => \N__8217\,
            I => \N__8201\
        );

    \I__2078\ : InMux
    port map (
            O => \N__8216\,
            I => \N__8201\
        );

    \I__2077\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8198\
        );

    \I__2076\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8192\
        );

    \I__2075\ : InMux
    port map (
            O => \N__8213\,
            I => \N__8192\
        );

    \I__2074\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8187\
        );

    \I__2073\ : InMux
    port map (
            O => \N__8211\,
            I => \N__8187\
        );

    \I__2072\ : InMux
    port map (
            O => \N__8210\,
            I => \N__8183\
        );

    \I__2071\ : InMux
    port map (
            O => \N__8209\,
            I => \N__8178\
        );

    \I__2070\ : InMux
    port map (
            O => \N__8208\,
            I => \N__8178\
        );

    \I__2069\ : InMux
    port map (
            O => \N__8207\,
            I => \N__8175\
        );

    \I__2068\ : InMux
    port map (
            O => \N__8206\,
            I => \N__8169\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__8201\,
            I => \N__8162\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__8198\,
            I => \N__8162\
        );

    \I__2065\ : InMux
    port map (
            O => \N__8197\,
            I => \N__8159\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__8192\,
            I => \N__8156\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__8187\,
            I => \N__8153\
        );

    \I__2062\ : InMux
    port map (
            O => \N__8186\,
            I => \N__8150\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__8183\,
            I => \N__8143\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__8178\,
            I => \N__8143\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__8175\,
            I => \N__8140\
        );

    \I__2058\ : InMux
    port map (
            O => \N__8174\,
            I => \N__8131\
        );

    \I__2057\ : InMux
    port map (
            O => \N__8173\,
            I => \N__8126\
        );

    \I__2056\ : InMux
    port map (
            O => \N__8172\,
            I => \N__8123\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__8169\,
            I => \N__8120\
        );

    \I__2054\ : InMux
    port map (
            O => \N__8168\,
            I => \N__8115\
        );

    \I__2053\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8115\
        );

    \I__2052\ : Span4Mux_v
    port map (
            O => \N__8162\,
            I => \N__8110\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__8159\,
            I => \N__8110\
        );

    \I__2050\ : Span4Mux_h
    port map (
            O => \N__8156\,
            I => \N__8103\
        );

    \I__2049\ : Span4Mux_h
    port map (
            O => \N__8153\,
            I => \N__8103\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__8150\,
            I => \N__8103\
        );

    \I__2047\ : InMux
    port map (
            O => \N__8149\,
            I => \N__8098\
        );

    \I__2046\ : InMux
    port map (
            O => \N__8148\,
            I => \N__8098\
        );

    \I__2045\ : Span4Mux_v
    port map (
            O => \N__8143\,
            I => \N__8093\
        );

    \I__2044\ : Span4Mux_v
    port map (
            O => \N__8140\,
            I => \N__8093\
        );

    \I__2043\ : InMux
    port map (
            O => \N__8139\,
            I => \N__8090\
        );

    \I__2042\ : InMux
    port map (
            O => \N__8138\,
            I => \N__8085\
        );

    \I__2041\ : InMux
    port map (
            O => \N__8137\,
            I => \N__8085\
        );

    \I__2040\ : InMux
    port map (
            O => \N__8136\,
            I => \N__8080\
        );

    \I__2039\ : InMux
    port map (
            O => \N__8135\,
            I => \N__8080\
        );

    \I__2038\ : InMux
    port map (
            O => \N__8134\,
            I => \N__8077\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__8131\,
            I => \N__8074\
        );

    \I__2036\ : InMux
    port map (
            O => \N__8130\,
            I => \N__8071\
        );

    \I__2035\ : InMux
    port map (
            O => \N__8129\,
            I => \N__8068\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__8126\,
            I => \N__8062\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__8123\,
            I => \N__8062\
        );

    \I__2032\ : Span4Mux_h
    port map (
            O => \N__8120\,
            I => \N__8057\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__8115\,
            I => \N__8057\
        );

    \I__2030\ : Span4Mux_v
    port map (
            O => \N__8110\,
            I => \N__8054\
        );

    \I__2029\ : Span4Mux_v
    port map (
            O => \N__8103\,
            I => \N__8049\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__8098\,
            I => \N__8049\
        );

    \I__2027\ : Span4Mux_v
    port map (
            O => \N__8093\,
            I => \N__8044\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__8090\,
            I => \N__8044\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__8085\,
            I => \N__8037\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__8080\,
            I => \N__8037\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__8077\,
            I => \N__8037\
        );

    \I__2022\ : Span4Mux_v
    port map (
            O => \N__8074\,
            I => \N__8030\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__8071\,
            I => \N__8030\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__8068\,
            I => \N__8030\
        );

    \I__2019\ : InMux
    port map (
            O => \N__8067\,
            I => \N__8027\
        );

    \I__2018\ : Span12Mux_v
    port map (
            O => \N__8062\,
            I => \N__8021\
        );

    \I__2017\ : Span4Mux_v
    port map (
            O => \N__8057\,
            I => \N__8018\
        );

    \I__2016\ : Span4Mux_h
    port map (
            O => \N__8054\,
            I => \N__8013\
        );

    \I__2015\ : Span4Mux_v
    port map (
            O => \N__8049\,
            I => \N__8013\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__8044\,
            I => \N__8006\
        );

    \I__2013\ : Span4Mux_v
    port map (
            O => \N__8037\,
            I => \N__8006\
        );

    \I__2012\ : Span4Mux_v
    port map (
            O => \N__8030\,
            I => \N__8006\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__8027\,
            I => \N__8003\
        );

    \I__2010\ : InMux
    port map (
            O => \N__8026\,
            I => \N__7998\
        );

    \I__2009\ : InMux
    port map (
            O => \N__8025\,
            I => \N__7998\
        );

    \I__2008\ : InMux
    port map (
            O => \N__8024\,
            I => \N__7995\
        );

    \I__2007\ : Odrv12
    port map (
            O => \N__8021\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__2006\ : Odrv4
    port map (
            O => \N__8018\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__8013\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__8006\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__8003\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__7998\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__7995\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__2000\ : IoInMux
    port map (
            O => \N__7980\,
            I => \N__7977\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__7977\,
            I => \N__7974\
        );

    \I__1998\ : Span12Mux_s6_v
    port map (
            O => \N__7974\,
            I => \N__7971\
        );

    \I__1997\ : Span12Mux_h
    port map (
            O => \N__7971\,
            I => \N__7968\
        );

    \I__1996\ : Odrv12
    port map (
            O => \N__7968\,
            I => \un1_D_UM_040_5\
        );

    \I__1995\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7962\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__7962\,
            I => \N__7959\
        );

    \I__1993\ : Sp12to4
    port map (
            O => \N__7959\,
            I => \N__7956\
        );

    \I__1992\ : Odrv12
    port map (
            O => \N__7956\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\
        );

    \I__1991\ : InMux
    port map (
            O => \N__7953\,
            I => \N__7949\
        );

    \I__1990\ : InMux
    port map (
            O => \N__7952\,
            I => \N__7946\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__7949\,
            I => \N__7943\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__7946\,
            I => \N__7939\
        );

    \I__1987\ : Span4Mux_v
    port map (
            O => \N__7943\,
            I => \N__7936\
        );

    \I__1986\ : InMux
    port map (
            O => \N__7942\,
            I => \N__7933\
        );

    \I__1985\ : Span4Mux_v
    port map (
            O => \N__7939\,
            I => \N__7930\
        );

    \I__1984\ : Span4Mux_v
    port map (
            O => \N__7936\,
            I => \N__7925\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__7933\,
            I => \N__7925\
        );

    \I__1982\ : Sp12to4
    port map (
            O => \N__7930\,
            I => \N__7922\
        );

    \I__1981\ : Span4Mux_v
    port map (
            O => \N__7925\,
            I => \N__7919\
        );

    \I__1980\ : Span12Mux_h
    port map (
            O => \N__7922\,
            I => \N__7916\
        );

    \I__1979\ : Sp12to4
    port map (
            O => \N__7919\,
            I => \N__7913\
        );

    \I__1978\ : Span12Mux_v
    port map (
            O => \N__7916\,
            I => \N__7910\
        );

    \I__1977\ : Span12Mux_h
    port map (
            O => \N__7913\,
            I => \N__7907\
        );

    \I__1976\ : Odrv12
    port map (
            O => \N__7910\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1975\ : Odrv12
    port map (
            O => \N__7907\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1974\ : IoInMux
    port map (
            O => \N__7902\,
            I => \N__7899\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__7899\,
            I => \N__7896\
        );

    \I__1972\ : Span12Mux_s11_v
    port map (
            O => \N__7896\,
            I => \N__7893\
        );

    \I__1971\ : Span12Mux_h
    port map (
            O => \N__7893\,
            I => \N__7890\
        );

    \I__1970\ : Odrv12
    port map (
            O => \N__7890\,
            I => \un1_D_UM_AMIGA_5\
        );

    \I__1969\ : InMux
    port map (
            O => \N__7887\,
            I => \N__7884\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__7884\,
            I => \N__7877\
        );

    \I__1967\ : InMux
    port map (
            O => \N__7883\,
            I => \N__7867\
        );

    \I__1966\ : InMux
    port map (
            O => \N__7882\,
            I => \N__7867\
        );

    \I__1965\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7867\
        );

    \I__1964\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7867\
        );

    \I__1963\ : Span4Mux_v
    port map (
            O => \N__7877\,
            I => \N__7858\
        );

    \I__1962\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7855\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__7867\,
            I => \N__7852\
        );

    \I__1960\ : InMux
    port map (
            O => \N__7866\,
            I => \N__7845\
        );

    \I__1959\ : InMux
    port map (
            O => \N__7865\,
            I => \N__7845\
        );

    \I__1958\ : InMux
    port map (
            O => \N__7864\,
            I => \N__7845\
        );

    \I__1957\ : InMux
    port map (
            O => \N__7863\,
            I => \N__7842\
        );

    \I__1956\ : InMux
    port map (
            O => \N__7862\,
            I => \N__7837\
        );

    \I__1955\ : InMux
    port map (
            O => \N__7861\,
            I => \N__7837\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__7858\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__7855\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__7852\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__7845\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__7842\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__7837\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1948\ : IoInMux
    port map (
            O => \N__7824\,
            I => \N__7821\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__7821\,
            I => \N__7817\
        );

    \I__1946\ : IoInMux
    port map (
            O => \N__7820\,
            I => \N__7814\
        );

    \I__1945\ : Span4Mux_s0_h
    port map (
            O => \N__7817\,
            I => \N__7811\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__7814\,
            I => \N__7808\
        );

    \I__1943\ : Span4Mux_h
    port map (
            O => \N__7811\,
            I => \N__7802\
        );

    \I__1942\ : IoSpan4Mux
    port map (
            O => \N__7808\,
            I => \N__7799\
        );

    \I__1941\ : InMux
    port map (
            O => \N__7807\,
            I => \N__7792\
        );

    \I__1940\ : InMux
    port map (
            O => \N__7806\,
            I => \N__7792\
        );

    \I__1939\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7792\
        );

    \I__1938\ : Span4Mux_h
    port map (
            O => \N__7802\,
            I => \N__7788\
        );

    \I__1937\ : Span4Mux_s2_v
    port map (
            O => \N__7799\,
            I => \N__7785\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__7792\,
            I => \N__7782\
        );

    \I__1935\ : InMux
    port map (
            O => \N__7791\,
            I => \N__7779\
        );

    \I__1934\ : Span4Mux_h
    port map (
            O => \N__7788\,
            I => \N__7776\
        );

    \I__1933\ : Span4Mux_v
    port map (
            O => \N__7785\,
            I => \N__7770\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__7782\,
            I => \N__7770\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__7779\,
            I => \N__7766\
        );

    \I__1930\ : Span4Mux_h
    port map (
            O => \N__7776\,
            I => \N__7763\
        );

    \I__1929\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7760\
        );

    \I__1928\ : Span4Mux_v
    port map (
            O => \N__7770\,
            I => \N__7757\
        );

    \I__1927\ : InMux
    port map (
            O => \N__7769\,
            I => \N__7754\
        );

    \I__1926\ : Span4Mux_h
    port map (
            O => \N__7766\,
            I => \N__7751\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__7763\,
            I => \N__7746\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__7760\,
            I => \N__7746\
        );

    \I__1923\ : Span4Mux_v
    port map (
            O => \N__7757\,
            I => \N__7741\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__7754\,
            I => \N__7741\
        );

    \I__1921\ : Sp12to4
    port map (
            O => \N__7751\,
            I => \N__7738\
        );

    \I__1920\ : Span4Mux_v
    port map (
            O => \N__7746\,
            I => \N__7735\
        );

    \I__1919\ : Span4Mux_h
    port map (
            O => \N__7741\,
            I => \N__7732\
        );

    \I__1918\ : Odrv12
    port map (
            O => \N__7738\,
            I => \CPUBGn_c\
        );

    \I__1917\ : Odrv4
    port map (
            O => \N__7735\,
            I => \CPUBGn_c\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__7732\,
            I => \CPUBGn_c\
        );

    \I__1915\ : InMux
    port map (
            O => \N__7725\,
            I => \N__7721\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__7724\,
            I => \N__7716\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__7721\,
            I => \N__7713\
        );

    \I__1912\ : CascadeMux
    port map (
            O => \N__7720\,
            I => \N__7710\
        );

    \I__1911\ : InMux
    port map (
            O => \N__7719\,
            I => \N__7705\
        );

    \I__1910\ : InMux
    port map (
            O => \N__7716\,
            I => \N__7705\
        );

    \I__1909\ : Span4Mux_v
    port map (
            O => \N__7713\,
            I => \N__7701\
        );

    \I__1908\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7698\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__7705\,
            I => \N__7695\
        );

    \I__1906\ : InMux
    port map (
            O => \N__7704\,
            I => \N__7692\
        );

    \I__1905\ : Span4Mux_h
    port map (
            O => \N__7701\,
            I => \N__7689\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__7698\,
            I => \N__7686\
        );

    \I__1903\ : Span4Mux_h
    port map (
            O => \N__7695\,
            I => \N__7681\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__7692\,
            I => \N__7681\
        );

    \I__1901\ : Span4Mux_v
    port map (
            O => \N__7689\,
            I => \N__7676\
        );

    \I__1900\ : Span4Mux_v
    port map (
            O => \N__7686\,
            I => \N__7676\
        );

    \I__1899\ : Span4Mux_v
    port map (
            O => \N__7681\,
            I => \N__7673\
        );

    \I__1898\ : Sp12to4
    port map (
            O => \N__7676\,
            I => \N__7670\
        );

    \I__1897\ : Sp12to4
    port map (
            O => \N__7673\,
            I => \N__7667\
        );

    \I__1896\ : Span12Mux_h
    port map (
            O => \N__7670\,
            I => \N__7664\
        );

    \I__1895\ : Span12Mux_h
    port map (
            O => \N__7667\,
            I => \N__7661\
        );

    \I__1894\ : Odrv12
    port map (
            O => \N__7664\,
            I => \RnW_c\
        );

    \I__1893\ : Odrv12
    port map (
            O => \N__7661\,
            I => \RnW_c\
        );

    \I__1892\ : IoInMux
    port map (
            O => \N__7656\,
            I => \N__7650\
        );

    \I__1891\ : IoInMux
    port map (
            O => \N__7655\,
            I => \N__7647\
        );

    \I__1890\ : IoInMux
    port map (
            O => \N__7654\,
            I => \N__7641\
        );

    \I__1889\ : IoInMux
    port map (
            O => \N__7653\,
            I => \N__7638\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__7650\,
            I => \N__7624\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__7647\,
            I => \N__7624\
        );

    \I__1886\ : IoInMux
    port map (
            O => \N__7646\,
            I => \N__7621\
        );

    \I__1885\ : IoInMux
    port map (
            O => \N__7645\,
            I => \N__7618\
        );

    \I__1884\ : IoInMux
    port map (
            O => \N__7644\,
            I => \N__7615\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__7641\,
            I => \N__7611\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__7638\,
            I => \N__7607\
        );

    \I__1881\ : IoInMux
    port map (
            O => \N__7637\,
            I => \N__7604\
        );

    \I__1880\ : IoInMux
    port map (
            O => \N__7636\,
            I => \N__7601\
        );

    \I__1879\ : IoInMux
    port map (
            O => \N__7635\,
            I => \N__7597\
        );

    \I__1878\ : IoInMux
    port map (
            O => \N__7634\,
            I => \N__7594\
        );

    \I__1877\ : IoInMux
    port map (
            O => \N__7633\,
            I => \N__7591\
        );

    \I__1876\ : IoInMux
    port map (
            O => \N__7632\,
            I => \N__7588\
        );

    \I__1875\ : IoInMux
    port map (
            O => \N__7631\,
            I => \N__7585\
        );

    \I__1874\ : IoInMux
    port map (
            O => \N__7630\,
            I => \N__7582\
        );

    \I__1873\ : IoInMux
    port map (
            O => \N__7629\,
            I => \N__7579\
        );

    \I__1872\ : IoSpan4Mux
    port map (
            O => \N__7624\,
            I => \N__7570\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__7621\,
            I => \N__7570\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__7618\,
            I => \N__7570\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__7615\,
            I => \N__7570\
        );

    \I__1868\ : IoInMux
    port map (
            O => \N__7614\,
            I => \N__7567\
        );

    \I__1867\ : Span4Mux_s2_h
    port map (
            O => \N__7611\,
            I => \N__7564\
        );

    \I__1866\ : IoInMux
    port map (
            O => \N__7610\,
            I => \N__7561\
        );

    \I__1865\ : IoSpan4Mux
    port map (
            O => \N__7607\,
            I => \N__7551\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__7604\,
            I => \N__7551\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__7601\,
            I => \N__7551\
        );

    \I__1862\ : IoInMux
    port map (
            O => \N__7600\,
            I => \N__7548\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__7597\,
            I => \N__7541\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__7594\,
            I => \N__7541\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__7591\,
            I => \N__7530\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__7588\,
            I => \N__7530\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__7585\,
            I => \N__7530\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__7582\,
            I => \N__7530\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__7579\,
            I => \N__7530\
        );

    \I__1854\ : IoSpan4Mux
    port map (
            O => \N__7570\,
            I => \N__7524\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__7567\,
            I => \N__7521\
        );

    \I__1852\ : Span4Mux_v
    port map (
            O => \N__7564\,
            I => \N__7516\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__7561\,
            I => \N__7516\
        );

    \I__1850\ : IoInMux
    port map (
            O => \N__7560\,
            I => \N__7513\
        );

    \I__1849\ : IoInMux
    port map (
            O => \N__7559\,
            I => \N__7510\
        );

    \I__1848\ : IoInMux
    port map (
            O => \N__7558\,
            I => \N__7507\
        );

    \I__1847\ : IoSpan4Mux
    port map (
            O => \N__7551\,
            I => \N__7502\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__7548\,
            I => \N__7502\
        );

    \I__1845\ : IoInMux
    port map (
            O => \N__7547\,
            I => \N__7499\
        );

    \I__1844\ : IoInMux
    port map (
            O => \N__7546\,
            I => \N__7496\
        );

    \I__1843\ : Span4Mux_s3_h
    port map (
            O => \N__7541\,
            I => \N__7491\
        );

    \I__1842\ : IoSpan4Mux
    port map (
            O => \N__7530\,
            I => \N__7488\
        );

    \I__1841\ : IoInMux
    port map (
            O => \N__7529\,
            I => \N__7485\
        );

    \I__1840\ : IoInMux
    port map (
            O => \N__7528\,
            I => \N__7482\
        );

    \I__1839\ : IoInMux
    port map (
            O => \N__7527\,
            I => \N__7476\
        );

    \I__1838\ : Span4Mux_s2_v
    port map (
            O => \N__7524\,
            I => \N__7473\
        );

    \I__1837\ : Span4Mux_s2_v
    port map (
            O => \N__7521\,
            I => \N__7470\
        );

    \I__1836\ : IoSpan4Mux
    port map (
            O => \N__7516\,
            I => \N__7461\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__7513\,
            I => \N__7461\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__7510\,
            I => \N__7461\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__7507\,
            I => \N__7461\
        );

    \I__1832\ : IoSpan4Mux
    port map (
            O => \N__7502\,
            I => \N__7454\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__7499\,
            I => \N__7454\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__7496\,
            I => \N__7454\
        );

    \I__1829\ : IoInMux
    port map (
            O => \N__7495\,
            I => \N__7451\
        );

    \I__1828\ : IoInMux
    port map (
            O => \N__7494\,
            I => \N__7448\
        );

    \I__1827\ : Span4Mux_v
    port map (
            O => \N__7491\,
            I => \N__7443\
        );

    \I__1826\ : Span4Mux_s3_h
    port map (
            O => \N__7488\,
            I => \N__7443\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__7485\,
            I => \N__7440\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__7482\,
            I => \N__7437\
        );

    \I__1823\ : IoInMux
    port map (
            O => \N__7481\,
            I => \N__7434\
        );

    \I__1822\ : IoInMux
    port map (
            O => \N__7480\,
            I => \N__7431\
        );

    \I__1821\ : IoInMux
    port map (
            O => \N__7479\,
            I => \N__7428\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__7476\,
            I => \N__7425\
        );

    \I__1819\ : Span4Mux_v
    port map (
            O => \N__7473\,
            I => \N__7420\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__7470\,
            I => \N__7420\
        );

    \I__1817\ : IoSpan4Mux
    port map (
            O => \N__7461\,
            I => \N__7415\
        );

    \I__1816\ : IoSpan4Mux
    port map (
            O => \N__7454\,
            I => \N__7415\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__7451\,
            I => \N__7410\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__7448\,
            I => \N__7410\
        );

    \I__1813\ : Sp12to4
    port map (
            O => \N__7443\,
            I => \N__7403\
        );

    \I__1812\ : Sp12to4
    port map (
            O => \N__7440\,
            I => \N__7403\
        );

    \I__1811\ : Span12Mux_s1_h
    port map (
            O => \N__7437\,
            I => \N__7403\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__7434\,
            I => \N__7398\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__7431\,
            I => \N__7398\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__7428\,
            I => \N__7395\
        );

    \I__1807\ : Span4Mux_s3_v
    port map (
            O => \N__7425\,
            I => \N__7392\
        );

    \I__1806\ : Span4Mux_v
    port map (
            O => \N__7420\,
            I => \N__7389\
        );

    \I__1805\ : Span4Mux_s2_h
    port map (
            O => \N__7415\,
            I => \N__7386\
        );

    \I__1804\ : Span12Mux_s8_h
    port map (
            O => \N__7410\,
            I => \N__7383\
        );

    \I__1803\ : Span12Mux_h
    port map (
            O => \N__7403\,
            I => \N__7380\
        );

    \I__1802\ : Span12Mux_s3_v
    port map (
            O => \N__7398\,
            I => \N__7373\
        );

    \I__1801\ : Sp12to4
    port map (
            O => \N__7395\,
            I => \N__7373\
        );

    \I__1800\ : Sp12to4
    port map (
            O => \N__7392\,
            I => \N__7373\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__7389\,
            I => \N__7368\
        );

    \I__1798\ : Span4Mux_h
    port map (
            O => \N__7386\,
            I => \N__7368\
        );

    \I__1797\ : Span12Mux_v
    port map (
            O => \N__7383\,
            I => \N__7365\
        );

    \I__1796\ : Span12Mux_v
    port map (
            O => \N__7380\,
            I => \N__7360\
        );

    \I__1795\ : Span12Mux_h
    port map (
            O => \N__7373\,
            I => \N__7360\
        );

    \I__1794\ : Span4Mux_h
    port map (
            O => \N__7368\,
            I => \N__7357\
        );

    \I__1793\ : Odrv12
    port map (
            O => \N__7365\,
            I => \N_60_i\
        );

    \I__1792\ : Odrv12
    port map (
            O => \N__7360\,
            I => \N_60_i\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__7357\,
            I => \N_60_i\
        );

    \I__1790\ : InMux
    port map (
            O => \N__7350\,
            I => \N__7345\
        );

    \I__1789\ : InMux
    port map (
            O => \N__7349\,
            I => \N__7334\
        );

    \I__1788\ : InMux
    port map (
            O => \N__7348\,
            I => \N__7334\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__7345\,
            I => \N__7330\
        );

    \I__1786\ : InMux
    port map (
            O => \N__7344\,
            I => \N__7327\
        );

    \I__1785\ : InMux
    port map (
            O => \N__7343\,
            I => \N__7324\
        );

    \I__1784\ : InMux
    port map (
            O => \N__7342\,
            I => \N__7310\
        );

    \I__1783\ : InMux
    port map (
            O => \N__7341\,
            I => \N__7310\
        );

    \I__1782\ : InMux
    port map (
            O => \N__7340\,
            I => \N__7310\
        );

    \I__1781\ : InMux
    port map (
            O => \N__7339\,
            I => \N__7310\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__7334\,
            I => \N__7306\
        );

    \I__1779\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7303\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__7330\,
            I => \N__7298\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__7327\,
            I => \N__7298\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__7324\,
            I => \N__7295\
        );

    \I__1775\ : InMux
    port map (
            O => \N__7323\,
            I => \N__7292\
        );

    \I__1774\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7289\
        );

    \I__1773\ : InMux
    port map (
            O => \N__7321\,
            I => \N__7286\
        );

    \I__1772\ : InMux
    port map (
            O => \N__7320\,
            I => \N__7281\
        );

    \I__1771\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7281\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__7310\,
            I => \N__7277\
        );

    \I__1769\ : InMux
    port map (
            O => \N__7309\,
            I => \N__7274\
        );

    \I__1768\ : Span4Mux_v
    port map (
            O => \N__7306\,
            I => \N__7269\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__7303\,
            I => \N__7269\
        );

    \I__1766\ : Span4Mux_v
    port map (
            O => \N__7298\,
            I => \N__7258\
        );

    \I__1765\ : Span4Mux_h
    port map (
            O => \N__7295\,
            I => \N__7258\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__7292\,
            I => \N__7258\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__7289\,
            I => \N__7258\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__7286\,
            I => \N__7258\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__7281\,
            I => \N__7255\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__7280\,
            I => \N__7252\
        );

    \I__1759\ : Sp12to4
    port map (
            O => \N__7277\,
            I => \N__7247\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__7274\,
            I => \N__7247\
        );

    \I__1757\ : Span4Mux_v
    port map (
            O => \N__7269\,
            I => \N__7244\
        );

    \I__1756\ : Span4Mux_v
    port map (
            O => \N__7258\,
            I => \N__7239\
        );

    \I__1755\ : Span4Mux_v
    port map (
            O => \N__7255\,
            I => \N__7239\
        );

    \I__1754\ : InMux
    port map (
            O => \N__7252\,
            I => \N__7236\
        );

    \I__1753\ : Odrv12
    port map (
            O => \N__7247\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__7244\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1751\ : Odrv4
    port map (
            O => \N__7239\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__7236\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1749\ : InMux
    port map (
            O => \N__7227\,
            I => \N__7224\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__7224\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\
        );

    \I__1747\ : InMux
    port map (
            O => \N__7221\,
            I => \N__7218\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__7218\,
            I => \N__7215\
        );

    \I__1745\ : Span4Mux_v
    port map (
            O => \N__7215\,
            I => \N__7212\
        );

    \I__1744\ : Span4Mux_v
    port map (
            O => \N__7212\,
            I => \N__7207\
        );

    \I__1743\ : InMux
    port map (
            O => \N__7211\,
            I => \N__7204\
        );

    \I__1742\ : InMux
    port map (
            O => \N__7210\,
            I => \N__7201\
        );

    \I__1741\ : Sp12to4
    port map (
            O => \N__7207\,
            I => \N__7194\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__7204\,
            I => \N__7194\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__7201\,
            I => \N__7194\
        );

    \I__1738\ : Span12Mux_h
    port map (
            O => \N__7194\,
            I => \N__7191\
        );

    \I__1737\ : Span12Mux_v
    port map (
            O => \N__7191\,
            I => \N__7188\
        );

    \I__1736\ : Odrv12
    port map (
            O => \N__7188\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__1735\ : InMux
    port map (
            O => \N__7185\,
            I => \N__7182\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__7182\,
            I => \N__7179\
        );

    \I__1733\ : Span4Mux_v
    port map (
            O => \N__7179\,
            I => \N__7174\
        );

    \I__1732\ : InMux
    port map (
            O => \N__7178\,
            I => \N__7171\
        );

    \I__1731\ : InMux
    port map (
            O => \N__7177\,
            I => \N__7168\
        );

    \I__1730\ : Span4Mux_v
    port map (
            O => \N__7174\,
            I => \N__7161\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__7171\,
            I => \N__7161\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__7168\,
            I => \N__7161\
        );

    \I__1727\ : Span4Mux_v
    port map (
            O => \N__7161\,
            I => \N__7158\
        );

    \I__1726\ : Sp12to4
    port map (
            O => \N__7158\,
            I => \N__7155\
        );

    \I__1725\ : Span12Mux_h
    port map (
            O => \N__7155\,
            I => \N__7152\
        );

    \I__1724\ : Odrv12
    port map (
            O => \N__7152\,
            I => \D_UM_AMIGA_in_0\
        );

    \I__1723\ : InMux
    port map (
            O => \N__7149\,
            I => \N__7146\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__7146\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\
        );

    \I__1721\ : InMux
    port map (
            O => \N__7143\,
            I => \N__7140\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__7140\,
            I => \N__7137\
        );

    \I__1719\ : Glb2LocalMux
    port map (
            O => \N__7137\,
            I => \N__7089\
        );

    \I__1718\ : ClkMux
    port map (
            O => \N__7136\,
            I => \N__7089\
        );

    \I__1717\ : ClkMux
    port map (
            O => \N__7135\,
            I => \N__7089\
        );

    \I__1716\ : ClkMux
    port map (
            O => \N__7134\,
            I => \N__7089\
        );

    \I__1715\ : ClkMux
    port map (
            O => \N__7133\,
            I => \N__7089\
        );

    \I__1714\ : ClkMux
    port map (
            O => \N__7132\,
            I => \N__7089\
        );

    \I__1713\ : ClkMux
    port map (
            O => \N__7131\,
            I => \N__7089\
        );

    \I__1712\ : ClkMux
    port map (
            O => \N__7130\,
            I => \N__7089\
        );

    \I__1711\ : ClkMux
    port map (
            O => \N__7129\,
            I => \N__7089\
        );

    \I__1710\ : ClkMux
    port map (
            O => \N__7128\,
            I => \N__7089\
        );

    \I__1709\ : ClkMux
    port map (
            O => \N__7127\,
            I => \N__7089\
        );

    \I__1708\ : ClkMux
    port map (
            O => \N__7126\,
            I => \N__7089\
        );

    \I__1707\ : ClkMux
    port map (
            O => \N__7125\,
            I => \N__7089\
        );

    \I__1706\ : ClkMux
    port map (
            O => \N__7124\,
            I => \N__7089\
        );

    \I__1705\ : ClkMux
    port map (
            O => \N__7123\,
            I => \N__7089\
        );

    \I__1704\ : ClkMux
    port map (
            O => \N__7122\,
            I => \N__7089\
        );

    \I__1703\ : GlobalMux
    port map (
            O => \N__7089\,
            I => \CLK40\
        );

    \I__1702\ : CEMux
    port map (
            O => \N__7086\,
            I => \N__7082\
        );

    \I__1701\ : CEMux
    port map (
            O => \N__7085\,
            I => \N__7079\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__7082\,
            I => \N__7076\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__7079\,
            I => \N__7072\
        );

    \I__1698\ : Span4Mux_v
    port map (
            O => \N__7076\,
            I => \N__7069\
        );

    \I__1697\ : CEMux
    port map (
            O => \N__7075\,
            I => \N__7066\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__7072\,
            I => \N__7063\
        );

    \I__1695\ : Span4Mux_h
    port map (
            O => \N__7069\,
            I => \N__7060\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__7066\,
            I => \N__7057\
        );

    \I__1693\ : Span4Mux_h
    port map (
            O => \N__7063\,
            I => \N__7054\
        );

    \I__1692\ : Odrv4
    port map (
            O => \N__7060\,
            I => \U111_CYCLE_SM.N_99_i_0\
        );

    \I__1691\ : Odrv12
    port map (
            O => \N__7057\,
            I => \U111_CYCLE_SM.N_99_i_0\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__7054\,
            I => \U111_CYCLE_SM.N_99_i_0\
        );

    \I__1689\ : SRMux
    port map (
            O => \N__7047\,
            I => \N__7043\
        );

    \I__1688\ : SRMux
    port map (
            O => \N__7046\,
            I => \N__7040\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__7043\,
            I => \N__7036\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__7040\,
            I => \N__7033\
        );

    \I__1685\ : SRMux
    port map (
            O => \N__7039\,
            I => \N__7030\
        );

    \I__1684\ : Span4Mux_h
    port map (
            O => \N__7036\,
            I => \N__7027\
        );

    \I__1683\ : Span4Mux_h
    port map (
            O => \N__7033\,
            I => \N__7024\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__7030\,
            I => \N__7021\
        );

    \I__1681\ : Odrv4
    port map (
            O => \N__7027\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__7024\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\
        );

    \I__1679\ : Odrv12
    port map (
            O => \N__7021\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\
        );

    \I__1678\ : InMux
    port map (
            O => \N__7014\,
            I => \N__7011\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__7011\,
            I => \N__7008\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__7008\,
            I => \N__7003\
        );

    \I__1675\ : InMux
    port map (
            O => \N__7007\,
            I => \N__7000\
        );

    \I__1674\ : InMux
    port map (
            O => \N__7006\,
            I => \N__6997\
        );

    \I__1673\ : Sp12to4
    port map (
            O => \N__7003\,
            I => \N__6994\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__7000\,
            I => \N__6989\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__6997\,
            I => \N__6989\
        );

    \I__1670\ : Span12Mux_h
    port map (
            O => \N__6994\,
            I => \N__6986\
        );

    \I__1669\ : Span12Mux_v
    port map (
            O => \N__6989\,
            I => \N__6983\
        );

    \I__1668\ : Span12Mux_v
    port map (
            O => \N__6986\,
            I => \N__6980\
        );

    \I__1667\ : Span12Mux_h
    port map (
            O => \N__6983\,
            I => \N__6977\
        );

    \I__1666\ : Odrv12
    port map (
            O => \N__6980\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__1665\ : Odrv12
    port map (
            O => \N__6977\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__1664\ : InMux
    port map (
            O => \N__6972\,
            I => \N__6969\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__6969\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\
        );

    \I__1662\ : IoInMux
    port map (
            O => \N__6966\,
            I => \N__6963\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__6963\,
            I => \N__6960\
        );

    \I__1660\ : Span4Mux_s2_h
    port map (
            O => \N__6960\,
            I => \N__6957\
        );

    \I__1659\ : Sp12to4
    port map (
            O => \N__6957\,
            I => \N__6954\
        );

    \I__1658\ : Span12Mux_s11_v
    port map (
            O => \N__6954\,
            I => \N__6951\
        );

    \I__1657\ : Span12Mux_h
    port map (
            O => \N__6951\,
            I => \N__6948\
        );

    \I__1656\ : Odrv12
    port map (
            O => \N__6948\,
            I => \un1_D_UM_AMIGA_1\
        );

    \I__1655\ : InMux
    port map (
            O => \N__6945\,
            I => \N__6942\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__6942\,
            I => \N__6937\
        );

    \I__1653\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6934\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__6940\,
            I => \N__6931\
        );

    \I__1651\ : Span4Mux_v
    port map (
            O => \N__6937\,
            I => \N__6926\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__6934\,
            I => \N__6926\
        );

    \I__1649\ : InMux
    port map (
            O => \N__6931\,
            I => \N__6923\
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__6926\,
            I => \U111_CYCLE_SM.TA_DISZ0\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__6923\,
            I => \U111_CYCLE_SM.TA_DISZ0\
        );

    \I__1646\ : IoInMux
    port map (
            O => \N__6918\,
            I => \N__6915\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__6915\,
            I => \N__6912\
        );

    \I__1644\ : Span4Mux_s1_v
    port map (
            O => \N__6912\,
            I => \N__6909\
        );

    \I__1643\ : Span4Mux_v
    port map (
            O => \N__6909\,
            I => \N__6906\
        );

    \I__1642\ : Span4Mux_v
    port map (
            O => \N__6906\,
            I => \N__6903\
        );

    \I__1641\ : Span4Mux_v
    port map (
            O => \N__6903\,
            I => \N__6900\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__6900\,
            I => \N_64\
        );

    \I__1639\ : InMux
    port map (
            O => \N__6897\,
            I => \N__6894\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__6894\,
            I => \N__6891\
        );

    \I__1637\ : Span4Mux_v
    port map (
            O => \N__6891\,
            I => \N__6888\
        );

    \I__1636\ : Sp12to4
    port map (
            O => \N__6888\,
            I => \N__6885\
        );

    \I__1635\ : Span12Mux_h
    port map (
            O => \N__6885\,
            I => \N__6882\
        );

    \I__1634\ : Span12Mux_v
    port map (
            O => \N__6882\,
            I => \N__6879\
        );

    \I__1633\ : Odrv12
    port map (
            O => \N__6879\,
            I => \TCIn_c\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__6876\,
            I => \N__6872\
        );

    \I__1631\ : InMux
    port map (
            O => \N__6875\,
            I => \N__6869\
        );

    \I__1630\ : InMux
    port map (
            O => \N__6872\,
            I => \N__6866\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__6869\,
            I => \N__6863\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__6866\,
            I => \N__6858\
        );

    \I__1627\ : Span4Mux_v
    port map (
            O => \N__6863\,
            I => \N__6855\
        );

    \I__1626\ : InMux
    port map (
            O => \N__6862\,
            I => \N__6850\
        );

    \I__1625\ : InMux
    port map (
            O => \N__6861\,
            I => \N__6850\
        );

    \I__1624\ : Span4Mux_v
    port map (
            O => \N__6858\,
            I => \N__6846\
        );

    \I__1623\ : Span4Mux_v
    port map (
            O => \N__6855\,
            I => \N__6843\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__6850\,
            I => \N__6840\
        );

    \I__1621\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6836\
        );

    \I__1620\ : Span4Mux_v
    port map (
            O => \N__6846\,
            I => \N__6832\
        );

    \I__1619\ : Sp12to4
    port map (
            O => \N__6843\,
            I => \N__6829\
        );

    \I__1618\ : Span4Mux_h
    port map (
            O => \N__6840\,
            I => \N__6826\
        );

    \I__1617\ : InMux
    port map (
            O => \N__6839\,
            I => \N__6823\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__6836\,
            I => \N__6820\
        );

    \I__1615\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6817\
        );

    \I__1614\ : Sp12to4
    port map (
            O => \N__6832\,
            I => \N__6814\
        );

    \I__1613\ : Span12Mux_h
    port map (
            O => \N__6829\,
            I => \N__6807\
        );

    \I__1612\ : Sp12to4
    port map (
            O => \N__6826\,
            I => \N__6807\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__6823\,
            I => \N__6807\
        );

    \I__1610\ : Span4Mux_h
    port map (
            O => \N__6820\,
            I => \N__6802\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__6817\,
            I => \N__6802\
        );

    \I__1608\ : Span12Mux_h
    port map (
            O => \N__6814\,
            I => \N__6797\
        );

    \I__1607\ : Span12Mux_v
    port map (
            O => \N__6807\,
            I => \N__6797\
        );

    \I__1606\ : Span4Mux_v
    port map (
            O => \N__6802\,
            I => \N__6794\
        );

    \I__1605\ : Odrv12
    port map (
            O => \N__6797\,
            I => \LBENn_c\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__6794\,
            I => \LBENn_c\
        );

    \I__1603\ : IoInMux
    port map (
            O => \N__6789\,
            I => \N__6786\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__6786\,
            I => \N__6783\
        );

    \I__1601\ : Span4Mux_s3_h
    port map (
            O => \N__6783\,
            I => \N__6780\
        );

    \I__1600\ : Span4Mux_v
    port map (
            O => \N__6780\,
            I => \N__6777\
        );

    \I__1599\ : Span4Mux_v
    port map (
            O => \N__6777\,
            I => \N__6774\
        );

    \I__1598\ : Sp12to4
    port map (
            O => \N__6774\,
            I => \N__6771\
        );

    \I__1597\ : Odrv12
    port map (
            O => \N__6771\,
            I => \U111_CYCLE_SM_TCI_CPUn_0_i\
        );

    \I__1596\ : IoInMux
    port map (
            O => \N__6768\,
            I => \N__6765\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__6765\,
            I => \N__6762\
        );

    \I__1594\ : Span4Mux_s2_v
    port map (
            O => \N__6762\,
            I => \N__6759\
        );

    \I__1593\ : Span4Mux_h
    port map (
            O => \N__6759\,
            I => \N__6756\
        );

    \I__1592\ : Span4Mux_h
    port map (
            O => \N__6756\,
            I => \N__6753\
        );

    \I__1591\ : Span4Mux_v
    port map (
            O => \N__6753\,
            I => \N__6750\
        );

    \I__1590\ : Odrv4
    port map (
            O => \N__6750\,
            I => \un1_D_UU_AMIGA_0\
        );

    \I__1589\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6744\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__6744\,
            I => \N__6740\
        );

    \I__1587\ : InMux
    port map (
            O => \N__6743\,
            I => \N__6737\
        );

    \I__1586\ : Odrv12
    port map (
            O => \N__6740\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__6737\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__6732\,
            I => \N__6729\
        );

    \I__1583\ : InMux
    port map (
            O => \N__6729\,
            I => \N__6725\
        );

    \I__1582\ : InMux
    port map (
            O => \N__6728\,
            I => \N__6722\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__6725\,
            I => \N__6719\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__6722\,
            I => \N__6715\
        );

    \I__1579\ : Span4Mux_v
    port map (
            O => \N__6719\,
            I => \N__6712\
        );

    \I__1578\ : InMux
    port map (
            O => \N__6718\,
            I => \N__6709\
        );

    \I__1577\ : Span4Mux_v
    port map (
            O => \N__6715\,
            I => \N__6706\
        );

    \I__1576\ : Span4Mux_v
    port map (
            O => \N__6712\,
            I => \N__6701\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__6709\,
            I => \N__6701\
        );

    \I__1574\ : Span4Mux_v
    port map (
            O => \N__6706\,
            I => \N__6698\
        );

    \I__1573\ : Span4Mux_v
    port map (
            O => \N__6701\,
            I => \N__6695\
        );

    \I__1572\ : Span4Mux_v
    port map (
            O => \N__6698\,
            I => \N__6692\
        );

    \I__1571\ : Span4Mux_h
    port map (
            O => \N__6695\,
            I => \N__6689\
        );

    \I__1570\ : Sp12to4
    port map (
            O => \N__6692\,
            I => \N__6684\
        );

    \I__1569\ : Sp12to4
    port map (
            O => \N__6689\,
            I => \N__6684\
        );

    \I__1568\ : Span12Mux_h
    port map (
            O => \N__6684\,
            I => \N__6681\
        );

    \I__1567\ : Odrv12
    port map (
            O => \N__6681\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__1566\ : IoInMux
    port map (
            O => \N__6678\,
            I => \N__6675\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__6675\,
            I => \N__6672\
        );

    \I__1564\ : IoSpan4Mux
    port map (
            O => \N__6672\,
            I => \N__6669\
        );

    \I__1563\ : IoSpan4Mux
    port map (
            O => \N__6669\,
            I => \N__6666\
        );

    \I__1562\ : IoSpan4Mux
    port map (
            O => \N__6666\,
            I => \N__6663\
        );

    \I__1561\ : Span4Mux_s2_v
    port map (
            O => \N__6663\,
            I => \N__6660\
        );

    \I__1560\ : Span4Mux_v
    port map (
            O => \N__6660\,
            I => \N__6657\
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__6657\,
            I => \N_117\
        );

    \I__1558\ : InMux
    port map (
            O => \N__6654\,
            I => \N__6651\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__6651\,
            I => \N__6648\
        );

    \I__1556\ : Span12Mux_v
    port map (
            O => \N__6648\,
            I => \N__6645\
        );

    \I__1555\ : Span12Mux_h
    port map (
            O => \N__6645\,
            I => \N__6642\
        );

    \I__1554\ : Odrv12
    port map (
            O => \N__6642\,
            I => \D_LL_AMIGA_in_0\
        );

    \I__1553\ : IoInMux
    port map (
            O => \N__6639\,
            I => \N__6636\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__6636\,
            I => \N__6633\
        );

    \I__1551\ : Span4Mux_s2_h
    port map (
            O => \N__6633\,
            I => \N__6630\
        );

    \I__1550\ : Span4Mux_h
    port map (
            O => \N__6630\,
            I => \N__6627\
        );

    \I__1549\ : Sp12to4
    port map (
            O => \N__6627\,
            I => \N__6624\
        );

    \I__1548\ : Span12Mux_s6_v
    port map (
            O => \N__6624\,
            I => \N__6621\
        );

    \I__1547\ : Odrv12
    port map (
            O => \N__6621\,
            I => \un2_D_LL_AMIGA_0\
        );

    \I__1546\ : InMux
    port map (
            O => \N__6618\,
            I => \N__6615\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__6615\,
            I => \N__6612\
        );

    \I__1544\ : Span4Mux_h
    port map (
            O => \N__6612\,
            I => \N__6609\
        );

    \I__1543\ : Span4Mux_h
    port map (
            O => \N__6609\,
            I => \N__6605\
        );

    \I__1542\ : InMux
    port map (
            O => \N__6608\,
            I => \N__6602\
        );

    \I__1541\ : Sp12to4
    port map (
            O => \N__6605\,
            I => \N__6599\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__6602\,
            I => \N__6596\
        );

    \I__1539\ : Span12Mux_v
    port map (
            O => \N__6599\,
            I => \N__6591\
        );

    \I__1538\ : Span12Mux_h
    port map (
            O => \N__6596\,
            I => \N__6591\
        );

    \I__1537\ : Odrv12
    port map (
            O => \N__6591\,
            I => \TBIn_c\
        );

    \I__1536\ : IoInMux
    port map (
            O => \N__6588\,
            I => \N__6585\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__6585\,
            I => \N__6582\
        );

    \I__1534\ : Span12Mux_s6_v
    port map (
            O => \N__6582\,
            I => \N__6579\
        );

    \I__1533\ : Odrv12
    port map (
            O => \N__6579\,
            I => \U111_CYCLE_SM_TBI_CPUn_0_i\
        );

    \I__1532\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6573\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__6573\,
            I => \N__6570\
        );

    \I__1530\ : Span4Mux_v
    port map (
            O => \N__6570\,
            I => \N__6567\
        );

    \I__1529\ : Sp12to4
    port map (
            O => \N__6567\,
            I => \N__6564\
        );

    \I__1528\ : Span12Mux_h
    port map (
            O => \N__6564\,
            I => \N__6561\
        );

    \I__1527\ : Odrv12
    port map (
            O => \N__6561\,
            I => \D_LL_AMIGA_in_6\
        );

    \I__1526\ : IoInMux
    port map (
            O => \N__6558\,
            I => \N__6555\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__6555\,
            I => \N__6552\
        );

    \I__1524\ : Span4Mux_s3_h
    port map (
            O => \N__6552\,
            I => \N__6549\
        );

    \I__1523\ : Span4Mux_v
    port map (
            O => \N__6549\,
            I => \N__6546\
        );

    \I__1522\ : Span4Mux_v
    port map (
            O => \N__6546\,
            I => \N__6543\
        );

    \I__1521\ : Sp12to4
    port map (
            O => \N__6543\,
            I => \N__6540\
        );

    \I__1520\ : Odrv12
    port map (
            O => \N__6540\,
            I => \un2_D_LL_AMIGA_6\
        );

    \I__1519\ : IoInMux
    port map (
            O => \N__6537\,
            I => \N__6534\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__6534\,
            I => \N__6531\
        );

    \I__1517\ : Span12Mux_s3_h
    port map (
            O => \N__6531\,
            I => \N__6528\
        );

    \I__1516\ : Odrv12
    port map (
            O => \N__6528\,
            I => \un1_D_UM_AMIGA_2\
        );

    \I__1515\ : IoInMux
    port map (
            O => \N__6525\,
            I => \N__6522\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__6522\,
            I => \N__6519\
        );

    \I__1513\ : IoSpan4Mux
    port map (
            O => \N__6519\,
            I => \N__6516\
        );

    \I__1512\ : Span4Mux_s3_h
    port map (
            O => \N__6516\,
            I => \N__6513\
        );

    \I__1511\ : Span4Mux_h
    port map (
            O => \N__6513\,
            I => \N__6510\
        );

    \I__1510\ : Span4Mux_h
    port map (
            O => \N__6510\,
            I => \N__6507\
        );

    \I__1509\ : Odrv4
    port map (
            O => \N__6507\,
            I => \un1_D_UM_AMIGA_0\
        );

    \I__1508\ : InMux
    port map (
            O => \N__6504\,
            I => \N__6499\
        );

    \I__1507\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6495\
        );

    \I__1506\ : InMux
    port map (
            O => \N__6502\,
            I => \N__6492\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__6499\,
            I => \N__6488\
        );

    \I__1504\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6485\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__6495\,
            I => \N__6481\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__6492\,
            I => \N__6478\
        );

    \I__1501\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6475\
        );

    \I__1500\ : Span4Mux_v
    port map (
            O => \N__6488\,
            I => \N__6472\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__6485\,
            I => \N__6469\
        );

    \I__1498\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6466\
        );

    \I__1497\ : Span4Mux_v
    port map (
            O => \N__6481\,
            I => \N__6459\
        );

    \I__1496\ : Span4Mux_h
    port map (
            O => \N__6478\,
            I => \N__6459\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__6475\,
            I => \N__6459\
        );

    \I__1494\ : Span4Mux_h
    port map (
            O => \N__6472\,
            I => \N__6452\
        );

    \I__1493\ : Span4Mux_v
    port map (
            O => \N__6469\,
            I => \N__6452\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__6466\,
            I => \N__6452\
        );

    \I__1491\ : Span4Mux_v
    port map (
            O => \N__6459\,
            I => \N__6449\
        );

    \I__1490\ : Span4Mux_v
    port map (
            O => \N__6452\,
            I => \N__6446\
        );

    \I__1489\ : Sp12to4
    port map (
            O => \N__6449\,
            I => \N__6443\
        );

    \I__1488\ : Span4Mux_h
    port map (
            O => \N__6446\,
            I => \N__6440\
        );

    \I__1487\ : Span12Mux_h
    port map (
            O => \N__6443\,
            I => \N__6435\
        );

    \I__1486\ : Sp12to4
    port map (
            O => \N__6440\,
            I => \N__6435\
        );

    \I__1485\ : Odrv12
    port map (
            O => \N__6435\,
            I => \TEAn_c\
        );

    \I__1484\ : IoInMux
    port map (
            O => \N__6432\,
            I => \N__6429\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__6429\,
            I => \N__6426\
        );

    \I__1482\ : IoSpan4Mux
    port map (
            O => \N__6426\,
            I => \N__6423\
        );

    \I__1481\ : Span4Mux_s3_v
    port map (
            O => \N__6423\,
            I => \N__6420\
        );

    \I__1480\ : Sp12to4
    port map (
            O => \N__6420\,
            I => \N__6417\
        );

    \I__1479\ : Span12Mux_v
    port map (
            O => \N__6417\,
            I => \N__6414\
        );

    \I__1478\ : Odrv12
    port map (
            O => \N__6414\,
            I => \U111_CYCLE_SM_TEA_CPUn_0_i\
        );

    \I__1477\ : InMux
    port map (
            O => \N__6411\,
            I => \N__6408\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__6408\,
            I => \N__6405\
        );

    \I__1475\ : Span4Mux_v
    port map (
            O => \N__6405\,
            I => \N__6402\
        );

    \I__1474\ : Span4Mux_v
    port map (
            O => \N__6402\,
            I => \N__6397\
        );

    \I__1473\ : InMux
    port map (
            O => \N__6401\,
            I => \N__6394\
        );

    \I__1472\ : InMux
    port map (
            O => \N__6400\,
            I => \N__6391\
        );

    \I__1471\ : Span4Mux_v
    port map (
            O => \N__6397\,
            I => \N__6388\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__6394\,
            I => \N__6383\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__6391\,
            I => \N__6383\
        );

    \I__1468\ : Sp12to4
    port map (
            O => \N__6388\,
            I => \N__6378\
        );

    \I__1467\ : Span12Mux_v
    port map (
            O => \N__6383\,
            I => \N__6378\
        );

    \I__1466\ : Span12Mux_h
    port map (
            O => \N__6378\,
            I => \N__6375\
        );

    \I__1465\ : Odrv12
    port map (
            O => \N__6375\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__1464\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6369\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__6369\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\
        );

    \I__1462\ : InMux
    port map (
            O => \N__6366\,
            I => \N__6362\
        );

    \I__1461\ : InMux
    port map (
            O => \N__6365\,
            I => \N__6358\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__6362\,
            I => \N__6355\
        );

    \I__1459\ : InMux
    port map (
            O => \N__6361\,
            I => \N__6352\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__6358\,
            I => \U111_CYCLE_SM.un4_TS_OUT_i_0\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__6355\,
            I => \U111_CYCLE_SM.un4_TS_OUT_i_0\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__6352\,
            I => \U111_CYCLE_SM.un4_TS_OUT_i_0\
        );

    \I__1455\ : InMux
    port map (
            O => \N__6345\,
            I => \N__6341\
        );

    \I__1454\ : InMux
    port map (
            O => \N__6344\,
            I => \N__6338\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__6341\,
            I => \N__6330\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__6338\,
            I => \N__6327\
        );

    \I__1451\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6324\
        );

    \I__1450\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6321\
        );

    \I__1449\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6318\
        );

    \I__1448\ : InMux
    port map (
            O => \N__6334\,
            I => \N__6313\
        );

    \I__1447\ : InMux
    port map (
            O => \N__6333\,
            I => \N__6313\
        );

    \I__1446\ : Odrv4
    port map (
            O => \N__6330\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1445\ : Odrv4
    port map (
            O => \N__6327\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__6324\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__6321\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__6318\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__6313\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1440\ : SRMux
    port map (
            O => \N__6300\,
            I => \N__6276\
        );

    \I__1439\ : SRMux
    port map (
            O => \N__6299\,
            I => \N__6276\
        );

    \I__1438\ : SRMux
    port map (
            O => \N__6298\,
            I => \N__6276\
        );

    \I__1437\ : SRMux
    port map (
            O => \N__6297\,
            I => \N__6276\
        );

    \I__1436\ : SRMux
    port map (
            O => \N__6296\,
            I => \N__6276\
        );

    \I__1435\ : SRMux
    port map (
            O => \N__6295\,
            I => \N__6276\
        );

    \I__1434\ : SRMux
    port map (
            O => \N__6294\,
            I => \N__6276\
        );

    \I__1433\ : SRMux
    port map (
            O => \N__6293\,
            I => \N__6276\
        );

    \I__1432\ : GlobalMux
    port map (
            O => \N__6276\,
            I => \N__6273\
        );

    \I__1431\ : gio2CtrlBuf
    port map (
            O => \N__6273\,
            I => \RESETn_c_i_g\
        );

    \I__1430\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6264\
        );

    \I__1429\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6264\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__6264\,
            I => \N__6259\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6263\,
            I => \N__6256\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6262\,
            I => \N__6249\
        );

    \I__1425\ : Span4Mux_v
    port map (
            O => \N__6259\,
            I => \N__6244\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__6256\,
            I => \N__6244\
        );

    \I__1423\ : InMux
    port map (
            O => \N__6255\,
            I => \N__6239\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6254\,
            I => \N__6239\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6253\,
            I => \N__6234\
        );

    \I__1420\ : InMux
    port map (
            O => \N__6252\,
            I => \N__6234\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__6249\,
            I => \N__6231\
        );

    \I__1418\ : Span4Mux_h
    port map (
            O => \N__6244\,
            I => \N__6224\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__6239\,
            I => \N__6224\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__6234\,
            I => \N__6224\
        );

    \I__1415\ : Span4Mux_v
    port map (
            O => \N__6231\,
            I => \N__6221\
        );

    \I__1414\ : Span4Mux_v
    port map (
            O => \N__6224\,
            I => \N__6218\
        );

    \I__1413\ : Span4Mux_h
    port map (
            O => \N__6221\,
            I => \N__6215\
        );

    \I__1412\ : Span4Mux_h
    port map (
            O => \N__6218\,
            I => \N__6211\
        );

    \I__1411\ : Span4Mux_h
    port map (
            O => \N__6215\,
            I => \N__6208\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6205\
        );

    \I__1409\ : Span4Mux_h
    port map (
            O => \N__6211\,
            I => \N__6202\
        );

    \I__1408\ : Sp12to4
    port map (
            O => \N__6208\,
            I => \N__6197\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__6205\,
            I => \N__6197\
        );

    \I__1406\ : Sp12to4
    port map (
            O => \N__6202\,
            I => \N__6192\
        );

    \I__1405\ : Span12Mux_s7_h
    port map (
            O => \N__6197\,
            I => \N__6192\
        );

    \I__1404\ : Span12Mux_v
    port map (
            O => \N__6192\,
            I => \N__6189\
        );

    \I__1403\ : Odrv12
    port map (
            O => \N__6189\,
            I => \RESETn_c\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6186\,
            I => \N__6180\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6177\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6174\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6183\,
            I => \N__6171\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6180\,
            I => \U111_CYCLE_SM.N_99\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__6177\,
            I => \U111_CYCLE_SM.N_99\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__6174\,
            I => \U111_CYCLE_SM.N_99\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__6171\,
            I => \U111_CYCLE_SM.N_99\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__6162\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6159\,
            I => \N__6152\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6139\
        );

    \I__1391\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6139\
        );

    \I__1390\ : InMux
    port map (
            O => \N__6156\,
            I => \N__6139\
        );

    \I__1389\ : InMux
    port map (
            O => \N__6155\,
            I => \N__6139\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__6152\,
            I => \N__6136\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6151\,
            I => \N__6129\
        );

    \I__1386\ : InMux
    port map (
            O => \N__6150\,
            I => \N__6129\
        );

    \I__1385\ : InMux
    port map (
            O => \N__6149\,
            I => \N__6129\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6148\,
            I => \N__6126\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__6139\,
            I => \U111_CYCLE_SM.N_99_i\
        );

    \I__1382\ : Odrv4
    port map (
            O => \N__6136\,
            I => \U111_CYCLE_SM.N_99_i\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__6129\,
            I => \U111_CYCLE_SM.N_99_i\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__6126\,
            I => \U111_CYCLE_SM.N_99_i\
        );

    \I__1379\ : InMux
    port map (
            O => \N__6117\,
            I => \N__6114\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6114\,
            I => \N__6111\
        );

    \I__1377\ : Sp12to4
    port map (
            O => \N__6111\,
            I => \N__6108\
        );

    \I__1376\ : Span12Mux_v
    port map (
            O => \N__6108\,
            I => \N__6105\
        );

    \I__1375\ : Span12Mux_h
    port map (
            O => \N__6105\,
            I => \N__6102\
        );

    \I__1374\ : Odrv12
    port map (
            O => \N__6102\,
            I => \D_UM_040_in_1\
        );

    \I__1373\ : IoInMux
    port map (
            O => \N__6099\,
            I => \N__6095\
        );

    \I__1372\ : InMux
    port map (
            O => \N__6098\,
            I => \N__6092\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__6095\,
            I => \N__6089\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__6092\,
            I => \N__6086\
        );

    \I__1369\ : Span4Mux_s3_h
    port map (
            O => \N__6089\,
            I => \N__6083\
        );

    \I__1368\ : Span4Mux_v
    port map (
            O => \N__6086\,
            I => \N__6080\
        );

    \I__1367\ : Sp12to4
    port map (
            O => \N__6083\,
            I => \N__6077\
        );

    \I__1366\ : Span4Mux_v
    port map (
            O => \N__6080\,
            I => \N__6074\
        );

    \I__1365\ : Span12Mux_v
    port map (
            O => \N__6077\,
            I => \N__6071\
        );

    \I__1364\ : Sp12to4
    port map (
            O => \N__6074\,
            I => \N__6068\
        );

    \I__1363\ : Span12Mux_h
    port map (
            O => \N__6071\,
            I => \N__6065\
        );

    \I__1362\ : Span12Mux_h
    port map (
            O => \N__6068\,
            I => \N__6062\
        );

    \I__1361\ : Span12Mux_h
    port map (
            O => \N__6065\,
            I => \N__6057\
        );

    \I__1360\ : Span12Mux_v
    port map (
            O => \N__6062\,
            I => \N__6057\
        );

    \I__1359\ : Odrv12
    port map (
            O => \N__6057\,
            I => \D_LL_040_in_1\
        );

    \I__1358\ : IoInMux
    port map (
            O => \N__6054\,
            I => \N__6051\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__6051\,
            I => \N__6048\
        );

    \I__1356\ : Span12Mux_s4_h
    port map (
            O => \N__6048\,
            I => \N__6045\
        );

    \I__1355\ : Span12Mux_h
    port map (
            O => \N__6045\,
            I => \N__6042\
        );

    \I__1354\ : Odrv12
    port map (
            O => \N__6042\,
            I => \un1_D_UM_040_1\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__6039\,
            I => \N__6035\
        );

    \I__1352\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6032\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6029\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6032\,
            I => \N__6025\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6029\,
            I => \N__6022\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6019\
        );

    \I__1347\ : Span4Mux_v
    port map (
            O => \N__6025\,
            I => \N__6016\
        );

    \I__1346\ : Span4Mux_v
    port map (
            O => \N__6022\,
            I => \N__6011\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__6019\,
            I => \N__6011\
        );

    \I__1344\ : Span4Mux_v
    port map (
            O => \N__6016\,
            I => \N__6008\
        );

    \I__1343\ : Span4Mux_v
    port map (
            O => \N__6011\,
            I => \N__6005\
        );

    \I__1342\ : Span4Mux_v
    port map (
            O => \N__6008\,
            I => \N__6000\
        );

    \I__1341\ : Span4Mux_v
    port map (
            O => \N__6005\,
            I => \N__6000\
        );

    \I__1340\ : Sp12to4
    port map (
            O => \N__6000\,
            I => \N__5997\
        );

    \I__1339\ : Span12Mux_h
    port map (
            O => \N__5997\,
            I => \N__5994\
        );

    \I__1338\ : Odrv12
    port map (
            O => \N__5994\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__1337\ : InMux
    port map (
            O => \N__5991\,
            I => \N__5988\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__5988\,
            I => \N__5984\
        );

    \I__1335\ : InMux
    port map (
            O => \N__5987\,
            I => \N__5981\
        );

    \I__1334\ : Odrv12
    port map (
            O => \N__5984\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__5981\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__1332\ : IoInMux
    port map (
            O => \N__5976\,
            I => \N__5973\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__5973\,
            I => \N__5970\
        );

    \I__1330\ : Span4Mux_s3_h
    port map (
            O => \N__5970\,
            I => \N__5967\
        );

    \I__1329\ : Sp12to4
    port map (
            O => \N__5967\,
            I => \N__5964\
        );

    \I__1328\ : Span12Mux_v
    port map (
            O => \N__5964\,
            I => \N__5961\
        );

    \I__1327\ : Span12Mux_h
    port map (
            O => \N__5961\,
            I => \N__5958\
        );

    \I__1326\ : Odrv12
    port map (
            O => \N__5958\,
            I => \N_119\
        );

    \I__1325\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5952\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__5952\,
            I => \N__5949\
        );

    \I__1323\ : Span12Mux_v
    port map (
            O => \N__5949\,
            I => \N__5946\
        );

    \I__1322\ : Odrv12
    port map (
            O => \N__5946\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\
        );

    \I__1321\ : InMux
    port map (
            O => \N__5943\,
            I => \N__5939\
        );

    \I__1320\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5936\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__5939\,
            I => \N__5933\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__5936\,
            I => \N__5929\
        );

    \I__1317\ : Span4Mux_h
    port map (
            O => \N__5933\,
            I => \N__5926\
        );

    \I__1316\ : InMux
    port map (
            O => \N__5932\,
            I => \N__5923\
        );

    \I__1315\ : Sp12to4
    port map (
            O => \N__5929\,
            I => \N__5920\
        );

    \I__1314\ : Span4Mux_v
    port map (
            O => \N__5926\,
            I => \N__5915\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5923\,
            I => \N__5915\
        );

    \I__1312\ : Span12Mux_v
    port map (
            O => \N__5920\,
            I => \N__5912\
        );

    \I__1311\ : Sp12to4
    port map (
            O => \N__5915\,
            I => \N__5909\
        );

    \I__1310\ : Span12Mux_h
    port map (
            O => \N__5912\,
            I => \N__5906\
        );

    \I__1309\ : Span12Mux_v
    port map (
            O => \N__5909\,
            I => \N__5903\
        );

    \I__1308\ : Span12Mux_v
    port map (
            O => \N__5906\,
            I => \N__5900\
        );

    \I__1307\ : Span12Mux_h
    port map (
            O => \N__5903\,
            I => \N__5897\
        );

    \I__1306\ : Odrv12
    port map (
            O => \N__5900\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__1305\ : Odrv12
    port map (
            O => \N__5897\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__1304\ : IoInMux
    port map (
            O => \N__5892\,
            I => \N__5889\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__5889\,
            I => \N__5886\
        );

    \I__1302\ : IoSpan4Mux
    port map (
            O => \N__5886\,
            I => \N__5883\
        );

    \I__1301\ : IoSpan4Mux
    port map (
            O => \N__5883\,
            I => \N__5880\
        );

    \I__1300\ : Span4Mux_s2_v
    port map (
            O => \N__5880\,
            I => \N__5877\
        );

    \I__1299\ : Sp12to4
    port map (
            O => \N__5877\,
            I => \N__5874\
        );

    \I__1298\ : Span12Mux_s8_v
    port map (
            O => \N__5874\,
            I => \N__5871\
        );

    \I__1297\ : Odrv12
    port map (
            O => \N__5871\,
            I => \un1_D_UM_AMIGA_4\
        );

    \I__1296\ : InMux
    port map (
            O => \N__5868\,
            I => \N__5865\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__5865\,
            I => \N__5862\
        );

    \I__1294\ : Glb2LocalMux
    port map (
            O => \N__5862\,
            I => \N__5859\
        );

    \I__1293\ : GlobalMux
    port map (
            O => \N__5859\,
            I => \CLK80\
        );

    \I__1292\ : IoInMux
    port map (
            O => \N__5856\,
            I => \N__5852\
        );

    \I__1291\ : IoInMux
    port map (
            O => \N__5855\,
            I => \N__5849\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__5852\,
            I => \N__5846\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5849\,
            I => \N__5843\
        );

    \I__1288\ : Span12Mux_s4_v
    port map (
            O => \N__5846\,
            I => \N__5840\
        );

    \I__1287\ : Span12Mux_s3_h
    port map (
            O => \N__5843\,
            I => \N__5837\
        );

    \I__1286\ : Span12Mux_v
    port map (
            O => \N__5840\,
            I => \N__5832\
        );

    \I__1285\ : Span12Mux_h
    port map (
            O => \N__5837\,
            I => \N__5832\
        );

    \I__1284\ : Odrv12
    port map (
            O => \N__5832\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5829\,
            I => \N__5826\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__5826\,
            I => \N__5823\
        );

    \I__1281\ : Span12Mux_s11_v
    port map (
            O => \N__5823\,
            I => \N__5819\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5822\,
            I => \N__5816\
        );

    \I__1279\ : Odrv12
    port map (
            O => \N__5819\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5816\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__1277\ : InMux
    port map (
            O => \N__5811\,
            I => \N__5807\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__5810\,
            I => \N__5804\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__5807\,
            I => \N__5801\
        );

    \I__1274\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5798\
        );

    \I__1273\ : Span4Mux_v
    port map (
            O => \N__5801\,
            I => \N__5794\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__5798\,
            I => \N__5791\
        );

    \I__1271\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5788\
        );

    \I__1270\ : Span4Mux_v
    port map (
            O => \N__5794\,
            I => \N__5785\
        );

    \I__1269\ : Span4Mux_v
    port map (
            O => \N__5791\,
            I => \N__5782\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__5788\,
            I => \N__5779\
        );

    \I__1267\ : Span4Mux_v
    port map (
            O => \N__5785\,
            I => \N__5776\
        );

    \I__1266\ : Span4Mux_v
    port map (
            O => \N__5782\,
            I => \N__5771\
        );

    \I__1265\ : Span4Mux_v
    port map (
            O => \N__5779\,
            I => \N__5771\
        );

    \I__1264\ : Sp12to4
    port map (
            O => \N__5776\,
            I => \N__5766\
        );

    \I__1263\ : Sp12to4
    port map (
            O => \N__5771\,
            I => \N__5766\
        );

    \I__1262\ : Span12Mux_h
    port map (
            O => \N__5766\,
            I => \N__5763\
        );

    \I__1261\ : Odrv12
    port map (
            O => \N__5763\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1260\ : IoInMux
    port map (
            O => \N__5760\,
            I => \N__5757\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__5757\,
            I => \N__5754\
        );

    \I__1258\ : IoSpan4Mux
    port map (
            O => \N__5754\,
            I => \N__5750\
        );

    \I__1257\ : InMux
    port map (
            O => \N__5753\,
            I => \N__5747\
        );

    \I__1256\ : Span4Mux_s3_v
    port map (
            O => \N__5750\,
            I => \N__5744\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__5747\,
            I => \N__5741\
        );

    \I__1254\ : Sp12to4
    port map (
            O => \N__5744\,
            I => \N__5738\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__5741\,
            I => \N__5735\
        );

    \I__1252\ : Span12Mux_v
    port map (
            O => \N__5738\,
            I => \N__5732\
        );

    \I__1251\ : Span4Mux_v
    port map (
            O => \N__5735\,
            I => \N__5729\
        );

    \I__1250\ : Odrv12
    port map (
            O => \N__5732\,
            I => \TS_OUT\
        );

    \I__1249\ : Odrv4
    port map (
            O => \N__5729\,
            I => \TS_OUT\
        );

    \I__1248\ : IoInMux
    port map (
            O => \N__5724\,
            I => \N__5721\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__5721\,
            I => \N__5718\
        );

    \I__1246\ : Span4Mux_s0_v
    port map (
            O => \N__5718\,
            I => \N__5715\
        );

    \I__1245\ : Span4Mux_v
    port map (
            O => \N__5715\,
            I => \N__5712\
        );

    \I__1244\ : Span4Mux_v
    port map (
            O => \N__5712\,
            I => \N__5709\
        );

    \I__1243\ : Odrv4
    port map (
            O => \N__5709\,
            I => \TSnz\
        );

    \I__1242\ : IoInMux
    port map (
            O => \N__5706\,
            I => \N__5703\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5703\,
            I => \N__5700\
        );

    \I__1240\ : IoSpan4Mux
    port map (
            O => \N__5700\,
            I => \N__5696\
        );

    \I__1239\ : InMux
    port map (
            O => \N__5699\,
            I => \N__5693\
        );

    \I__1238\ : Span4Mux_s2_h
    port map (
            O => \N__5696\,
            I => \N__5690\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__5693\,
            I => \N__5687\
        );

    \I__1236\ : Sp12to4
    port map (
            O => \N__5690\,
            I => \N__5684\
        );

    \I__1235\ : Span4Mux_v
    port map (
            O => \N__5687\,
            I => \N__5681\
        );

    \I__1234\ : Span12Mux_h
    port map (
            O => \N__5684\,
            I => \N__5678\
        );

    \I__1233\ : Sp12to4
    port map (
            O => \N__5681\,
            I => \N__5675\
        );

    \I__1232\ : Span12Mux_h
    port map (
            O => \N__5678\,
            I => \N__5672\
        );

    \I__1231\ : Span12Mux_h
    port map (
            O => \N__5675\,
            I => \N__5669\
        );

    \I__1230\ : Odrv12
    port map (
            O => \N__5672\,
            I => \D_LM_040_in_7\
        );

    \I__1229\ : Odrv12
    port map (
            O => \N__5669\,
            I => \D_LM_040_in_7\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5661\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__5661\,
            I => \N__5658\
        );

    \I__1226\ : Span4Mux_v
    port map (
            O => \N__5658\,
            I => \N__5655\
        );

    \I__1225\ : Sp12to4
    port map (
            O => \N__5655\,
            I => \N__5652\
        );

    \I__1224\ : Span12Mux_h
    port map (
            O => \N__5652\,
            I => \N__5649\
        );

    \I__1223\ : Odrv12
    port map (
            O => \N__5649\,
            I => \D_UU_040_in_7\
        );

    \I__1222\ : IoInMux
    port map (
            O => \N__5646\,
            I => \N__5643\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5643\,
            I => \N__5640\
        );

    \I__1220\ : Span12Mux_s9_v
    port map (
            O => \N__5640\,
            I => \N__5637\
        );

    \I__1219\ : Span12Mux_h
    port map (
            O => \N__5637\,
            I => \N__5634\
        );

    \I__1218\ : Odrv12
    port map (
            O => \N__5634\,
            I => \un1_D_UU_040_7\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5631\,
            I => \N__5628\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__5628\,
            I => \N__5625\
        );

    \I__1215\ : Sp12to4
    port map (
            O => \N__5625\,
            I => \N__5621\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5624\,
            I => \N__5618\
        );

    \I__1213\ : Odrv12
    port map (
            O => \N__5621\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5618\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5613\,
            I => \N__5610\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__5610\,
            I => \N__5606\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__5609\,
            I => \N__5603\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__5606\,
            I => \N__5599\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5596\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5602\,
            I => \N__5593\
        );

    \I__1205\ : Span4Mux_v
    port map (
            O => \N__5599\,
            I => \N__5590\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__5596\,
            I => \N__5585\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__5593\,
            I => \N__5585\
        );

    \I__1202\ : Sp12to4
    port map (
            O => \N__5590\,
            I => \N__5580\
        );

    \I__1201\ : Span12Mux_v
    port map (
            O => \N__5585\,
            I => \N__5580\
        );

    \I__1200\ : Span12Mux_h
    port map (
            O => \N__5580\,
            I => \N__5577\
        );

    \I__1199\ : Odrv12
    port map (
            O => \N__5577\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__1198\ : IoInMux
    port map (
            O => \N__5574\,
            I => \N__5571\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5571\,
            I => \N__5568\
        );

    \I__1196\ : Span4Mux_s3_v
    port map (
            O => \N__5568\,
            I => \N__5565\
        );

    \I__1195\ : Span4Mux_h
    port map (
            O => \N__5565\,
            I => \N__5562\
        );

    \I__1194\ : Span4Mux_h
    port map (
            O => \N__5562\,
            I => \N__5559\
        );

    \I__1193\ : Span4Mux_h
    port map (
            O => \N__5559\,
            I => \N__5556\
        );

    \I__1192\ : Odrv4
    port map (
            O => \N__5556\,
            I => \N_114\
        );

    \I__1191\ : IoInMux
    port map (
            O => \N__5553\,
            I => \N__5550\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__5550\,
            I => \N__5547\
        );

    \I__1189\ : Span4Mux_s2_v
    port map (
            O => \N__5547\,
            I => \N__5544\
        );

    \I__1188\ : Span4Mux_v
    port map (
            O => \N__5544\,
            I => \N__5541\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__5541\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5538\,
            I => \N__5534\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5531\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__5534\,
            I => \N__5526\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5531\,
            I => \N__5526\
        );

    \I__1182\ : Span4Mux_v
    port map (
            O => \N__5526\,
            I => \N__5523\
        );

    \I__1181\ : Sp12to4
    port map (
            O => \N__5523\,
            I => \N__5520\
        );

    \I__1180\ : Span12Mux_h
    port map (
            O => \N__5520\,
            I => \N__5517\
        );

    \I__1179\ : Odrv12
    port map (
            O => \N__5517\,
            I => \BGn_c\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__5514\,
            I => \N__5511\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5511\,
            I => \N__5508\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__5508\,
            I => \N__5505\
        );

    \I__1175\ : Span4Mux_v
    port map (
            O => \N__5505\,
            I => \N__5500\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5504\,
            I => \N__5497\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5503\,
            I => \N__5494\
        );

    \I__1172\ : Odrv4
    port map (
            O => \N__5500\,
            I => \U111_CYCLE_SM.CYCLE_ENZ0\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__5497\,
            I => \U111_CYCLE_SM.CYCLE_ENZ0\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5494\,
            I => \U111_CYCLE_SM.CYCLE_ENZ0\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5483\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5486\,
            I => \N__5480\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__5483\,
            I => \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5480\,
            I => \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0\
        );

    \I__1165\ : IoInMux
    port map (
            O => \N__5475\,
            I => \N__5472\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__5472\,
            I => \N__5469\
        );

    \I__1163\ : IoSpan4Mux
    port map (
            O => \N__5469\,
            I => \N__5458\
        );

    \I__1162\ : IoInMux
    port map (
            O => \N__5468\,
            I => \N__5454\
        );

    \I__1161\ : IoInMux
    port map (
            O => \N__5467\,
            I => \N__5451\
        );

    \I__1160\ : IoInMux
    port map (
            O => \N__5466\,
            I => \N__5448\
        );

    \I__1159\ : IoInMux
    port map (
            O => \N__5465\,
            I => \N__5445\
        );

    \I__1158\ : IoInMux
    port map (
            O => \N__5464\,
            I => \N__5442\
        );

    \I__1157\ : IoInMux
    port map (
            O => \N__5463\,
            I => \N__5439\
        );

    \I__1156\ : IoInMux
    port map (
            O => \N__5462\,
            I => \N__5436\
        );

    \I__1155\ : IoInMux
    port map (
            O => \N__5461\,
            I => \N__5427\
        );

    \I__1154\ : Span4Mux_s3_h
    port map (
            O => \N__5458\,
            I => \N__5424\
        );

    \I__1153\ : IoInMux
    port map (
            O => \N__5457\,
            I => \N__5421\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5454\,
            I => \N__5408\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5451\,
            I => \N__5408\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5448\,
            I => \N__5408\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5445\,
            I => \N__5408\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__5442\,
            I => \N__5408\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__5439\,
            I => \N__5408\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5436\,
            I => \N__5405\
        );

    \I__1145\ : IoInMux
    port map (
            O => \N__5435\,
            I => \N__5402\
        );

    \I__1144\ : IoInMux
    port map (
            O => \N__5434\,
            I => \N__5399\
        );

    \I__1143\ : IoInMux
    port map (
            O => \N__5433\,
            I => \N__5392\
        );

    \I__1142\ : IoInMux
    port map (
            O => \N__5432\,
            I => \N__5389\
        );

    \I__1141\ : IoInMux
    port map (
            O => \N__5431\,
            I => \N__5386\
        );

    \I__1140\ : IoInMux
    port map (
            O => \N__5430\,
            I => \N__5383\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5427\,
            I => \N__5374\
        );

    \I__1138\ : IoSpan4Mux
    port map (
            O => \N__5424\,
            I => \N__5374\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5421\,
            I => \N__5374\
        );

    \I__1136\ : IoSpan4Mux
    port map (
            O => \N__5408\,
            I => \N__5374\
        );

    \I__1135\ : IoSpan4Mux
    port map (
            O => \N__5405\,
            I => \N__5363\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__5402\,
            I => \N__5363\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__5399\,
            I => \N__5363\
        );

    \I__1132\ : IoInMux
    port map (
            O => \N__5398\,
            I => \N__5360\
        );

    \I__1131\ : IoInMux
    port map (
            O => \N__5397\,
            I => \N__5357\
        );

    \I__1130\ : IoInMux
    port map (
            O => \N__5396\,
            I => \N__5354\
        );

    \I__1129\ : IoInMux
    port map (
            O => \N__5395\,
            I => \N__5351\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5392\,
            I => \N__5340\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5389\,
            I => \N__5340\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5386\,
            I => \N__5340\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__5383\,
            I => \N__5340\
        );

    \I__1124\ : IoSpan4Mux
    port map (
            O => \N__5374\,
            I => \N__5340\
        );

    \I__1123\ : IoInMux
    port map (
            O => \N__5373\,
            I => \N__5337\
        );

    \I__1122\ : IoInMux
    port map (
            O => \N__5372\,
            I => \N__5334\
        );

    \I__1121\ : IoInMux
    port map (
            O => \N__5371\,
            I => \N__5331\
        );

    \I__1120\ : IoInMux
    port map (
            O => \N__5370\,
            I => \N__5328\
        );

    \I__1119\ : IoSpan4Mux
    port map (
            O => \N__5363\,
            I => \N__5312\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5360\,
            I => \N__5312\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__5357\,
            I => \N__5312\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5354\,
            I => \N__5312\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__5351\,
            I => \N__5312\
        );

    \I__1114\ : IoSpan4Mux
    port map (
            O => \N__5340\,
            I => \N__5301\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__5337\,
            I => \N__5301\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__5334\,
            I => \N__5301\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__5331\,
            I => \N__5301\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__5328\,
            I => \N__5301\
        );

    \I__1109\ : IoInMux
    port map (
            O => \N__5327\,
            I => \N__5298\
        );

    \I__1108\ : IoInMux
    port map (
            O => \N__5326\,
            I => \N__5295\
        );

    \I__1107\ : IoInMux
    port map (
            O => \N__5325\,
            I => \N__5292\
        );

    \I__1106\ : IoInMux
    port map (
            O => \N__5324\,
            I => \N__5289\
        );

    \I__1105\ : IoInMux
    port map (
            O => \N__5323\,
            I => \N__5286\
        );

    \I__1104\ : IoSpan4Mux
    port map (
            O => \N__5312\,
            I => \N__5281\
        );

    \I__1103\ : IoSpan4Mux
    port map (
            O => \N__5301\,
            I => \N__5270\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5298\,
            I => \N__5270\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5295\,
            I => \N__5270\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5292\,
            I => \N__5270\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5289\,
            I => \N__5270\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5286\,
            I => \N__5267\
        );

    \I__1097\ : IoInMux
    port map (
            O => \N__5285\,
            I => \N__5263\
        );

    \I__1096\ : IoInMux
    port map (
            O => \N__5284\,
            I => \N__5260\
        );

    \I__1095\ : Span4Mux_s3_h
    port map (
            O => \N__5281\,
            I => \N__5257\
        );

    \I__1094\ : IoSpan4Mux
    port map (
            O => \N__5270\,
            I => \N__5252\
        );

    \I__1093\ : IoSpan4Mux
    port map (
            O => \N__5267\,
            I => \N__5252\
        );

    \I__1092\ : IoInMux
    port map (
            O => \N__5266\,
            I => \N__5249\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5263\,
            I => \N__5244\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__5260\,
            I => \N__5244\
        );

    \I__1089\ : Span4Mux_v
    port map (
            O => \N__5257\,
            I => \N__5239\
        );

    \I__1088\ : Span4Mux_s3_h
    port map (
            O => \N__5252\,
            I => \N__5239\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__5249\,
            I => \N__5236\
        );

    \I__1086\ : Span12Mux_s4_h
    port map (
            O => \N__5244\,
            I => \N__5233\
        );

    \I__1085\ : Sp12to4
    port map (
            O => \N__5239\,
            I => \N__5228\
        );

    \I__1084\ : Span12Mux_s4_h
    port map (
            O => \N__5236\,
            I => \N__5228\
        );

    \I__1083\ : Span12Mux_h
    port map (
            O => \N__5233\,
            I => \N__5223\
        );

    \I__1082\ : Span12Mux_h
    port map (
            O => \N__5228\,
            I => \N__5223\
        );

    \I__1081\ : Odrv12
    port map (
            O => \N__5223\,
            I => \U111_CYCLE_SM_OFFBOARD_EN_0\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5216\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5219\,
            I => \N__5213\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__5216\,
            I => \U111_CYCLE_SM.TS_DELAYZ0\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5213\,
            I => \U111_CYCLE_SM.TS_DELAYZ0\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__5208\,
            I => \U111_CYCLE_SM.un4_TS_OUT_i_0_cascade_\
        );

    \I__1075\ : IoInMux
    port map (
            O => \N__5205\,
            I => \N__5202\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__5202\,
            I => \N__5199\
        );

    \I__1073\ : Span4Mux_s1_v
    port map (
            O => \N__5199\,
            I => \N__5196\
        );

    \I__1072\ : Span4Mux_h
    port map (
            O => \N__5196\,
            I => \N__5193\
        );

    \I__1071\ : Span4Mux_v
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__1070\ : Span4Mux_v
    port map (
            O => \N__5190\,
            I => \N__5186\
        );

    \I__1069\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5183\
        );

    \I__1068\ : Span4Mux_v
    port map (
            O => \N__5186\,
            I => \N__5176\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__5183\,
            I => \N__5176\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5173\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5170\
        );

    \I__1064\ : Span4Mux_v
    port map (
            O => \N__5176\,
            I => \N__5163\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__5173\,
            I => \N__5163\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__5170\,
            I => \N__5163\
        );

    \I__1061\ : Span4Mux_v
    port map (
            O => \N__5163\,
            I => \N__5159\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__5162\,
            I => \N__5155\
        );

    \I__1059\ : Sp12to4
    port map (
            O => \N__5159\,
            I => \N__5151\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5146\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5146\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5154\,
            I => \N__5143\
        );

    \I__1055\ : Span12Mux_h
    port map (
            O => \N__5151\,
            I => \N__5136\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5146\,
            I => \N__5136\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__5143\,
            I => \N__5136\
        );

    \I__1052\ : Span12Mux_v
    port map (
            O => \N__5136\,
            I => \N__5133\
        );

    \I__1051\ : Odrv12
    port map (
            O => \N__5133\,
            I => \TACKn_in\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5130\,
            I => \N__5123\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5120\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5128\,
            I => \N__5115\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5127\,
            I => \N__5115\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5126\,
            I => \N__5112\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5123\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__5120\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5115\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5112\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__5103\,
            I => \U111_CYCLE_SM.N_99_cascade_\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__5100\,
            I => \N__5097\
        );

    \I__1039\ : InMux
    port map (
            O => \N__5097\,
            I => \N__5088\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5088\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5095\,
            I => \N__5085\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5081\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5093\,
            I => \N__5078\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5088\,
            I => \N__5075\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__5085\,
            I => \N__5072\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5084\,
            I => \N__5069\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__5081\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5078\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1029\ : Odrv4
    port map (
            O => \N__5075\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1028\ : Odrv4
    port map (
            O => \N__5072\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5069\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5058\,
            I => \N__5055\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5055\,
            I => \U111_CYCLE_SM.N_51\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__5052\,
            I => \N__5045\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5040\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5037\
        );

    \I__1021\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5026\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5048\,
            I => \N__5026\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5045\,
            I => \N__5026\
        );

    \I__1018\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5026\
        );

    \I__1017\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5026\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5040\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5037\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5026\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1013\ : IoInMux
    port map (
            O => \N__5019\,
            I => \N__5016\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5016\,
            I => \N__5013\
        );

    \I__1011\ : Span4Mux_s3_h
    port map (
            O => \N__5013\,
            I => \N__5009\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5012\,
            I => \N__5006\
        );

    \I__1009\ : Sp12to4
    port map (
            O => \N__5009\,
            I => \N__5003\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5006\,
            I => \N__5000\
        );

    \I__1007\ : Span12Mux_v
    port map (
            O => \N__5003\,
            I => \N__4997\
        );

    \I__1006\ : Span12Mux_v
    port map (
            O => \N__5000\,
            I => \N__4994\
        );

    \I__1005\ : Span12Mux_h
    port map (
            O => \N__4997\,
            I => \N__4989\
        );

    \I__1004\ : Span12Mux_v
    port map (
            O => \N__4994\,
            I => \N__4989\
        );

    \I__1003\ : Span12Mux_h
    port map (
            O => \N__4989\,
            I => \N__4986\
        );

    \I__1002\ : Odrv12
    port map (
            O => \N__4986\,
            I => \D_LM_040_in_1\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4983\,
            I => \N__4980\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4980\,
            I => \N__4977\
        );

    \I__999\ : Span12Mux_v
    port map (
            O => \N__4977\,
            I => \N__4974\
        );

    \I__998\ : Span12Mux_h
    port map (
            O => \N__4974\,
            I => \N__4971\
        );

    \I__997\ : Odrv12
    port map (
            O => \N__4971\,
            I => \D_UU_040_in_1\
        );

    \I__996\ : IoInMux
    port map (
            O => \N__4968\,
            I => \N__4965\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__4965\,
            I => \N__4962\
        );

    \I__994\ : IoSpan4Mux
    port map (
            O => \N__4962\,
            I => \N__4959\
        );

    \I__993\ : Span4Mux_s0_h
    port map (
            O => \N__4959\,
            I => \N__4956\
        );

    \I__992\ : Sp12to4
    port map (
            O => \N__4956\,
            I => \N__4953\
        );

    \I__991\ : Span12Mux_s11_h
    port map (
            O => \N__4953\,
            I => \N__4950\
        );

    \I__990\ : Odrv12
    port map (
            O => \N__4950\,
            I => \un1_D_UU_040_1\
        );

    \I__989\ : InMux
    port map (
            O => \N__4947\,
            I => \N__4944\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__4944\,
            I => \N__4941\
        );

    \I__987\ : Span4Mux_v
    port map (
            O => \N__4941\,
            I => \N__4938\
        );

    \I__986\ : Span4Mux_v
    port map (
            O => \N__4938\,
            I => \N__4934\
        );

    \I__985\ : InMux
    port map (
            O => \N__4937\,
            I => \N__4931\
        );

    \I__984\ : Odrv4
    port map (
            O => \N__4934\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4931\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__982\ : IoInMux
    port map (
            O => \N__4926\,
            I => \N__4923\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4923\,
            I => \N__4920\
        );

    \I__980\ : Span4Mux_s2_v
    port map (
            O => \N__4920\,
            I => \N__4917\
        );

    \I__979\ : Span4Mux_h
    port map (
            O => \N__4917\,
            I => \N__4914\
        );

    \I__978\ : Span4Mux_v
    port map (
            O => \N__4914\,
            I => \N__4911\
        );

    \I__977\ : Sp12to4
    port map (
            O => \N__4911\,
            I => \N__4908\
        );

    \I__976\ : Odrv12
    port map (
            O => \N__4908\,
            I => \N_115\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__4905\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_i_o2_0_5_cascade_\
        );

    \I__974\ : InMux
    port map (
            O => \N__4902\,
            I => \N__4899\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4899\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__4896\,
            I => \N__4893\
        );

    \I__971\ : InMux
    port map (
            O => \N__4893\,
            I => \N__4887\
        );

    \I__970\ : InMux
    port map (
            O => \N__4892\,
            I => \N__4884\
        );

    \I__969\ : InMux
    port map (
            O => \N__4891\,
            I => \N__4879\
        );

    \I__968\ : InMux
    port map (
            O => \N__4890\,
            I => \N__4879\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4887\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4884\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__4879\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__964\ : InMux
    port map (
            O => \N__4872\,
            I => \N__4866\
        );

    \I__963\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4863\
        );

    \I__962\ : InMux
    port map (
            O => \N__4870\,
            I => \N__4858\
        );

    \I__961\ : InMux
    port map (
            O => \N__4869\,
            I => \N__4858\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4866\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4863\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4858\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__957\ : InMux
    port map (
            O => \N__4851\,
            I => \N__4843\
        );

    \I__956\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4840\
        );

    \I__955\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4837\
        );

    \I__954\ : InMux
    port map (
            O => \N__4848\,
            I => \N__4834\
        );

    \I__953\ : InMux
    port map (
            O => \N__4847\,
            I => \N__4829\
        );

    \I__952\ : InMux
    port map (
            O => \N__4846\,
            I => \N__4829\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4843\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__4840\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4837\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4834\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4829\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__4818\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_a3_2_0_0_cascade_\
        );

    \I__945\ : InMux
    port map (
            O => \N__4815\,
            I => \N__4812\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4812\,
            I => \U111_CYCLE_SM.N_133\
        );

    \I__943\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4806\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4806\,
            I => \U111_CYCLE_SM.N_131\
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__4803\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_2_0_cascade_\
        );

    \I__940\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4797\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4797\,
            I => \N__4794\
        );

    \I__938\ : Span4Mux_h
    port map (
            O => \N__4794\,
            I => \N__4791\
        );

    \I__937\ : Sp12to4
    port map (
            O => \N__4791\,
            I => \N__4788\
        );

    \I__936\ : Span12Mux_v
    port map (
            O => \N__4788\,
            I => \N__4785\
        );

    \I__935\ : Odrv12
    port map (
            O => \N__4785\,
            I => \TS_CPUn_in\
        );

    \I__934\ : InMux
    port map (
            O => \N__4782\,
            I => \N__4779\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4779\,
            I => \N__4776\
        );

    \I__932\ : Span4Mux_v
    port map (
            O => \N__4776\,
            I => \N__4773\
        );

    \I__931\ : Sp12to4
    port map (
            O => \N__4773\,
            I => \N__4770\
        );

    \I__930\ : Span12Mux_h
    port map (
            O => \N__4770\,
            I => \N__4767\
        );

    \I__929\ : Odrv12
    port map (
            O => \N__4767\,
            I => \D_LM_AMIGA_in_4\
        );

    \I__928\ : IoInMux
    port map (
            O => \N__4764\,
            I => \N__4761\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4761\,
            I => \N__4758\
        );

    \I__926\ : IoSpan4Mux
    port map (
            O => \N__4758\,
            I => \N__4755\
        );

    \I__925\ : Span4Mux_s3_h
    port map (
            O => \N__4755\,
            I => \N__4752\
        );

    \I__924\ : Sp12to4
    port map (
            O => \N__4752\,
            I => \N__4749\
        );

    \I__923\ : Span12Mux_h
    port map (
            O => \N__4749\,
            I => \N__4746\
        );

    \I__922\ : Odrv12
    port map (
            O => \N__4746\,
            I => \N_109\
        );

    \I__921\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4740\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4740\,
            I => \N__4737\
        );

    \I__919\ : Span4Mux_v
    port map (
            O => \N__4737\,
            I => \N__4734\
        );

    \I__918\ : Sp12to4
    port map (
            O => \N__4734\,
            I => \N__4731\
        );

    \I__917\ : Span12Mux_h
    port map (
            O => \N__4731\,
            I => \N__4728\
        );

    \I__916\ : Odrv12
    port map (
            O => \N__4728\,
            I => \D_UU_040_in_2\
        );

    \I__915\ : IoInMux
    port map (
            O => \N__4725\,
            I => \N__4721\
        );

    \I__914\ : InMux
    port map (
            O => \N__4724\,
            I => \N__4718\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4721\,
            I => \N__4715\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__4718\,
            I => \N__4712\
        );

    \I__911\ : Span4Mux_s2_h
    port map (
            O => \N__4715\,
            I => \N__4709\
        );

    \I__910\ : Span4Mux_h
    port map (
            O => \N__4712\,
            I => \N__4706\
        );

    \I__909\ : Sp12to4
    port map (
            O => \N__4709\,
            I => \N__4703\
        );

    \I__908\ : Sp12to4
    port map (
            O => \N__4706\,
            I => \N__4700\
        );

    \I__907\ : Span12Mux_h
    port map (
            O => \N__4703\,
            I => \N__4697\
        );

    \I__906\ : Span12Mux_v
    port map (
            O => \N__4700\,
            I => \N__4694\
        );

    \I__905\ : Span12Mux_h
    port map (
            O => \N__4697\,
            I => \N__4691\
        );

    \I__904\ : Span12Mux_v
    port map (
            O => \N__4694\,
            I => \N__4688\
        );

    \I__903\ : Span12Mux_v
    port map (
            O => \N__4691\,
            I => \N__4685\
        );

    \I__902\ : Span12Mux_h
    port map (
            O => \N__4688\,
            I => \N__4682\
        );

    \I__901\ : Odrv12
    port map (
            O => \N__4685\,
            I => \D_LM_040_in_2\
        );

    \I__900\ : Odrv12
    port map (
            O => \N__4682\,
            I => \D_LM_040_in_2\
        );

    \I__899\ : IoInMux
    port map (
            O => \N__4677\,
            I => \N__4674\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4674\,
            I => \N__4671\
        );

    \I__897\ : Span4Mux_s2_v
    port map (
            O => \N__4671\,
            I => \N__4668\
        );

    \I__896\ : Span4Mux_h
    port map (
            O => \N__4668\,
            I => \N__4665\
        );

    \I__895\ : Span4Mux_h
    port map (
            O => \N__4665\,
            I => \N__4662\
        );

    \I__894\ : Span4Mux_v
    port map (
            O => \N__4662\,
            I => \N__4659\
        );

    \I__893\ : Odrv4
    port map (
            O => \N__4659\,
            I => \un1_D_UU_040_2\
        );

    \I__892\ : InMux
    port map (
            O => \N__4656\,
            I => \N__4653\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__4653\,
            I => \N__4649\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__4652\,
            I => \N__4645\
        );

    \I__889\ : Span4Mux_v
    port map (
            O => \N__4649\,
            I => \N__4642\
        );

    \I__888\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4639\
        );

    \I__887\ : InMux
    port map (
            O => \N__4645\,
            I => \N__4636\
        );

    \I__886\ : Span4Mux_v
    port map (
            O => \N__4642\,
            I => \N__4633\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4639\,
            I => \N__4630\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4636\,
            I => \N__4627\
        );

    \I__883\ : Span4Mux_v
    port map (
            O => \N__4633\,
            I => \N__4624\
        );

    \I__882\ : Span4Mux_v
    port map (
            O => \N__4630\,
            I => \N__4621\
        );

    \I__881\ : Span12Mux_h
    port map (
            O => \N__4627\,
            I => \N__4618\
        );

    \I__880\ : Sp12to4
    port map (
            O => \N__4624\,
            I => \N__4613\
        );

    \I__879\ : Sp12to4
    port map (
            O => \N__4621\,
            I => \N__4613\
        );

    \I__878\ : Span12Mux_v
    port map (
            O => \N__4618\,
            I => \N__4608\
        );

    \I__877\ : Span12Mux_h
    port map (
            O => \N__4613\,
            I => \N__4608\
        );

    \I__876\ : Odrv12
    port map (
            O => \N__4608\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__875\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4602\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__4602\,
            I => \N__4598\
        );

    \I__873\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4595\
        );

    \I__872\ : Odrv12
    port map (
            O => \N__4598\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4595\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__870\ : IoInMux
    port map (
            O => \N__4590\,
            I => \N__4587\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4587\,
            I => \N__4584\
        );

    \I__868\ : Span12Mux_s8_v
    port map (
            O => \N__4584\,
            I => \N__4581\
        );

    \I__867\ : Span12Mux_h
    port map (
            O => \N__4581\,
            I => \N__4578\
        );

    \I__866\ : Odrv12
    port map (
            O => \N__4578\,
            I => \N_118\
        );

    \I__865\ : InMux
    port map (
            O => \N__4575\,
            I => \N__4572\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4572\,
            I => \N__4569\
        );

    \I__863\ : Span12Mux_s8_v
    port map (
            O => \N__4569\,
            I => \N__4565\
        );

    \I__862\ : InMux
    port map (
            O => \N__4568\,
            I => \N__4562\
        );

    \I__861\ : Odrv12
    port map (
            O => \N__4565\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4562\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__4557\,
            I => \N__4554\
        );

    \I__858\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4551\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4551\,
            I => \N__4547\
        );

    \I__856\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4544\
        );

    \I__855\ : Span4Mux_h
    port map (
            O => \N__4547\,
            I => \N__4539\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4544\,
            I => \N__4539\
        );

    \I__853\ : Span4Mux_v
    port map (
            O => \N__4539\,
            I => \N__4535\
        );

    \I__852\ : InMux
    port map (
            O => \N__4538\,
            I => \N__4532\
        );

    \I__851\ : Span4Mux_v
    port map (
            O => \N__4535\,
            I => \N__4527\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4532\,
            I => \N__4527\
        );

    \I__849\ : Span4Mux_v
    port map (
            O => \N__4527\,
            I => \N__4524\
        );

    \I__848\ : IoSpan4Mux
    port map (
            O => \N__4524\,
            I => \N__4521\
        );

    \I__847\ : IoSpan4Mux
    port map (
            O => \N__4521\,
            I => \N__4518\
        );

    \I__846\ : Odrv4
    port map (
            O => \N__4518\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__845\ : IoInMux
    port map (
            O => \N__4515\,
            I => \N__4512\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4512\,
            I => \N__4509\
        );

    \I__843\ : Span4Mux_s2_v
    port map (
            O => \N__4509\,
            I => \N__4506\
        );

    \I__842\ : Span4Mux_h
    port map (
            O => \N__4506\,
            I => \N__4503\
        );

    \I__841\ : Span4Mux_h
    port map (
            O => \N__4503\,
            I => \N__4500\
        );

    \I__840\ : Span4Mux_v
    port map (
            O => \N__4500\,
            I => \N__4497\
        );

    \I__839\ : Odrv4
    port map (
            O => \N__4497\,
            I => \N_116\
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__4494\,
            I => \N__4490\
        );

    \I__837\ : InMux
    port map (
            O => \N__4493\,
            I => \N__4487\
        );

    \I__836\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4483\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4487\,
            I => \N__4480\
        );

    \I__834\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4477\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4483\,
            I => \N__4474\
        );

    \I__832\ : Span4Mux_v
    port map (
            O => \N__4480\,
            I => \N__4469\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4477\,
            I => \N__4469\
        );

    \I__830\ : Sp12to4
    port map (
            O => \N__4474\,
            I => \N__4466\
        );

    \I__829\ : Span4Mux_v
    port map (
            O => \N__4469\,
            I => \N__4463\
        );

    \I__828\ : Span12Mux_v
    port map (
            O => \N__4466\,
            I => \N__4458\
        );

    \I__827\ : Sp12to4
    port map (
            O => \N__4463\,
            I => \N__4458\
        );

    \I__826\ : Span12Mux_h
    port map (
            O => \N__4458\,
            I => \N__4455\
        );

    \I__825\ : Odrv12
    port map (
            O => \N__4455\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__824\ : InMux
    port map (
            O => \N__4452\,
            I => \N__4449\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__4449\,
            I => \N__4446\
        );

    \I__822\ : Span12Mux_v
    port map (
            O => \N__4446\,
            I => \N__4442\
        );

    \I__821\ : InMux
    port map (
            O => \N__4445\,
            I => \N__4439\
        );

    \I__820\ : Odrv12
    port map (
            O => \N__4442\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4439\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__818\ : IoInMux
    port map (
            O => \N__4434\,
            I => \N__4431\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4431\,
            I => \N__4428\
        );

    \I__816\ : IoSpan4Mux
    port map (
            O => \N__4428\,
            I => \N__4425\
        );

    \I__815\ : Span4Mux_s2_v
    port map (
            O => \N__4425\,
            I => \N__4422\
        );

    \I__814\ : Span4Mux_v
    port map (
            O => \N__4422\,
            I => \N__4419\
        );

    \I__813\ : Sp12to4
    port map (
            O => \N__4419\,
            I => \N__4416\
        );

    \I__812\ : Odrv12
    port map (
            O => \N__4416\,
            I => \N_113\
        );

    \I__811\ : IoInMux
    port map (
            O => \N__4413\,
            I => \N__4410\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__4410\,
            I => \N__4407\
        );

    \I__809\ : IoSpan4Mux
    port map (
            O => \N__4407\,
            I => \N__4403\
        );

    \I__808\ : InMux
    port map (
            O => \N__4406\,
            I => \N__4400\
        );

    \I__807\ : IoSpan4Mux
    port map (
            O => \N__4403\,
            I => \N__4397\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4400\,
            I => \N__4394\
        );

    \I__805\ : Span4Mux_s2_h
    port map (
            O => \N__4397\,
            I => \N__4391\
        );

    \I__804\ : Span4Mux_v
    port map (
            O => \N__4394\,
            I => \N__4388\
        );

    \I__803\ : Sp12to4
    port map (
            O => \N__4391\,
            I => \N__4385\
        );

    \I__802\ : Sp12to4
    port map (
            O => \N__4388\,
            I => \N__4382\
        );

    \I__801\ : Span12Mux_h
    port map (
            O => \N__4385\,
            I => \N__4379\
        );

    \I__800\ : Span12Mux_h
    port map (
            O => \N__4382\,
            I => \N__4376\
        );

    \I__799\ : Span12Mux_h
    port map (
            O => \N__4379\,
            I => \N__4373\
        );

    \I__798\ : Span12Mux_v
    port map (
            O => \N__4376\,
            I => \N__4370\
        );

    \I__797\ : Odrv12
    port map (
            O => \N__4373\,
            I => \D_LM_040_in_3\
        );

    \I__796\ : Odrv12
    port map (
            O => \N__4370\,
            I => \D_LM_040_in_3\
        );

    \I__795\ : InMux
    port map (
            O => \N__4365\,
            I => \N__4362\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4362\,
            I => \N__4359\
        );

    \I__793\ : Span4Mux_v
    port map (
            O => \N__4359\,
            I => \N__4356\
        );

    \I__792\ : Span4Mux_h
    port map (
            O => \N__4356\,
            I => \N__4353\
        );

    \I__791\ : Sp12to4
    port map (
            O => \N__4353\,
            I => \N__4350\
        );

    \I__790\ : Span12Mux_h
    port map (
            O => \N__4350\,
            I => \N__4347\
        );

    \I__789\ : Odrv12
    port map (
            O => \N__4347\,
            I => \D_UU_040_in_3\
        );

    \I__788\ : IoInMux
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4341\,
            I => \N__4338\
        );

    \I__786\ : Span12Mux_s1_v
    port map (
            O => \N__4338\,
            I => \N__4335\
        );

    \I__785\ : Span12Mux_h
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__784\ : Odrv12
    port map (
            O => \N__4332\,
            I => \un1_D_UU_040_3\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__4329\,
            I => \N__4326\
        );

    \I__782\ : InMux
    port map (
            O => \N__4326\,
            I => \N__4323\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__4323\,
            I => \N__4319\
        );

    \I__780\ : InMux
    port map (
            O => \N__4322\,
            I => \N__4316\
        );

    \I__779\ : Span4Mux_v
    port map (
            O => \N__4319\,
            I => \N__4313\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4316\,
            I => \N__4310\
        );

    \I__777\ : Span4Mux_h
    port map (
            O => \N__4313\,
            I => \N__4304\
        );

    \I__776\ : Span4Mux_v
    port map (
            O => \N__4310\,
            I => \N__4304\
        );

    \I__775\ : InMux
    port map (
            O => \N__4309\,
            I => \N__4301\
        );

    \I__774\ : Span4Mux_v
    port map (
            O => \N__4304\,
            I => \N__4298\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4301\,
            I => \N__4295\
        );

    \I__772\ : Span4Mux_v
    port map (
            O => \N__4298\,
            I => \N__4290\
        );

    \I__771\ : Span4Mux_h
    port map (
            O => \N__4295\,
            I => \N__4290\
        );

    \I__770\ : Span4Mux_v
    port map (
            O => \N__4290\,
            I => \N__4287\
        );

    \I__769\ : Span4Mux_h
    port map (
            O => \N__4287\,
            I => \N__4284\
        );

    \I__768\ : Span4Mux_h
    port map (
            O => \N__4284\,
            I => \N__4281\
        );

    \I__767\ : Odrv4
    port map (
            O => \N__4281\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__766\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4274\
        );

    \I__765\ : InMux
    port map (
            O => \N__4277\,
            I => \N__4271\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4274\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__4271\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\
        );

    \I__762\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4260\
        );

    \I__761\ : InMux
    port map (
            O => \N__4265\,
            I => \N__4260\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4260\,
            I => \N__4257\
        );

    \I__759\ : Span4Mux_v
    port map (
            O => \N__4257\,
            I => \N__4254\
        );

    \I__758\ : Sp12to4
    port map (
            O => \N__4254\,
            I => \N__4251\
        );

    \I__757\ : Span12Mux_h
    port map (
            O => \N__4251\,
            I => \N__4248\
        );

    \I__756\ : Span12Mux_v
    port map (
            O => \N__4248\,
            I => \N__4245\
        );

    \I__755\ : Odrv12
    port map (
            O => \N__4245\,
            I => \SIZ_c_0\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__4242\,
            I => \N__4238\
        );

    \I__753\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4233\
        );

    \I__752\ : InMux
    port map (
            O => \N__4238\,
            I => \N__4233\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4233\,
            I => \N__4230\
        );

    \I__750\ : Span4Mux_v
    port map (
            O => \N__4230\,
            I => \N__4227\
        );

    \I__749\ : Sp12to4
    port map (
            O => \N__4227\,
            I => \N__4224\
        );

    \I__748\ : Span12Mux_h
    port map (
            O => \N__4224\,
            I => \N__4221\
        );

    \I__747\ : Span12Mux_v
    port map (
            O => \N__4221\,
            I => \N__4218\
        );

    \I__746\ : Odrv12
    port map (
            O => \N__4218\,
            I => \SIZ_c_1\
        );

    \I__745\ : CascadeMux
    port map (
            O => \N__4215\,
            I => \N__4210\
        );

    \I__744\ : InMux
    port map (
            O => \N__4214\,
            I => \N__4205\
        );

    \I__743\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4205\
        );

    \I__742\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4202\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4205\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4202\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__4197\,
            I => \N__4194\
        );

    \I__738\ : InMux
    port map (
            O => \N__4194\,
            I => \N__4187\
        );

    \I__737\ : InMux
    port map (
            O => \N__4193\,
            I => \N__4187\
        );

    \I__736\ : InMux
    port map (
            O => \N__4192\,
            I => \N__4184\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__4187\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__4184\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__733\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4170\
        );

    \I__732\ : InMux
    port map (
            O => \N__4178\,
            I => \N__4170\
        );

    \I__731\ : InMux
    port map (
            O => \N__4177\,
            I => \N__4167\
        );

    \I__730\ : InMux
    port map (
            O => \N__4176\,
            I => \N__4162\
        );

    \I__729\ : InMux
    port map (
            O => \N__4175\,
            I => \N__4162\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4170\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__4167\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4162\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__725\ : InMux
    port map (
            O => \N__4155\,
            I => \N__4151\
        );

    \I__724\ : InMux
    port map (
            O => \N__4154\,
            I => \N__4148\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__4151\,
            I => \N__4143\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4148\,
            I => \N__4143\
        );

    \I__721\ : Span4Mux_v
    port map (
            O => \N__4143\,
            I => \N__4139\
        );

    \I__720\ : InMux
    port map (
            O => \N__4142\,
            I => \N__4136\
        );

    \I__719\ : Sp12to4
    port map (
            O => \N__4139\,
            I => \N__4131\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__4136\,
            I => \N__4131\
        );

    \I__717\ : Span12Mux_h
    port map (
            O => \N__4131\,
            I => \N__4128\
        );

    \I__716\ : Span12Mux_v
    port map (
            O => \N__4128\,
            I => \N__4125\
        );

    \I__715\ : Odrv12
    port map (
            O => \N__4125\,
            I => \PORTSIZE_c\
        );

    \I__714\ : InMux
    port map (
            O => \N__4122\,
            I => \N__4119\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__4119\,
            I => \U111_CYCLE_SM.N_179\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__4116\,
            I => \U111_CYCLE_SM.N_179_cascade_\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__4113\,
            I => \U111_CYCLE_SM.N_101_cascade_\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__4110\,
            I => \N__4107\
        );

    \I__709\ : InMux
    port map (
            O => \N__4107\,
            I => \N__4100\
        );

    \I__708\ : InMux
    port map (
            O => \N__4106\,
            I => \N__4100\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__4105\,
            I => \N__4097\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4100\,
            I => \N__4094\
        );

    \I__705\ : InMux
    port map (
            O => \N__4097\,
            I => \N__4091\
        );

    \I__704\ : Odrv12
    port map (
            O => \N__4094\,
            I => \U111_CYCLE_SM.N_98\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4091\,
            I => \U111_CYCLE_SM.N_98\
        );

    \I__702\ : InMux
    port map (
            O => \N__4086\,
            I => \N__4083\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__4083\,
            I => \U111_CYCLE_SM.N_10\
        );

    \I__700\ : InMux
    port map (
            O => \N__4080\,
            I => \N__4077\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__4077\,
            I => \U111_CYCLE_SM.N_101\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__4074\,
            I => \U111_CYCLE_SM.N_12_i_1_cascade_\
        );

    \I__697\ : InMux
    port map (
            O => \N__4071\,
            I => \N__4068\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__4068\,
            I => \U111_CYCLE_SM.N_55\
        );

    \I__695\ : InMux
    port map (
            O => \N__4065\,
            I => \N__4061\
        );

    \I__694\ : InMux
    port map (
            O => \N__4064\,
            I => \N__4058\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4061\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4058\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__691\ : InMux
    port map (
            O => \N__4053\,
            I => \N__4050\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4050\,
            I => \N__4047\
        );

    \I__689\ : Span4Mux_v
    port map (
            O => \N__4047\,
            I => \N__4044\
        );

    \I__688\ : Sp12to4
    port map (
            O => \N__4044\,
            I => \N__4041\
        );

    \I__687\ : Span12Mux_h
    port map (
            O => \N__4041\,
            I => \N__4038\
        );

    \I__686\ : Odrv12
    port map (
            O => \N__4038\,
            I => \D_LM_AMIGA_in_7\
        );

    \I__685\ : IoInMux
    port map (
            O => \N__4035\,
            I => \N__4032\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__4032\,
            I => \N__4029\
        );

    \I__683\ : IoSpan4Mux
    port map (
            O => \N__4029\,
            I => \N__4026\
        );

    \I__682\ : Span4Mux_s3_h
    port map (
            O => \N__4026\,
            I => \N__4023\
        );

    \I__681\ : Span4Mux_h
    port map (
            O => \N__4023\,
            I => \N__4020\
        );

    \I__680\ : Sp12to4
    port map (
            O => \N__4020\,
            I => \N__4017\
        );

    \I__679\ : Odrv12
    port map (
            O => \N__4017\,
            I => \N_106\
        );

    \I__678\ : InMux
    port map (
            O => \N__4014\,
            I => \N__4011\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4011\,
            I => \N__4008\
        );

    \I__676\ : Span12Mux_v
    port map (
            O => \N__4008\,
            I => \N__4005\
        );

    \I__675\ : Span12Mux_h
    port map (
            O => \N__4005\,
            I => \N__4002\
        );

    \I__674\ : Odrv12
    port map (
            O => \N__4002\,
            I => \D_LM_AMIGA_in_6\
        );

    \I__673\ : IoInMux
    port map (
            O => \N__3999\,
            I => \N__3996\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3996\,
            I => \N__3993\
        );

    \I__671\ : IoSpan4Mux
    port map (
            O => \N__3993\,
            I => \N__3990\
        );

    \I__670\ : Sp12to4
    port map (
            O => \N__3990\,
            I => \N__3987\
        );

    \I__669\ : Span12Mux_s9_h
    port map (
            O => \N__3987\,
            I => \N__3984\
        );

    \I__668\ : Odrv12
    port map (
            O => \N__3984\,
            I => \N_107\
        );

    \I__667\ : InMux
    port map (
            O => \N__3981\,
            I => \N__3978\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__3978\,
            I => \N__3975\
        );

    \I__665\ : Span12Mux_v
    port map (
            O => \N__3975\,
            I => \N__3972\
        );

    \I__664\ : Span12Mux_h
    port map (
            O => \N__3972\,
            I => \N__3969\
        );

    \I__663\ : Odrv12
    port map (
            O => \N__3969\,
            I => \D_UM_040_in_3\
        );

    \I__662\ : InMux
    port map (
            O => \N__3966\,
            I => \N__3962\
        );

    \I__661\ : IoInMux
    port map (
            O => \N__3965\,
            I => \N__3959\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3962\,
            I => \N__3956\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3959\,
            I => \N__3953\
        );

    \I__658\ : Span4Mux_v
    port map (
            O => \N__3956\,
            I => \N__3950\
        );

    \I__657\ : Span4Mux_s3_h
    port map (
            O => \N__3953\,
            I => \N__3947\
        );

    \I__656\ : Sp12to4
    port map (
            O => \N__3950\,
            I => \N__3944\
        );

    \I__655\ : Sp12to4
    port map (
            O => \N__3947\,
            I => \N__3941\
        );

    \I__654\ : Span12Mux_h
    port map (
            O => \N__3944\,
            I => \N__3938\
        );

    \I__653\ : Span12Mux_v
    port map (
            O => \N__3941\,
            I => \N__3935\
        );

    \I__652\ : Span12Mux_v
    port map (
            O => \N__3938\,
            I => \N__3932\
        );

    \I__651\ : Span12Mux_h
    port map (
            O => \N__3935\,
            I => \N__3929\
        );

    \I__650\ : Span12Mux_v
    port map (
            O => \N__3932\,
            I => \N__3924\
        );

    \I__649\ : Span12Mux_h
    port map (
            O => \N__3929\,
            I => \N__3924\
        );

    \I__648\ : Odrv12
    port map (
            O => \N__3924\,
            I => \D_LL_040_in_3\
        );

    \I__647\ : IoInMux
    port map (
            O => \N__3921\,
            I => \N__3918\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3918\,
            I => \N__3915\
        );

    \I__645\ : IoSpan4Mux
    port map (
            O => \N__3915\,
            I => \N__3912\
        );

    \I__644\ : Span4Mux_s2_h
    port map (
            O => \N__3912\,
            I => \N__3909\
        );

    \I__643\ : Sp12to4
    port map (
            O => \N__3909\,
            I => \N__3906\
        );

    \I__642\ : Odrv12
    port map (
            O => \N__3906\,
            I => \un1_D_UM_040_3\
        );

    \I__641\ : InMux
    port map (
            O => \N__3903\,
            I => \N__3900\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3900\,
            I => \N__3897\
        );

    \I__639\ : Span4Mux_v
    port map (
            O => \N__3897\,
            I => \N__3894\
        );

    \I__638\ : Span4Mux_h
    port map (
            O => \N__3894\,
            I => \N__3891\
        );

    \I__637\ : Sp12to4
    port map (
            O => \N__3891\,
            I => \N__3888\
        );

    \I__636\ : Odrv12
    port map (
            O => \N__3888\,
            I => \D_LL_AMIGA_in_3\
        );

    \I__635\ : IoInMux
    port map (
            O => \N__3885\,
            I => \N__3882\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3882\,
            I => \N__3879\
        );

    \I__633\ : Span4Mux_s2_h
    port map (
            O => \N__3879\,
            I => \N__3876\
        );

    \I__632\ : Span4Mux_v
    port map (
            O => \N__3876\,
            I => \N__3873\
        );

    \I__631\ : Span4Mux_h
    port map (
            O => \N__3873\,
            I => \N__3870\
        );

    \I__630\ : Sp12to4
    port map (
            O => \N__3870\,
            I => \N__3867\
        );

    \I__629\ : Span12Mux_h
    port map (
            O => \N__3867\,
            I => \N__3864\
        );

    \I__628\ : Odrv12
    port map (
            O => \N__3864\,
            I => \un2_D_LL_AMIGA_3\
        );

    \I__627\ : IoInMux
    port map (
            O => \N__3861\,
            I => \N__3858\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3858\,
            I => \N__3855\
        );

    \I__625\ : Odrv12
    port map (
            O => \N__3855\,
            I => \LBENn_c_i\
        );

    \I__624\ : InMux
    port map (
            O => \N__3852\,
            I => \N__3849\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3849\,
            I => \N__3846\
        );

    \I__622\ : Span4Mux_v
    port map (
            O => \N__3846\,
            I => \N__3843\
        );

    \I__621\ : Sp12to4
    port map (
            O => \N__3843\,
            I => \N__3840\
        );

    \I__620\ : Span12Mux_h
    port map (
            O => \N__3840\,
            I => \N__3837\
        );

    \I__619\ : Odrv12
    port map (
            O => \N__3837\,
            I => \D_LM_AMIGA_in_0\
        );

    \I__618\ : IoInMux
    port map (
            O => \N__3834\,
            I => \N__3831\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__3831\,
            I => \N__3828\
        );

    \I__616\ : IoSpan4Mux
    port map (
            O => \N__3828\,
            I => \N__3825\
        );

    \I__615\ : Span4Mux_s3_h
    port map (
            O => \N__3825\,
            I => \N__3822\
        );

    \I__614\ : Sp12to4
    port map (
            O => \N__3822\,
            I => \N__3819\
        );

    \I__613\ : Span12Mux_h
    port map (
            O => \N__3819\,
            I => \N__3816\
        );

    \I__612\ : Odrv12
    port map (
            O => \N__3816\,
            I => \un2_D_LM_AMIGA_0\
        );

    \I__611\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3807\
        );

    \I__610\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3807\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3807\,
            I => \N__3804\
        );

    \I__608\ : Span4Mux_h
    port map (
            O => \N__3804\,
            I => \N__3801\
        );

    \I__607\ : Span4Mux_v
    port map (
            O => \N__3801\,
            I => \N__3798\
        );

    \I__606\ : Span4Mux_h
    port map (
            O => \N__3798\,
            I => \N__3794\
        );

    \I__605\ : InMux
    port map (
            O => \N__3797\,
            I => \N__3791\
        );

    \I__604\ : Odrv4
    port map (
            O => \N__3794\,
            I => \U111_CYCLE_SM.A2_ENZ0\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3791\,
            I => \U111_CYCLE_SM.A2_ENZ0\
        );

    \I__602\ : InMux
    port map (
            O => \N__3786\,
            I => \N__3783\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3783\,
            I => \N__3780\
        );

    \I__600\ : Span4Mux_v
    port map (
            O => \N__3780\,
            I => \N__3777\
        );

    \I__599\ : Sp12to4
    port map (
            O => \N__3777\,
            I => \N__3774\
        );

    \I__598\ : Span12Mux_h
    port map (
            O => \N__3774\,
            I => \N__3771\
        );

    \I__597\ : Odrv12
    port map (
            O => \N__3771\,
            I => \D_LL_AMIGA_in_2\
        );

    \I__596\ : IoInMux
    port map (
            O => \N__3768\,
            I => \N__3765\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3765\,
            I => \N__3762\
        );

    \I__594\ : Span12Mux_s7_h
    port map (
            O => \N__3762\,
            I => \N__3759\
        );

    \I__593\ : Span12Mux_h
    port map (
            O => \N__3759\,
            I => \N__3756\
        );

    \I__592\ : Odrv12
    port map (
            O => \N__3756\,
            I => \un2_D_LL_AMIGA_2\
        );

    \I__591\ : IoInMux
    port map (
            O => \N__3753\,
            I => \N__3750\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3750\,
            I => \N__3746\
        );

    \I__589\ : InMux
    port map (
            O => \N__3749\,
            I => \N__3743\
        );

    \I__588\ : IoSpan4Mux
    port map (
            O => \N__3746\,
            I => \N__3740\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3743\,
            I => \N__3737\
        );

    \I__586\ : Span4Mux_s2_h
    port map (
            O => \N__3740\,
            I => \N__3734\
        );

    \I__585\ : Span4Mux_v
    port map (
            O => \N__3737\,
            I => \N__3731\
        );

    \I__584\ : Sp12to4
    port map (
            O => \N__3734\,
            I => \N__3728\
        );

    \I__583\ : Sp12to4
    port map (
            O => \N__3731\,
            I => \N__3725\
        );

    \I__582\ : Span12Mux_h
    port map (
            O => \N__3728\,
            I => \N__3720\
        );

    \I__581\ : Span12Mux_v
    port map (
            O => \N__3725\,
            I => \N__3720\
        );

    \I__580\ : Span12Mux_h
    port map (
            O => \N__3720\,
            I => \N__3717\
        );

    \I__579\ : Odrv12
    port map (
            O => \N__3717\,
            I => \D_LL_040_in_0\
        );

    \I__578\ : InMux
    port map (
            O => \N__3714\,
            I => \N__3711\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3711\,
            I => \N__3708\
        );

    \I__576\ : Span4Mux_v
    port map (
            O => \N__3708\,
            I => \N__3705\
        );

    \I__575\ : Sp12to4
    port map (
            O => \N__3705\,
            I => \N__3702\
        );

    \I__574\ : Span12Mux_h
    port map (
            O => \N__3702\,
            I => \N__3699\
        );

    \I__573\ : Span12Mux_h
    port map (
            O => \N__3699\,
            I => \N__3696\
        );

    \I__572\ : Odrv12
    port map (
            O => \N__3696\,
            I => \D_UM_040_in_0\
        );

    \I__571\ : IoInMux
    port map (
            O => \N__3693\,
            I => \N__3690\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3690\,
            I => \N__3687\
        );

    \I__569\ : IoSpan4Mux
    port map (
            O => \N__3687\,
            I => \N__3684\
        );

    \I__568\ : Sp12to4
    port map (
            O => \N__3684\,
            I => \N__3681\
        );

    \I__567\ : Span12Mux_h
    port map (
            O => \N__3681\,
            I => \N__3678\
        );

    \I__566\ : Odrv12
    port map (
            O => \N__3678\,
            I => \un1_D_UM_040_0\
        );

    \I__565\ : InMux
    port map (
            O => \N__3675\,
            I => \N__3672\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__3672\,
            I => \N__3669\
        );

    \I__563\ : Span12Mux_h
    port map (
            O => \N__3669\,
            I => \N__3666\
        );

    \I__562\ : Odrv12
    port map (
            O => \N__3666\,
            I => \D_LM_AMIGA_in_1\
        );

    \I__561\ : IoInMux
    port map (
            O => \N__3663\,
            I => \N__3660\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3660\,
            I => \N__3657\
        );

    \I__559\ : IoSpan4Mux
    port map (
            O => \N__3657\,
            I => \N__3654\
        );

    \I__558\ : Sp12to4
    port map (
            O => \N__3654\,
            I => \N__3651\
        );

    \I__557\ : Span12Mux_s7_h
    port map (
            O => \N__3651\,
            I => \N__3648\
        );

    \I__556\ : Span12Mux_h
    port map (
            O => \N__3648\,
            I => \N__3645\
        );

    \I__555\ : Odrv12
    port map (
            O => \N__3645\,
            I => \N_112\
        );

    \I__554\ : IoInMux
    port map (
            O => \N__3642\,
            I => \N__3639\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3639\,
            I => \N__3636\
        );

    \I__552\ : Span4Mux_s2_v
    port map (
            O => \N__3636\,
            I => \N__3633\
        );

    \I__551\ : Span4Mux_h
    port map (
            O => \N__3633\,
            I => \N__3630\
        );

    \I__550\ : Span4Mux_v
    port map (
            O => \N__3630\,
            I => \N__3627\
        );

    \I__549\ : Odrv4
    port map (
            O => \N__3627\,
            I => \N_96\
        );

    \I__548\ : IoInMux
    port map (
            O => \N__3624\,
            I => \N__3621\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3621\,
            I => \N__3618\
        );

    \I__546\ : Span4Mux_s2_v
    port map (
            O => \N__3618\,
            I => \N__3615\
        );

    \I__545\ : Span4Mux_h
    port map (
            O => \N__3615\,
            I => \N__3612\
        );

    \I__544\ : Span4Mux_v
    port map (
            O => \N__3612\,
            I => \N__3609\
        );

    \I__543\ : Odrv4
    port map (
            O => \N__3609\,
            I => \N_94_i\
        );

    \I__542\ : InMux
    port map (
            O => \N__3606\,
            I => \N__3601\
        );

    \I__541\ : InMux
    port map (
            O => \N__3605\,
            I => \N__3596\
        );

    \I__540\ : InMux
    port map (
            O => \N__3604\,
            I => \N__3596\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3601\,
            I => \N__3591\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3596\,
            I => \N__3591\
        );

    \I__537\ : Span4Mux_h
    port map (
            O => \N__3591\,
            I => \N__3588\
        );

    \I__536\ : Span4Mux_v
    port map (
            O => \N__3588\,
            I => \N__3585\
        );

    \I__535\ : Odrv4
    port map (
            O => \N__3585\,
            I => \BBn_c\
        );

    \I__534\ : IoInMux
    port map (
            O => \N__3582\,
            I => \N__3579\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3579\,
            I => \N__3576\
        );

    \I__532\ : IoSpan4Mux
    port map (
            O => \N__3576\,
            I => \N__3573\
        );

    \I__531\ : Span4Mux_s2_v
    port map (
            O => \N__3573\,
            I => \N__3570\
        );

    \I__530\ : Span4Mux_v
    port map (
            O => \N__3570\,
            I => \N__3567\
        );

    \I__529\ : Odrv4
    port map (
            O => \N__3567\,
            I => \BUFDIR_c\
        );

    \I__528\ : IoInMux
    port map (
            O => \N__3564\,
            I => \N__3560\
        );

    \I__527\ : IoInMux
    port map (
            O => \N__3563\,
            I => \N__3557\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3560\,
            I => \N__3553\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3557\,
            I => \N__3549\
        );

    \I__524\ : IoInMux
    port map (
            O => \N__3556\,
            I => \N__3546\
        );

    \I__523\ : IoSpan4Mux
    port map (
            O => \N__3553\,
            I => \N__3543\
        );

    \I__522\ : IoInMux
    port map (
            O => \N__3552\,
            I => \N__3540\
        );

    \I__521\ : Span4Mux_s2_h
    port map (
            O => \N__3549\,
            I => \N__3537\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3546\,
            I => \N__3534\
        );

    \I__519\ : IoSpan4Mux
    port map (
            O => \N__3543\,
            I => \N__3529\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3540\,
            I => \N__3529\
        );

    \I__517\ : Span4Mux_h
    port map (
            O => \N__3537\,
            I => \N__3526\
        );

    \I__516\ : Span4Mux_s1_h
    port map (
            O => \N__3534\,
            I => \N__3523\
        );

    \I__515\ : IoSpan4Mux
    port map (
            O => \N__3529\,
            I => \N__3520\
        );

    \I__514\ : Span4Mux_h
    port map (
            O => \N__3526\,
            I => \N__3517\
        );

    \I__513\ : Span4Mux_h
    port map (
            O => \N__3523\,
            I => \N__3514\
        );

    \I__512\ : Span4Mux_s3_v
    port map (
            O => \N__3520\,
            I => \N__3511\
        );

    \I__511\ : Span4Mux_h
    port map (
            O => \N__3517\,
            I => \N__3508\
        );

    \I__510\ : Span4Mux_h
    port map (
            O => \N__3514\,
            I => \N__3505\
        );

    \I__509\ : Sp12to4
    port map (
            O => \N__3511\,
            I => \N__3502\
        );

    \I__508\ : Span4Mux_h
    port map (
            O => \N__3508\,
            I => \N__3497\
        );

    \I__507\ : Span4Mux_h
    port map (
            O => \N__3505\,
            I => \N__3497\
        );

    \I__506\ : Odrv12
    port map (
            O => \N__3502\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__505\ : Odrv4
    port map (
            O => \N__3497\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__504\ : CascadeMux
    port map (
            O => \N__3492\,
            I => \N__3489\
        );

    \I__503\ : InMux
    port map (
            O => \N__3489\,
            I => \N__3486\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3486\,
            I => \N__3483\
        );

    \I__501\ : Span4Mux_v
    port map (
            O => \N__3483\,
            I => \N__3480\
        );

    \I__500\ : Odrv4
    port map (
            O => \N__3480\,
            I => \U111_CYCLE_SM.N_141\
        );

    \I__499\ : InMux
    port map (
            O => \N__3477\,
            I => \N__3474\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3474\,
            I => \N__3471\
        );

    \I__497\ : Span4Mux_v
    port map (
            O => \N__3471\,
            I => \N__3468\
        );

    \I__496\ : Span4Mux_v
    port map (
            O => \N__3468\,
            I => \N__3464\
        );

    \I__495\ : InMux
    port map (
            O => \N__3467\,
            I => \N__3461\
        );

    \I__494\ : Sp12to4
    port map (
            O => \N__3464\,
            I => \N__3456\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3461\,
            I => \N__3456\
        );

    \I__492\ : Span12Mux_h
    port map (
            O => \N__3456\,
            I => \N__3453\
        );

    \I__491\ : Odrv12
    port map (
            O => \N__3453\,
            I => \A_040_c_1\
        );

    \I__490\ : InMux
    port map (
            O => \N__3450\,
            I => \N__3447\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3447\,
            I => \N__3444\
        );

    \I__488\ : Span12Mux_v
    port map (
            O => \N__3444\,
            I => \N__3441\
        );

    \I__487\ : Odrv12
    port map (
            O => \N__3441\,
            I => \D_LM_AMIGA_in_5\
        );

    \I__486\ : IoInMux
    port map (
            O => \N__3438\,
            I => \N__3435\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3435\,
            I => \N__3432\
        );

    \I__484\ : Span12Mux_s8_h
    port map (
            O => \N__3432\,
            I => \N__3429\
        );

    \I__483\ : Span12Mux_h
    port map (
            O => \N__3429\,
            I => \N__3426\
        );

    \I__482\ : Odrv12
    port map (
            O => \N__3426\,
            I => \N_108\
        );

    \I__481\ : InMux
    port map (
            O => \N__3423\,
            I => \N__3420\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3420\,
            I => \N__3417\
        );

    \I__479\ : Span12Mux_h
    port map (
            O => \N__3417\,
            I => \N__3414\
        );

    \I__478\ : Odrv12
    port map (
            O => \N__3414\,
            I => \D_LM_AMIGA_in_3\
        );

    \I__477\ : IoInMux
    port map (
            O => \N__3411\,
            I => \N__3408\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3408\,
            I => \N__3405\
        );

    \I__475\ : IoSpan4Mux
    port map (
            O => \N__3405\,
            I => \N__3402\
        );

    \I__474\ : Span4Mux_s1_h
    port map (
            O => \N__3402\,
            I => \N__3399\
        );

    \I__473\ : Span4Mux_v
    port map (
            O => \N__3399\,
            I => \N__3396\
        );

    \I__472\ : Sp12to4
    port map (
            O => \N__3396\,
            I => \N__3393\
        );

    \I__471\ : Span12Mux_s10_h
    port map (
            O => \N__3393\,
            I => \N__3390\
        );

    \I__470\ : Odrv12
    port map (
            O => \N__3390\,
            I => \N_110\
        );

    \I__469\ : InMux
    port map (
            O => \N__3387\,
            I => \N__3384\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__3384\,
            I => \N__3381\
        );

    \I__467\ : Span12Mux_h
    port map (
            O => \N__3381\,
            I => \N__3378\
        );

    \I__466\ : Odrv12
    port map (
            O => \N__3378\,
            I => \D_LM_AMIGA_in_2\
        );

    \I__465\ : IoInMux
    port map (
            O => \N__3375\,
            I => \N__3372\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3372\,
            I => \N__3369\
        );

    \I__463\ : Span12Mux_s3_h
    port map (
            O => \N__3369\,
            I => \N__3366\
        );

    \I__462\ : Span12Mux_h
    port map (
            O => \N__3366\,
            I => \N__3363\
        );

    \I__461\ : Span12Mux_v
    port map (
            O => \N__3363\,
            I => \N__3360\
        );

    \I__460\ : Odrv12
    port map (
            O => \N__3360\,
            I => \N_111\
        );

    \I__459\ : InMux
    port map (
            O => \N__3357\,
            I => \N__3354\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3354\,
            I => \N__3351\
        );

    \I__457\ : Span4Mux_v
    port map (
            O => \N__3351\,
            I => \N__3348\
        );

    \I__456\ : Sp12to4
    port map (
            O => \N__3348\,
            I => \N__3345\
        );

    \I__455\ : Span12Mux_h
    port map (
            O => \N__3345\,
            I => \N__3342\
        );

    \I__454\ : Odrv12
    port map (
            O => \N__3342\,
            I => \D_UM_040_in_6\
        );

    \I__453\ : IoInMux
    port map (
            O => \N__3339\,
            I => \N__3336\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3336\,
            I => \N__3333\
        );

    \I__451\ : IoSpan4Mux
    port map (
            O => \N__3333\,
            I => \N__3329\
        );

    \I__450\ : InMux
    port map (
            O => \N__3332\,
            I => \N__3326\
        );

    \I__449\ : IoSpan4Mux
    port map (
            O => \N__3329\,
            I => \N__3323\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3326\,
            I => \N__3320\
        );

    \I__447\ : Span4Mux_s2_h
    port map (
            O => \N__3323\,
            I => \N__3317\
        );

    \I__446\ : Span4Mux_v
    port map (
            O => \N__3320\,
            I => \N__3314\
        );

    \I__445\ : Sp12to4
    port map (
            O => \N__3317\,
            I => \N__3311\
        );

    \I__444\ : Sp12to4
    port map (
            O => \N__3314\,
            I => \N__3308\
        );

    \I__443\ : Span12Mux_h
    port map (
            O => \N__3311\,
            I => \N__3305\
        );

    \I__442\ : Span12Mux_h
    port map (
            O => \N__3308\,
            I => \N__3302\
        );

    \I__441\ : Span12Mux_h
    port map (
            O => \N__3305\,
            I => \N__3297\
        );

    \I__440\ : Span12Mux_v
    port map (
            O => \N__3302\,
            I => \N__3297\
        );

    \I__439\ : Odrv12
    port map (
            O => \N__3297\,
            I => \D_LL_040_in_6\
        );

    \I__438\ : IoInMux
    port map (
            O => \N__3294\,
            I => \N__3291\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__3291\,
            I => \N__3288\
        );

    \I__436\ : Span12Mux_s9_h
    port map (
            O => \N__3288\,
            I => \N__3285\
        );

    \I__435\ : Span12Mux_v
    port map (
            O => \N__3285\,
            I => \N__3282\
        );

    \I__434\ : Odrv12
    port map (
            O => \N__3282\,
            I => \un1_D_UM_040_6\
        );

    \I__433\ : InMux
    port map (
            O => \N__3279\,
            I => \N__3276\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__3276\,
            I => \N__3273\
        );

    \I__431\ : Span4Mux_v
    port map (
            O => \N__3273\,
            I => \N__3270\
        );

    \I__430\ : Span4Mux_h
    port map (
            O => \N__3270\,
            I => \N__3267\
        );

    \I__429\ : Sp12to4
    port map (
            O => \N__3267\,
            I => \N__3264\
        );

    \I__428\ : Span12Mux_h
    port map (
            O => \N__3264\,
            I => \N__3261\
        );

    \I__427\ : Odrv12
    port map (
            O => \N__3261\,
            I => \D_UU_040_in_0\
        );

    \I__426\ : IoInMux
    port map (
            O => \N__3258\,
            I => \N__3254\
        );

    \I__425\ : InMux
    port map (
            O => \N__3257\,
            I => \N__3251\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3254\,
            I => \N__3248\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__3251\,
            I => \N__3245\
        );

    \I__422\ : IoSpan4Mux
    port map (
            O => \N__3248\,
            I => \N__3242\
        );

    \I__421\ : Span4Mux_v
    port map (
            O => \N__3245\,
            I => \N__3239\
        );

    \I__420\ : Span4Mux_s2_h
    port map (
            O => \N__3242\,
            I => \N__3236\
        );

    \I__419\ : Sp12to4
    port map (
            O => \N__3239\,
            I => \N__3233\
        );

    \I__418\ : Span4Mux_v
    port map (
            O => \N__3236\,
            I => \N__3230\
        );

    \I__417\ : Span12Mux_h
    port map (
            O => \N__3233\,
            I => \N__3227\
        );

    \I__416\ : Sp12to4
    port map (
            O => \N__3230\,
            I => \N__3224\
        );

    \I__415\ : Span12Mux_v
    port map (
            O => \N__3227\,
            I => \N__3221\
        );

    \I__414\ : Span12Mux_s9_h
    port map (
            O => \N__3224\,
            I => \N__3218\
        );

    \I__413\ : Span12Mux_v
    port map (
            O => \N__3221\,
            I => \N__3213\
        );

    \I__412\ : Span12Mux_h
    port map (
            O => \N__3218\,
            I => \N__3213\
        );

    \I__411\ : Odrv12
    port map (
            O => \N__3213\,
            I => \D_LM_040_in_0\
        );

    \I__410\ : IoInMux
    port map (
            O => \N__3210\,
            I => \N__3207\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3207\,
            I => \N__3204\
        );

    \I__408\ : IoSpan4Mux
    port map (
            O => \N__3204\,
            I => \N__3201\
        );

    \I__407\ : Span4Mux_s2_v
    port map (
            O => \N__3201\,
            I => \N__3198\
        );

    \I__406\ : Span4Mux_v
    port map (
            O => \N__3198\,
            I => \N__3195\
        );

    \I__405\ : Odrv4
    port map (
            O => \N__3195\,
            I => \un1_D_UU_040_0\
        );

    \I__404\ : InMux
    port map (
            O => \N__3192\,
            I => \N__3189\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__3189\,
            I => \N__3186\
        );

    \I__402\ : Span4Mux_v
    port map (
            O => \N__3186\,
            I => \N__3183\
        );

    \I__401\ : Span4Mux_h
    port map (
            O => \N__3183\,
            I => \N__3180\
        );

    \I__400\ : Sp12to4
    port map (
            O => \N__3180\,
            I => \N__3177\
        );

    \I__399\ : Span12Mux_h
    port map (
            O => \N__3177\,
            I => \N__3174\
        );

    \I__398\ : Odrv12
    port map (
            O => \N__3174\,
            I => \D_UU_040_in_6\
        );

    \I__397\ : IoInMux
    port map (
            O => \N__3171\,
            I => \N__3168\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3168\,
            I => \N__3164\
        );

    \I__395\ : InMux
    port map (
            O => \N__3167\,
            I => \N__3161\
        );

    \I__394\ : Span4Mux_s2_h
    port map (
            O => \N__3164\,
            I => \N__3158\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3161\,
            I => \N__3155\
        );

    \I__392\ : Span4Mux_v
    port map (
            O => \N__3158\,
            I => \N__3152\
        );

    \I__391\ : Span4Mux_v
    port map (
            O => \N__3155\,
            I => \N__3149\
        );

    \I__390\ : Sp12to4
    port map (
            O => \N__3152\,
            I => \N__3146\
        );

    \I__389\ : Span4Mux_v
    port map (
            O => \N__3149\,
            I => \N__3143\
        );

    \I__388\ : Span12Mux_h
    port map (
            O => \N__3146\,
            I => \N__3138\
        );

    \I__387\ : Sp12to4
    port map (
            O => \N__3143\,
            I => \N__3138\
        );

    \I__386\ : Span12Mux_h
    port map (
            O => \N__3138\,
            I => \N__3135\
        );

    \I__385\ : Odrv12
    port map (
            O => \N__3135\,
            I => \D_LM_040_in_6\
        );

    \I__384\ : IoInMux
    port map (
            O => \N__3132\,
            I => \N__3129\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3129\,
            I => \N__3126\
        );

    \I__382\ : Span4Mux_s3_v
    port map (
            O => \N__3126\,
            I => \N__3123\
        );

    \I__381\ : Span4Mux_h
    port map (
            O => \N__3123\,
            I => \N__3120\
        );

    \I__380\ : Span4Mux_h
    port map (
            O => \N__3120\,
            I => \N__3117\
        );

    \I__379\ : Odrv4
    port map (
            O => \N__3117\,
            I => \un1_D_UU_040_6\
        );

    \I__378\ : InMux
    port map (
            O => \N__3114\,
            I => \N__3111\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__3111\,
            I => \N__3108\
        );

    \I__376\ : Span4Mux_v
    port map (
            O => \N__3108\,
            I => \N__3105\
        );

    \I__375\ : Sp12to4
    port map (
            O => \N__3105\,
            I => \N__3102\
        );

    \I__374\ : Odrv12
    port map (
            O => \N__3102\,
            I => \D_LL_AMIGA_in_4\
        );

    \I__373\ : IoInMux
    port map (
            O => \N__3099\,
            I => \N__3096\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3096\,
            I => \N__3093\
        );

    \I__371\ : Span4Mux_s2_h
    port map (
            O => \N__3093\,
            I => \N__3090\
        );

    \I__370\ : Sp12to4
    port map (
            O => \N__3090\,
            I => \N__3087\
        );

    \I__369\ : Span12Mux_s8_v
    port map (
            O => \N__3087\,
            I => \N__3084\
        );

    \I__368\ : Span12Mux_h
    port map (
            O => \N__3084\,
            I => \N__3081\
        );

    \I__367\ : Odrv12
    port map (
            O => \N__3081\,
            I => \un2_D_LL_AMIGA_4\
        );

    \I__366\ : IoInMux
    port map (
            O => \N__3078\,
            I => \N__3075\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__3075\,
            I => \N__3072\
        );

    \I__364\ : Odrv12
    port map (
            O => \N__3072\,
            I => \U111_CYCLE_SM_A_AMIGA_0_i_1\
        );

    \I__363\ : InMux
    port map (
            O => \N__3069\,
            I => \N__3066\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__3066\,
            I => \N__3063\
        );

    \I__361\ : Span4Mux_h
    port map (
            O => \N__3063\,
            I => \N__3060\
        );

    \I__360\ : Span4Mux_v
    port map (
            O => \N__3060\,
            I => \N__3057\
        );

    \I__359\ : Odrv4
    port map (
            O => \N__3057\,
            I => \A_040_c_0\
        );

    \I__358\ : IoInMux
    port map (
            O => \N__3054\,
            I => \N__3051\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__3051\,
            I => \N__3048\
        );

    \I__356\ : Span12Mux_s6_v
    port map (
            O => \N__3048\,
            I => \N__3045\
        );

    \I__355\ : Odrv12
    port map (
            O => \N__3045\,
            I => \A_AMIGA_c_0\
        );

    \I__354\ : InMux
    port map (
            O => \N__3042\,
            I => \N__3039\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__3039\,
            I => \N__3036\
        );

    \I__352\ : Span12Mux_h
    port map (
            O => \N__3036\,
            I => \N__3033\
        );

    \I__351\ : Span12Mux_h
    port map (
            O => \N__3033\,
            I => \N__3030\
        );

    \I__350\ : Odrv12
    port map (
            O => \N__3030\,
            I => \D_UM_040_in_2\
        );

    \I__349\ : IoInMux
    port map (
            O => \N__3027\,
            I => \N__3023\
        );

    \I__348\ : InMux
    port map (
            O => \N__3026\,
            I => \N__3020\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__3023\,
            I => \N__3017\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__3020\,
            I => \N__3014\
        );

    \I__345\ : IoSpan4Mux
    port map (
            O => \N__3017\,
            I => \N__3011\
        );

    \I__344\ : Span4Mux_v
    port map (
            O => \N__3014\,
            I => \N__3008\
        );

    \I__343\ : Span4Mux_s2_h
    port map (
            O => \N__3011\,
            I => \N__3005\
        );

    \I__342\ : Sp12to4
    port map (
            O => \N__3008\,
            I => \N__3002\
        );

    \I__341\ : Sp12to4
    port map (
            O => \N__3005\,
            I => \N__2999\
        );

    \I__340\ : Span12Mux_h
    port map (
            O => \N__3002\,
            I => \N__2996\
        );

    \I__339\ : Span12Mux_h
    port map (
            O => \N__2999\,
            I => \N__2993\
        );

    \I__338\ : Span12Mux_v
    port map (
            O => \N__2996\,
            I => \N__2990\
        );

    \I__337\ : Span12Mux_h
    port map (
            O => \N__2993\,
            I => \N__2987\
        );

    \I__336\ : Odrv12
    port map (
            O => \N__2990\,
            I => \D_LL_040_in_2\
        );

    \I__335\ : Odrv12
    port map (
            O => \N__2987\,
            I => \D_LL_040_in_2\
        );

    \I__334\ : IoInMux
    port map (
            O => \N__2982\,
            I => \N__2979\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2979\,
            I => \N__2976\
        );

    \I__332\ : Span4Mux_s3_h
    port map (
            O => \N__2976\,
            I => \N__2973\
        );

    \I__331\ : Span4Mux_h
    port map (
            O => \N__2973\,
            I => \N__2970\
        );

    \I__330\ : Span4Mux_v
    port map (
            O => \N__2970\,
            I => \N__2967\
        );

    \I__329\ : Odrv4
    port map (
            O => \N__2967\,
            I => \un1_D_UM_040_2\
        );

    \I__328\ : InMux
    port map (
            O => \N__2964\,
            I => \N__2961\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2961\,
            I => \N__2958\
        );

    \I__326\ : Span4Mux_h
    port map (
            O => \N__2958\,
            I => \N__2955\
        );

    \I__325\ : Span4Mux_v
    port map (
            O => \N__2955\,
            I => \N__2952\
        );

    \I__324\ : Span4Mux_h
    port map (
            O => \N__2952\,
            I => \N__2949\
        );

    \I__323\ : Span4Mux_h
    port map (
            O => \N__2949\,
            I => \N__2946\
        );

    \I__322\ : Span4Mux_h
    port map (
            O => \N__2946\,
            I => \N__2943\
        );

    \I__321\ : Odrv4
    port map (
            O => \N__2943\,
            I => \D_UU_040_in_4\
        );

    \I__320\ : IoInMux
    port map (
            O => \N__2940\,
            I => \N__2937\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2937\,
            I => \N__2934\
        );

    \I__318\ : Span4Mux_s1_h
    port map (
            O => \N__2934\,
            I => \N__2931\
        );

    \I__317\ : Span4Mux_h
    port map (
            O => \N__2931\,
            I => \N__2927\
        );

    \I__316\ : InMux
    port map (
            O => \N__2930\,
            I => \N__2924\
        );

    \I__315\ : Sp12to4
    port map (
            O => \N__2927\,
            I => \N__2921\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2924\,
            I => \N__2918\
        );

    \I__313\ : Span12Mux_v
    port map (
            O => \N__2921\,
            I => \N__2915\
        );

    \I__312\ : Span12Mux_h
    port map (
            O => \N__2918\,
            I => \N__2912\
        );

    \I__311\ : Span12Mux_h
    port map (
            O => \N__2915\,
            I => \N__2907\
        );

    \I__310\ : Span12Mux_v
    port map (
            O => \N__2912\,
            I => \N__2907\
        );

    \I__309\ : Span12Mux_h
    port map (
            O => \N__2907\,
            I => \N__2904\
        );

    \I__308\ : Odrv12
    port map (
            O => \N__2904\,
            I => \D_LM_040_in_4\
        );

    \I__307\ : IoInMux
    port map (
            O => \N__2901\,
            I => \N__2898\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2898\,
            I => \N__2895\
        );

    \I__305\ : Span4Mux_s3_v
    port map (
            O => \N__2895\,
            I => \N__2892\
        );

    \I__304\ : Span4Mux_h
    port map (
            O => \N__2892\,
            I => \N__2889\
        );

    \I__303\ : Odrv4
    port map (
            O => \N__2889\,
            I => \un1_D_UU_040_4\
        );

    \I__302\ : InMux
    port map (
            O => \N__2886\,
            I => \N__2883\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2883\,
            I => \N__2880\
        );

    \I__300\ : Span4Mux_v
    port map (
            O => \N__2880\,
            I => \N__2877\
        );

    \I__299\ : Sp12to4
    port map (
            O => \N__2877\,
            I => \N__2874\
        );

    \I__298\ : Span12Mux_h
    port map (
            O => \N__2874\,
            I => \N__2871\
        );

    \I__297\ : Span12Mux_h
    port map (
            O => \N__2871\,
            I => \N__2868\
        );

    \I__296\ : Odrv12
    port map (
            O => \N__2868\,
            I => \D_UM_040_in_4\
        );

    \I__295\ : IoInMux
    port map (
            O => \N__2865\,
            I => \N__2862\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2862\,
            I => \N__2858\
        );

    \I__293\ : InMux
    port map (
            O => \N__2861\,
            I => \N__2855\
        );

    \I__292\ : Span4Mux_s2_h
    port map (
            O => \N__2858\,
            I => \N__2852\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2855\,
            I => \N__2849\
        );

    \I__290\ : Span4Mux_v
    port map (
            O => \N__2852\,
            I => \N__2846\
        );

    \I__289\ : Span12Mux_h
    port map (
            O => \N__2849\,
            I => \N__2843\
        );

    \I__288\ : Sp12to4
    port map (
            O => \N__2846\,
            I => \N__2840\
        );

    \I__287\ : Span12Mux_v
    port map (
            O => \N__2843\,
            I => \N__2837\
        );

    \I__286\ : Span12Mux_h
    port map (
            O => \N__2840\,
            I => \N__2834\
        );

    \I__285\ : Span12Mux_v
    port map (
            O => \N__2837\,
            I => \N__2831\
        );

    \I__284\ : Span12Mux_h
    port map (
            O => \N__2834\,
            I => \N__2828\
        );

    \I__283\ : Odrv12
    port map (
            O => \N__2831\,
            I => \D_LL_040_in_4\
        );

    \I__282\ : Odrv12
    port map (
            O => \N__2828\,
            I => \D_LL_040_in_4\
        );

    \I__281\ : IoInMux
    port map (
            O => \N__2823\,
            I => \N__2820\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__2820\,
            I => \N__2817\
        );

    \I__279\ : Span4Mux_s2_h
    port map (
            O => \N__2817\,
            I => \N__2814\
        );

    \I__278\ : Span4Mux_h
    port map (
            O => \N__2814\,
            I => \N__2811\
        );

    \I__277\ : Span4Mux_h
    port map (
            O => \N__2811\,
            I => \N__2808\
        );

    \I__276\ : Odrv4
    port map (
            O => \N__2808\,
            I => \un1_D_UM_040_4\
        );

    \I__275\ : InMux
    port map (
            O => \N__2805\,
            I => \N__2802\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2802\,
            I => \N__2799\
        );

    \I__273\ : Span4Mux_v
    port map (
            O => \N__2799\,
            I => \N__2796\
        );

    \I__272\ : Sp12to4
    port map (
            O => \N__2796\,
            I => \N__2793\
        );

    \I__271\ : Span12Mux_h
    port map (
            O => \N__2793\,
            I => \N__2790\
        );

    \I__270\ : Odrv12
    port map (
            O => \N__2790\,
            I => \D_LL_AMIGA_in_1\
        );

    \I__269\ : IoInMux
    port map (
            O => \N__2787\,
            I => \N__2784\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2784\,
            I => \N__2781\
        );

    \I__267\ : IoSpan4Mux
    port map (
            O => \N__2781\,
            I => \N__2778\
        );

    \I__266\ : Span4Mux_s3_h
    port map (
            O => \N__2778\,
            I => \N__2775\
        );

    \I__265\ : Span4Mux_v
    port map (
            O => \N__2775\,
            I => \N__2772\
        );

    \I__264\ : Span4Mux_h
    port map (
            O => \N__2772\,
            I => \N__2769\
        );

    \I__263\ : Sp12to4
    port map (
            O => \N__2769\,
            I => \N__2766\
        );

    \I__262\ : Odrv12
    port map (
            O => \N__2766\,
            I => \un2_D_LL_AMIGA_1\
        );

    \I__261\ : IoInMux
    port map (
            O => \N__2763\,
            I => \N__2760\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2760\,
            I => \N__2757\
        );

    \I__259\ : Span12Mux_s1_v
    port map (
            O => \N__2757\,
            I => \N__2754\
        );

    \I__258\ : Odrv12
    port map (
            O => \N__2754\,
            I => \CPUBGn_c_i_0\
        );

    \I__257\ : InMux
    port map (
            O => \N__2751\,
            I => \N__2748\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__2748\,
            I => \N__2745\
        );

    \I__255\ : Span4Mux_v
    port map (
            O => \N__2745\,
            I => \N__2742\
        );

    \I__254\ : Sp12to4
    port map (
            O => \N__2742\,
            I => \N__2739\
        );

    \I__253\ : Span12Mux_h
    port map (
            O => \N__2739\,
            I => \N__2736\
        );

    \I__252\ : Odrv12
    port map (
            O => \N__2736\,
            I => \D_LL_AMIGA_in_5\
        );

    \I__251\ : IoInMux
    port map (
            O => \N__2733\,
            I => \N__2730\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2730\,
            I => \N__2727\
        );

    \I__249\ : Span12Mux_s8_h
    port map (
            O => \N__2727\,
            I => \N__2724\
        );

    \I__248\ : Span12Mux_h
    port map (
            O => \N__2724\,
            I => \N__2721\
        );

    \I__247\ : Odrv12
    port map (
            O => \N__2721\,
            I => \un2_D_LL_AMIGA_5\
        );

    \I__246\ : InMux
    port map (
            O => \N__2718\,
            I => \N__2715\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2715\,
            I => \N__2712\
        );

    \I__244\ : Span12Mux_v
    port map (
            O => \N__2712\,
            I => \N__2709\
        );

    \I__243\ : Odrv12
    port map (
            O => \N__2709\,
            I => \D_LL_AMIGA_in_7\
        );

    \I__242\ : IoInMux
    port map (
            O => \N__2706\,
            I => \N__2703\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__2703\,
            I => \N__2700\
        );

    \I__240\ : Span4Mux_s2_h
    port map (
            O => \N__2700\,
            I => \N__2697\
        );

    \I__239\ : Sp12to4
    port map (
            O => \N__2697\,
            I => \N__2694\
        );

    \I__238\ : Span12Mux_v
    port map (
            O => \N__2694\,
            I => \N__2691\
        );

    \I__237\ : Span12Mux_h
    port map (
            O => \N__2691\,
            I => \N__2688\
        );

    \I__236\ : Odrv12
    port map (
            O => \N__2688\,
            I => \un2_D_LL_AMIGA_7\
        );

    \I__235\ : IoInMux
    port map (
            O => \N__2685\,
            I => \N__2682\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2682\,
            I => \N__2679\
        );

    \I__233\ : Span4Mux_s0_v
    port map (
            O => \N__2679\,
            I => \N__2676\
        );

    \I__232\ : Sp12to4
    port map (
            O => \N__2676\,
            I => \N__2673\
        );

    \I__231\ : Span12Mux_h
    port map (
            O => \N__2673\,
            I => \N__2670\
        );

    \I__230\ : Span12Mux_v
    port map (
            O => \N__2670\,
            I => \N__2667\
        );

    \I__229\ : Span12Mux_v
    port map (
            O => \N__2667\,
            I => \N__2664\
        );

    \I__228\ : Odrv12
    port map (
            O => \N__2664\,
            I => \TAn_in\
        );

    \I__227\ : IoInMux
    port map (
            O => \N__2661\,
            I => \N__2658\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__2658\,
            I => \N__2655\
        );

    \I__225\ : Odrv12
    port map (
            O => \N__2655\,
            I => \RESETn_c_i\
        );

    \INVU111_CYCLE_SM.TS_OUTC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TS_OUTC_net\,
            I => \N__7133\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2661\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6214\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__3467\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3813\,
            lcout => \U111_CYCLE_SM_A_AMIGA_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__3069\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3812\,
            lcout => \A_AMIGA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8134\,
            in1 => \N__3042\,
            in2 => \_gnd_net_\,
            in3 => \N__3026\,
            lcout => \un1_D_UM_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8214\,
            in1 => \N__2964\,
            in2 => \_gnd_net_\,
            in3 => \N__2930\,
            lcout => \un1_D_UU_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2886\,
            in1 => \N__2861\,
            in2 => \_gnd_net_\,
            in3 => \N__8213\,
            lcout => \un1_D_UM_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7014\,
            in1 => \N__2805\,
            in2 => \_gnd_net_\,
            in3 => \N__8174\,
            lcout => \un2_D_LL_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TSn_obuft_RNO_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7791\,
            lcout => \CPUBGn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2751\,
            in1 => \N__7952\,
            in2 => \_gnd_net_\,
            in3 => \N__8130\,
            lcout => \un2_D_LL_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2718\,
            in1 => \N__8426\,
            in2 => \_gnd_net_\,
            in3 => \N__8129\,
            lcout => \un2_D_LL_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4142\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3477\,
            lcout => \U111_CYCLE_SM.N_141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3450\,
            in1 => \N__4322\,
            in2 => \_gnd_net_\,
            in3 => \N__8136\,
            lcout => \N_108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3423\,
            in1 => \N__6728\,
            in2 => \_gnd_net_\,
            in3 => \N__8135\,
            lcout => \N_110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3387\,
            in1 => \N__4656\,
            in2 => \_gnd_net_\,
            in3 => \N__8137\,
            lcout => \N_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8138\,
            in1 => \N__3357\,
            in2 => \_gnd_net_\,
            in3 => \N__3332\,
            lcout => \un1_D_UM_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8211\,
            in1 => \N__3279\,
            in2 => \_gnd_net_\,
            in3 => \N__3257\,
            lcout => \un1_D_UU_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8212\,
            in1 => \N__3192\,
            in2 => \_gnd_net_\,
            in3 => \N__3167\,
            lcout => \un1_D_UU_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8168\,
            in1 => \N__5942\,
            in2 => \_gnd_net_\,
            in3 => \N__3114\,
            lcout => \un2_D_LL_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3786\,
            in1 => \N__6411\,
            in2 => \_gnd_net_\,
            in3 => \N__8167\,
            lcout => \un2_D_LL_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3749\,
            in1 => \N__3714\,
            in2 => \_gnd_net_\,
            in3 => \N__8025\,
            lcout => \un1_D_UM_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8026\,
            in1 => \N__6038\,
            in2 => \_gnd_net_\,
            in3 => \N__3675\,
            lcout => \N_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_BUFFERS.DMA_EN_i_0_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__3604\,
            in1 => \N__7805\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_BUFFERS.N_94_i_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__7806\,
            in1 => \N__3605\,
            in2 => \_gnd_net_\,
            in3 => \N__6875\,
            lcout => \N_94_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_BUFFERS.un1_DMA_EN_0_0_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101010"
        )
    port map (
            in0 => \N__7725\,
            in1 => \N__3606\,
            in2 => \_gnd_net_\,
            in3 => \N__7807\,
            lcout => \BUFDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_THRU_LUT4_0_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7143\,
            lcout => \GB_BUFFER_CLK40_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000110010"
        )
    port map (
            in0 => \N__4122\,
            in1 => \N__4086\,
            in2 => \N__5100\,
            in3 => \N__4065\,
            lcout => \U111_CYCLE_SM.TS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7135\,
            ce => 'H',
            sr => \N__6294\
        );

    \U111_CYCLE_SM.FLIP_WORD_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__5096\,
            in1 => \N__8024\,
            in2 => \N__3492\,
            in3 => \N__4177\,
            lcout => \U111_CYCLE_SM.FLIP_WORDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7135\,
            ce => 'H',
            sr => \N__6294\
        );

    \U111_CYCLE_SM.TS_OUT_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101010111"
        )
    port map (
            in0 => \N__6263\,
            in1 => \N__4064\,
            in2 => \N__6876\,
            in3 => \N__5220\,
            lcout => \TS_OUT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TS_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8149\,
            in1 => \N__4493\,
            in2 => \_gnd_net_\,
            in3 => \N__4053\,
            lcout => \N_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4014\,
            in1 => \N__5613\,
            in2 => \_gnd_net_\,
            in3 => \N__8148\,
            lcout => \N_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3981\,
            in1 => \N__3966\,
            in2 => \_gnd_net_\,
            in3 => \N__8186\,
            lcout => \un1_D_UM_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3903\,
            in1 => \N__8206\,
            in2 => \_gnd_net_\,
            in3 => \N__8616\,
            lcout => \un2_D_LL_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LBENn_c_sbtinv_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6835\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \LBENn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8067\,
            in1 => \N__5811\,
            in2 => \_gnd_net_\,
            in3 => \N__3852\,
            lcout => \un2_D_LM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.un1_CYCLE_STATE_1_i_i_o2_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__6484\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5154\,
            lcout => \U111_CYCLE_SM.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__3797\,
            in1 => \N__5093\,
            in2 => \N__4105\,
            in3 => \N__4851\,
            lcout => \U111_CYCLE_SM.A2_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7136\,
            ce => 'H',
            sr => \N__6297\
        );

    \U111_CYCLE_SM.BURST_RNILNBJ_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4870\,
            in2 => \_gnd_net_\,
            in3 => \N__4848\,
            lcout => \U111_CYCLE_SM.N_179\,
            ltout => \U111_CYCLE_SM.N_179_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001000000"
        )
    port map (
            in0 => \N__4106\,
            in1 => \N__6252\,
            in2 => \N__4116\,
            in3 => \N__5051\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7134\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__4154\,
            in1 => \N__4192\,
            in2 => \_gnd_net_\,
            in3 => \N__4175\,
            lcout => \U111_CYCLE_SM.N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101110111"
        )
    port map (
            in0 => \N__4869\,
            in1 => \N__6618\,
            in2 => \N__4215\,
            in3 => \N__4277\,
            lcout => \U111_CYCLE_SM.N_101\,
            ltout => \U111_CYCLE_SM.N_101_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5158\,
            in1 => \N__4890\,
            in2 => \N__4113\,
            in3 => \N__5127\,
            lcout => \U111_CYCLE_SM.N_133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__5128\,
            in1 => \N__4849\,
            in2 => \N__4110\,
            in3 => \N__6335\,
            lcout => \U111_CYCLE_SM.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011101"
        )
    port map (
            in0 => \N__6498\,
            in1 => \N__4080\,
            in2 => \N__5162\,
            in3 => \N__4891\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_12_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_2_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000000000"
        )
    port map (
            in0 => \N__4176\,
            in1 => \N__5130\,
            in2 => \N__4074\,
            in3 => \N__6253\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7134\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_DIS_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000011111110"
        )
    port map (
            in0 => \N__5094\,
            in1 => \N__4179\,
            in2 => \N__6940\,
            in3 => \N__4071\,
            lcout => \U111_CYCLE_SM.TA_DISZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7129\,
            ce => 'H',
            sr => \N__6293\
        );

    \U111_CYCLE_SM.BURST_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__5048\,
            in1 => \N__4265\,
            in2 => \N__4242\,
            in3 => \N__4872\,
            lcout => \U111_CYCLE_SM.BURSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7129\,
            ce => 'H',
            sr => \N__6293\
        );

    \U111_CYCLE_SM.BURST_COUNT_1_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100100001100"
        )
    port map (
            in0 => \N__6185\,
            in1 => \N__4278\,
            in2 => \N__5052\,
            in3 => \N__4214\,
            lcout => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7129\,
            ce => 'H',
            sr => \N__6293\
        );

    \U111_CYCLE_SM.LW_TRANS_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__4266\,
            in1 => \N__4241\,
            in2 => \N__4197\,
            in3 => \N__5049\,
            lcout => \U111_CYCLE_SM.LW_TRANSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7129\,
            ce => 'H',
            sr => \N__6293\
        );

    \U111_CYCLE_SM.BURST_COUNT_0_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__5043\,
            in1 => \N__6184\,
            in2 => \_gnd_net_\,
            in3 => \N__4213\,
            lcout => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7129\,
            ce => 'H',
            sr => \N__6293\
        );

    \U111_CYCLE_SM.PORT_MISMATCH_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__4193\,
            in1 => \N__4178\,
            in2 => \N__4896\,
            in3 => \N__4155\,
            lcout => \U111_CYCLE_SM.PORT_MISMATCHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7129\,
            ce => 'H',
            sr => \N__6293\
        );

    \U111_CYCLE_SM.CYCLE_EN_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__5044\,
            in1 => \N__5503\,
            in2 => \_gnd_net_\,
            in3 => \N__6337\,
            lcout => \U111_CYCLE_SM.CYCLE_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7129\,
            ce => 'H',
            sr => \N__6293\
        );

    \U111_CYCLE_SM.UU_LATCHED_5_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7882\,
            in1 => \N__4937\,
            in2 => \N__4329\,
            in3 => \N__6157\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7125\,
            ce => 'H',
            sr => \N__6295\
        );

    \U111_CYCLE_SM.UU_LATCHED_2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7880\,
            in1 => \N__4601\,
            in2 => \N__4652\,
            in3 => \N__6155\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7125\,
            ce => 'H',
            sr => \N__6295\
        );

    \U111_CYCLE_SM.UU_LATCHED_7_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7883\,
            in1 => \N__4445\,
            in2 => \N__4494\,
            in3 => \N__6158\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7125\,
            ce => 'H',
            sr => \N__6295\
        );

    \U111_CYCLE_SM.TS_DELAY_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4800\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.TS_DELAYZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7125\,
            ce => 'H',
            sr => \N__6295\
        );

    \U111_CYCLE_SM.UU_LATCHED_4_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__6156\,
            in1 => \N__4568\,
            in2 => \N__4557\,
            in3 => \N__7881\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7125\,
            ce => 'H',
            sr => \N__6295\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4782\,
            in1 => \N__4550\,
            in2 => \_gnd_net_\,
            in3 => \N__8139\,
            lcout => \N_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8208\,
            in1 => \N__4743\,
            in2 => \_gnd_net_\,
            in3 => \N__4724\,
            lcout => \un1_D_UU_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNINJKT_2_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7340\,
            in1 => \N__4648\,
            in2 => \_gnd_net_\,
            in3 => \N__4605\,
            lcout => \N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNIRNKT_4_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4575\,
            in1 => \N__4538\,
            in2 => \_gnd_net_\,
            in3 => \N__7341\,
            lcout => \N_116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNI1UKT_7_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7339\,
            in1 => \N__4486\,
            in2 => \_gnd_net_\,
            in3 => \N__4452\,
            lcout => \N_113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4406\,
            in1 => \N__4365\,
            in2 => \_gnd_net_\,
            in3 => \N__8209\,
            lcout => \un1_D_UU_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNITPKT_5_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7342\,
            in1 => \N__4309\,
            in2 => \_gnd_net_\,
            in3 => \N__4947\,
            lcout => \N_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6491\,
            in2 => \_gnd_net_\,
            in3 => \N__5181\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_i_o2_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__6255\,
            in1 => \N__4902\,
            in2 => \N__4905\,
            in3 => \N__4850\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7132\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6254\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5084\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7132\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6269\,
            in1 => \N__4892\,
            in2 => \_gnd_net_\,
            in3 => \N__6186\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__6502\,
            in1 => \N__4846\,
            in2 => \_gnd_net_\,
            in3 => \N__5129\,
            lcout => \U111_CYCLE_SM.N_131\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5182\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4871\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_a3_2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110011"
        )
    port map (
            in0 => \N__4847\,
            in1 => \N__6270\,
            in2 => \N__4818\,
            in3 => \N__4815\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__6361\,
            in1 => \N__4809\,
            in2 => \N__4803\,
            in3 => \N__6336\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_DELAY_RNIDR7G_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__6839\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5219\,
            lcout => \U111_CYCLE_SM.un4_TS_OUT_i_0\,
            ltout => \U111_CYCLE_SM.un4_TS_OUT_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNI9UTM_0_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5208\,
            in3 => \N__6334\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__5189\,
            in1 => \N__6503\,
            in2 => \_gnd_net_\,
            in3 => \N__5126\,
            lcout => \U111_CYCLE_SM.N_99\,
            ltout => \U111_CYCLE_SM.N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_0_2_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5103\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.N_99_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6333\,
            in2 => \_gnd_net_\,
            in3 => \N__7863\,
            lcout => \U111_CYCLE_SM.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LATCH_EN_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101110010"
        )
    port map (
            in0 => \N__5095\,
            in1 => \N__5058\,
            in2 => \N__7280\,
            in3 => \N__5050\,
            lcout => \U111_CYCLE_SM.LATCH_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7123\,
            ce => 'H',
            sr => \N__6298\
        );

    \U111_CYCLE_SM.CYCLE_EN_RNI26B3_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__5538\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5504\,
            lcout => \CPUBGn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000101110"
        )
    port map (
            in0 => \N__5486\,
            in1 => \N__6344\,
            in2 => \N__7720\,
            in3 => \N__6366\,
            lcout => \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7122\,
            ce => 'H',
            sr => \N__6299\
        );

    \U111_CYCLE_SM.UU_LATCHED_6_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__5624\,
            in1 => \N__7876\,
            in2 => \N__5609\,
            in3 => \N__6159\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7122\,
            ce => 'H',
            sr => \N__6299\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5012\,
            in1 => \N__4983\,
            in2 => \_gnd_net_\,
            in3 => \N__8207\,
            lcout => \un1_D_UU_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TS_CPUn_iobuf_RNO_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7775\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5753\,
            lcout => \TSnz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5699\,
            in1 => \N__5664\,
            in2 => \_gnd_net_\,
            in3 => \N__8210\,
            lcout => \un1_D_UU_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNIVRKT_6_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5631\,
            in1 => \N__5602\,
            in2 => \_gnd_net_\,
            in3 => \N__7309\,
            lcout => \N_114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_1_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__5987\,
            in1 => \N__7865\,
            in2 => \N__6039\,
            in3 => \N__6150\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7130\,
            ce => 'H',
            sr => \N__6296\
        );

    \U111_CYCLE_SM.UU_LATCHED_3_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__6743\,
            in1 => \N__7866\,
            in2 => \N__6732\,
            in3 => \N__6151\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7130\,
            ce => 'H',
            sr => \N__6296\
        );

    \U111_CYCLE_SM.UU_LATCHED_0_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__5822\,
            in1 => \N__7864\,
            in2 => \N__5810\,
            in3 => \N__6149\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7130\,
            ce => 'H',
            sr => \N__6296\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNINRNR_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__7719\,
            in1 => \N__5537\,
            in2 => \N__5514\,
            in3 => \N__5487\,
            lcout => \U111_CYCLE_SM_OFFBOARD_EN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__7862\,
            in1 => \N__6365\,
            in2 => \N__7724\,
            in3 => \N__6345\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7126\,
            ce => 'H',
            sr => \N__6300\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__6262\,
            in1 => \N__7861\,
            in2 => \_gnd_net_\,
            in3 => \N__6183\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\,
            ltout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI0BVS1_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6162\,
            in3 => \N__6148\,
            lcout => \U111_CYCLE_SM.N_99_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5943\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7124\,
            ce => \N__7085\,
            sr => \N__7039\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6117\,
            in1 => \N__6098\,
            in2 => \_gnd_net_\,
            in3 => \N__8197\,
            lcout => \un1_D_UM_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNILHKT_1_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7343\,
            in1 => \N__6028\,
            in2 => \_gnd_net_\,
            in3 => \N__5991\,
            lcout => \N_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7333\,
            in1 => \N__5955\,
            in2 => \_gnd_net_\,
            in3 => \N__5932\,
            lcout => \un1_D_UM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5868\,
            lcout => \GB_BUFFER_CLK80_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNIJFKT_0_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5829\,
            in1 => \N__5797\,
            in2 => \_gnd_net_\,
            in3 => \N__7348\,
            lcout => \un1_D_UU_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNIPLKT_3_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6747\,
            in1 => \N__6718\,
            in2 => \_gnd_net_\,
            in3 => \N__7349\,
            lcout => \N_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_14_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6654\,
            in1 => \N__7185\,
            in2 => \_gnd_net_\,
            in3 => \N__8173\,
            lcout => \un2_D_LL_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TBI_CPUn_0_i_LC_14_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__6608\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6849\,
            lcout => \U111_CYCLE_SM_TBI_CPUn_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6576\,
            in1 => \N__7221\,
            in2 => \_gnd_net_\,
            in3 => \N__8172\,
            lcout => \un2_D_LL_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7320\,
            in1 => \N__6372\,
            in2 => \_gnd_net_\,
            in3 => \N__6401\,
            lcout => \un1_D_UM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7178\,
            in1 => \N__7149\,
            in2 => \_gnd_net_\,
            in3 => \N__7319\,
            lcout => \un1_D_UM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_DIS_RNI576J_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6504\,
            in2 => \_gnd_net_\,
            in3 => \N__6941\,
            lcout => \U111_CYCLE_SM_TEA_CPUn_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6400\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7131\,
            ce => \N__7075\,
            sr => \N__7046\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7177\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7131\,
            ce => \N__7075\,
            sr => \N__7046\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8615\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7127\,
            ce => \N__7086\,
            sr => \N__7047\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7127\,
            ce => \N__7086\,
            sr => \N__7047\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7210\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7127\,
            ce => \N__7086\,
            sr => \N__7047\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8430\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7127\,
            ce => \N__7086\,
            sr => \N__7047\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7953\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7127\,
            ce => \N__7086\,
            sr => \N__7047\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7006\,
            in1 => \N__6972\,
            in2 => \_gnd_net_\,
            in3 => \N__7321\,
            lcout => \un1_D_UM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__6861\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6945\,
            lcout => \N_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TCI_CPUn_0_i_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6897\,
            in2 => \_gnd_net_\,
            in3 => \N__6862\,
            lcout => \U111_CYCLE_SM_TCI_CPUn_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8608\,
            in1 => \N__8565\,
            in2 => \_gnd_net_\,
            in3 => \N__7323\,
            lcout => \un1_D_UM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8531\,
            in1 => \N__8484\,
            in2 => \_gnd_net_\,
            in3 => \N__8215\,
            lcout => \un1_D_UM_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8442\,
            in1 => \N__8422\,
            in2 => \_gnd_net_\,
            in3 => \N__7344\,
            lcout => \un1_D_UM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8348\,
            in1 => \N__8319\,
            in2 => \_gnd_net_\,
            in3 => \N__8217\,
            lcout => \un1_D_UU_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8283\,
            in1 => \N__8264\,
            in2 => \_gnd_net_\,
            in3 => \N__8216\,
            lcout => \un1_D_UM_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7350\,
            in1 => \N__7965\,
            in2 => \_gnd_net_\,
            in3 => \N__7942\,
            lcout => \un1_D_UM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI8QUM_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__7887\,
            in1 => \N__7769\,
            in2 => \_gnd_net_\,
            in3 => \N__7704\,
            lcout => \N_60_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7322\,
            in1 => \N__7227\,
            in2 => \_gnd_net_\,
            in3 => \N__7211\,
            lcout => \un1_D_UM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

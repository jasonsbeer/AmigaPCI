// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 8 2025 22:54:55

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    DRA,
    SIZ,
    CMA,
    A,
    TSn,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    VBENn,
    CUMBEn,
    CLKRAM,
    C3,
    ASn,
    LDSn,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40_OUT,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    DBRn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    TACKn,
    C1);

    input [9:0] DRA;
    input [1:0] SIZ;
    output [10:0] CMA;
    input [20:0] A;
    input TSn;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    input C3;
    output ASn;
    output LDSn;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40_OUT;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    input DBRn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    output TACKn;
    input C1;

    wire N__10288;
    wire N__10287;
    wire N__10286;
    wire N__10279;
    wire N__10278;
    wire N__10277;
    wire N__10270;
    wire N__10269;
    wire N__10268;
    wire N__10261;
    wire N__10260;
    wire N__10259;
    wire N__10252;
    wire N__10251;
    wire N__10250;
    wire N__10243;
    wire N__10242;
    wire N__10241;
    wire N__10234;
    wire N__10233;
    wire N__10232;
    wire N__10225;
    wire N__10224;
    wire N__10223;
    wire N__10216;
    wire N__10215;
    wire N__10214;
    wire N__10207;
    wire N__10206;
    wire N__10205;
    wire N__10198;
    wire N__10197;
    wire N__10196;
    wire N__10189;
    wire N__10188;
    wire N__10187;
    wire N__10180;
    wire N__10179;
    wire N__10178;
    wire N__10171;
    wire N__10170;
    wire N__10169;
    wire N__10162;
    wire N__10161;
    wire N__10160;
    wire N__10153;
    wire N__10152;
    wire N__10151;
    wire N__10144;
    wire N__10143;
    wire N__10142;
    wire N__10135;
    wire N__10134;
    wire N__10133;
    wire N__10126;
    wire N__10125;
    wire N__10124;
    wire N__10117;
    wire N__10116;
    wire N__10115;
    wire N__10108;
    wire N__10107;
    wire N__10106;
    wire N__10099;
    wire N__10098;
    wire N__10097;
    wire N__10090;
    wire N__10089;
    wire N__10088;
    wire N__10081;
    wire N__10080;
    wire N__10079;
    wire N__10072;
    wire N__10071;
    wire N__10070;
    wire N__10063;
    wire N__10062;
    wire N__10061;
    wire N__10054;
    wire N__10053;
    wire N__10052;
    wire N__10045;
    wire N__10044;
    wire N__10043;
    wire N__10036;
    wire N__10035;
    wire N__10034;
    wire N__10027;
    wire N__10026;
    wire N__10025;
    wire N__10018;
    wire N__10017;
    wire N__10016;
    wire N__10009;
    wire N__10008;
    wire N__10007;
    wire N__10000;
    wire N__9999;
    wire N__9998;
    wire N__9991;
    wire N__9990;
    wire N__9989;
    wire N__9982;
    wire N__9981;
    wire N__9980;
    wire N__9973;
    wire N__9972;
    wire N__9971;
    wire N__9964;
    wire N__9963;
    wire N__9962;
    wire N__9955;
    wire N__9954;
    wire N__9953;
    wire N__9946;
    wire N__9945;
    wire N__9944;
    wire N__9937;
    wire N__9936;
    wire N__9935;
    wire N__9928;
    wire N__9927;
    wire N__9926;
    wire N__9919;
    wire N__9918;
    wire N__9917;
    wire N__9910;
    wire N__9909;
    wire N__9908;
    wire N__9901;
    wire N__9900;
    wire N__9899;
    wire N__9892;
    wire N__9891;
    wire N__9890;
    wire N__9883;
    wire N__9882;
    wire N__9881;
    wire N__9874;
    wire N__9873;
    wire N__9872;
    wire N__9865;
    wire N__9864;
    wire N__9863;
    wire N__9856;
    wire N__9855;
    wire N__9854;
    wire N__9847;
    wire N__9846;
    wire N__9845;
    wire N__9838;
    wire N__9837;
    wire N__9836;
    wire N__9829;
    wire N__9828;
    wire N__9827;
    wire N__9820;
    wire N__9819;
    wire N__9818;
    wire N__9811;
    wire N__9810;
    wire N__9809;
    wire N__9802;
    wire N__9801;
    wire N__9800;
    wire N__9793;
    wire N__9792;
    wire N__9791;
    wire N__9784;
    wire N__9783;
    wire N__9782;
    wire N__9775;
    wire N__9774;
    wire N__9773;
    wire N__9766;
    wire N__9765;
    wire N__9764;
    wire N__9757;
    wire N__9756;
    wire N__9755;
    wire N__9748;
    wire N__9747;
    wire N__9746;
    wire N__9739;
    wire N__9738;
    wire N__9737;
    wire N__9730;
    wire N__9729;
    wire N__9728;
    wire N__9721;
    wire N__9720;
    wire N__9719;
    wire N__9712;
    wire N__9711;
    wire N__9710;
    wire N__9703;
    wire N__9702;
    wire N__9701;
    wire N__9694;
    wire N__9693;
    wire N__9692;
    wire N__9685;
    wire N__9684;
    wire N__9683;
    wire N__9676;
    wire N__9675;
    wire N__9674;
    wire N__9667;
    wire N__9666;
    wire N__9665;
    wire N__9658;
    wire N__9657;
    wire N__9656;
    wire N__9649;
    wire N__9648;
    wire N__9647;
    wire N__9640;
    wire N__9639;
    wire N__9638;
    wire N__9631;
    wire N__9630;
    wire N__9629;
    wire N__9622;
    wire N__9621;
    wire N__9620;
    wire N__9613;
    wire N__9612;
    wire N__9611;
    wire N__9604;
    wire N__9603;
    wire N__9602;
    wire N__9595;
    wire N__9594;
    wire N__9593;
    wire N__9586;
    wire N__9585;
    wire N__9584;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9555;
    wire N__9552;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9528;
    wire N__9525;
    wire N__9522;
    wire N__9519;
    wire N__9516;
    wire N__9513;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9503;
    wire N__9502;
    wire N__9501;
    wire N__9500;
    wire N__9499;
    wire N__9498;
    wire N__9495;
    wire N__9480;
    wire N__9477;
    wire N__9474;
    wire N__9471;
    wire N__9470;
    wire N__9469;
    wire N__9468;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9451;
    wire N__9446;
    wire N__9443;
    wire N__9438;
    wire N__9435;
    wire N__9430;
    wire N__9427;
    wire N__9424;
    wire N__9417;
    wire N__9416;
    wire N__9415;
    wire N__9414;
    wire N__9413;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9394;
    wire N__9393;
    wire N__9392;
    wire N__9391;
    wire N__9388;
    wire N__9387;
    wire N__9386;
    wire N__9385;
    wire N__9382;
    wire N__9381;
    wire N__9380;
    wire N__9379;
    wire N__9378;
    wire N__9377;
    wire N__9376;
    wire N__9375;
    wire N__9372;
    wire N__9371;
    wire N__9370;
    wire N__9369;
    wire N__9368;
    wire N__9367;
    wire N__9366;
    wire N__9365;
    wire N__9364;
    wire N__9363;
    wire N__9360;
    wire N__9359;
    wire N__9358;
    wire N__9357;
    wire N__9356;
    wire N__9355;
    wire N__9354;
    wire N__9351;
    wire N__9350;
    wire N__9349;
    wire N__9348;
    wire N__9347;
    wire N__9346;
    wire N__9345;
    wire N__9342;
    wire N__9341;
    wire N__9340;
    wire N__9339;
    wire N__9338;
    wire N__9337;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9219;
    wire N__9216;
    wire N__9213;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9159;
    wire N__9156;
    wire N__9153;
    wire N__9150;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9138;
    wire N__9135;
    wire N__9132;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9105;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9093;
    wire N__9090;
    wire N__9087;
    wire N__9084;
    wire N__9083;
    wire N__9082;
    wire N__9081;
    wire N__9078;
    wire N__9075;
    wire N__9072;
    wire N__9069;
    wire N__9066;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9038;
    wire N__9033;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9021;
    wire N__9018;
    wire N__9015;
    wire N__9012;
    wire N__9009;
    wire N__9006;
    wire N__9003;
    wire N__9000;
    wire N__8997;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8985;
    wire N__8982;
    wire N__8979;
    wire N__8976;
    wire N__8973;
    wire N__8970;
    wire N__8967;
    wire N__8964;
    wire N__8961;
    wire N__8958;
    wire N__8955;
    wire N__8952;
    wire N__8949;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8922;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8901;
    wire N__8898;
    wire N__8895;
    wire N__8892;
    wire N__8889;
    wire N__8888;
    wire N__8883;
    wire N__8880;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8870;
    wire N__8869;
    wire N__8868;
    wire N__8867;
    wire N__8866;
    wire N__8865;
    wire N__8862;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8840;
    wire N__8837;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8793;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8781;
    wire N__8778;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8754;
    wire N__8751;
    wire N__8748;
    wire N__8745;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8720;
    wire N__8719;
    wire N__8718;
    wire N__8715;
    wire N__8712;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8691;
    wire N__8688;
    wire N__8685;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8640;
    wire N__8637;
    wire N__8636;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8622;
    wire N__8619;
    wire N__8616;
    wire N__8613;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8595;
    wire N__8592;
    wire N__8589;
    wire N__8588;
    wire N__8585;
    wire N__8584;
    wire N__8583;
    wire N__8580;
    wire N__8579;
    wire N__8578;
    wire N__8577;
    wire N__8576;
    wire N__8573;
    wire N__8572;
    wire N__8571;
    wire N__8570;
    wire N__8569;
    wire N__8566;
    wire N__8563;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8552;
    wire N__8549;
    wire N__8548;
    wire N__8545;
    wire N__8544;
    wire N__8543;
    wire N__8540;
    wire N__8539;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8531;
    wire N__8530;
    wire N__8521;
    wire N__8518;
    wire N__8517;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8497;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8473;
    wire N__8468;
    wire N__8465;
    wire N__8456;
    wire N__8453;
    wire N__8444;
    wire N__8437;
    wire N__8432;
    wire N__8429;
    wire N__8424;
    wire N__8421;
    wire N__8412;
    wire N__8409;
    wire N__8406;
    wire N__8403;
    wire N__8400;
    wire N__8399;
    wire N__8398;
    wire N__8395;
    wire N__8394;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8386;
    wire N__8385;
    wire N__8382;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8365;
    wire N__8364;
    wire N__8361;
    wire N__8360;
    wire N__8359;
    wire N__8358;
    wire N__8357;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8343;
    wire N__8342;
    wire N__8341;
    wire N__8340;
    wire N__8339;
    wire N__8338;
    wire N__8337;
    wire N__8336;
    wire N__8335;
    wire N__8334;
    wire N__8331;
    wire N__8330;
    wire N__8327;
    wire N__8318;
    wire N__8315;
    wire N__8312;
    wire N__8307;
    wire N__8302;
    wire N__8291;
    wire N__8282;
    wire N__8275;
    wire N__8262;
    wire N__8259;
    wire N__8258;
    wire N__8257;
    wire N__8256;
    wire N__8253;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8245;
    wire N__8242;
    wire N__8239;
    wire N__8234;
    wire N__8231;
    wire N__8226;
    wire N__8225;
    wire N__8224;
    wire N__8219;
    wire N__8214;
    wire N__8211;
    wire N__8210;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8196;
    wire N__8187;
    wire N__8186;
    wire N__8185;
    wire N__8184;
    wire N__8183;
    wire N__8182;
    wire N__8179;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8151;
    wire N__8148;
    wire N__8145;
    wire N__8142;
    wire N__8139;
    wire N__8136;
    wire N__8133;
    wire N__8130;
    wire N__8127;
    wire N__8124;
    wire N__8123;
    wire N__8122;
    wire N__8121;
    wire N__8120;
    wire N__8119;
    wire N__8118;
    wire N__8117;
    wire N__8116;
    wire N__8115;
    wire N__8114;
    wire N__8113;
    wire N__8112;
    wire N__8111;
    wire N__8110;
    wire N__8109;
    wire N__8108;
    wire N__8107;
    wire N__8106;
    wire N__8105;
    wire N__8104;
    wire N__8103;
    wire N__8102;
    wire N__8101;
    wire N__8100;
    wire N__8099;
    wire N__8096;
    wire N__8095;
    wire N__8094;
    wire N__8093;
    wire N__8092;
    wire N__8091;
    wire N__8090;
    wire N__8089;
    wire N__8088;
    wire N__8019;
    wire N__8016;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8008;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7989;
    wire N__7986;
    wire N__7985;
    wire N__7984;
    wire N__7981;
    wire N__7978;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7959;
    wire N__7954;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7940;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7911;
    wire N__7908;
    wire N__7905;
    wire N__7902;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7890;
    wire N__7887;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7872;
    wire N__7869;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7854;
    wire N__7851;
    wire N__7850;
    wire N__7847;
    wire N__7844;
    wire N__7839;
    wire N__7836;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7824;
    wire N__7821;
    wire N__7818;
    wire N__7815;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7800;
    wire N__7797;
    wire N__7794;
    wire N__7791;
    wire N__7788;
    wire N__7785;
    wire N__7784;
    wire N__7783;
    wire N__7782;
    wire N__7781;
    wire N__7780;
    wire N__7779;
    wire N__7774;
    wire N__7773;
    wire N__7766;
    wire N__7761;
    wire N__7760;
    wire N__7759;
    wire N__7756;
    wire N__7753;
    wire N__7750;
    wire N__7747;
    wire N__7742;
    wire N__7737;
    wire N__7734;
    wire N__7729;
    wire N__7728;
    wire N__7725;
    wire N__7720;
    wire N__7717;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7683;
    wire N__7682;
    wire N__7681;
    wire N__7678;
    wire N__7675;
    wire N__7674;
    wire N__7673;
    wire N__7672;
    wire N__7671;
    wire N__7668;
    wire N__7663;
    wire N__7660;
    wire N__7653;
    wire N__7650;
    wire N__7641;
    wire N__7638;
    wire N__7635;
    wire N__7632;
    wire N__7629;
    wire N__7626;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7602;
    wire N__7599;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7581;
    wire N__7578;
    wire N__7575;
    wire N__7572;
    wire N__7569;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7551;
    wire N__7548;
    wire N__7545;
    wire N__7542;
    wire N__7539;
    wire N__7536;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7512;
    wire N__7509;
    wire N__7508;
    wire N__7505;
    wire N__7504;
    wire N__7501;
    wire N__7500;
    wire N__7499;
    wire N__7496;
    wire N__7495;
    wire N__7492;
    wire N__7489;
    wire N__7486;
    wire N__7483;
    wire N__7480;
    wire N__7477;
    wire N__7476;
    wire N__7473;
    wire N__7468;
    wire N__7465;
    wire N__7462;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7440;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7426;
    wire N__7425;
    wire N__7422;
    wire N__7419;
    wire N__7414;
    wire N__7407;
    wire N__7404;
    wire N__7401;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7389;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7374;
    wire N__7371;
    wire N__7368;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7356;
    wire N__7353;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7341;
    wire N__7338;
    wire N__7335;
    wire N__7334;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7317;
    wire N__7316;
    wire N__7313;
    wire N__7310;
    wire N__7305;
    wire N__7302;
    wire N__7299;
    wire N__7296;
    wire N__7293;
    wire N__7290;
    wire N__7287;
    wire N__7284;
    wire N__7281;
    wire N__7278;
    wire N__7275;
    wire N__7272;
    wire N__7269;
    wire N__7266;
    wire N__7263;
    wire N__7260;
    wire N__7259;
    wire N__7258;
    wire N__7255;
    wire N__7250;
    wire N__7247;
    wire N__7244;
    wire N__7243;
    wire N__7240;
    wire N__7237;
    wire N__7234;
    wire N__7227;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7219;
    wire N__7218;
    wire N__7213;
    wire N__7208;
    wire N__7207;
    wire N__7206;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7194;
    wire N__7185;
    wire N__7182;
    wire N__7179;
    wire N__7176;
    wire N__7173;
    wire N__7170;
    wire N__7167;
    wire N__7164;
    wire N__7161;
    wire N__7158;
    wire N__7155;
    wire N__7152;
    wire N__7149;
    wire N__7148;
    wire N__7147;
    wire N__7146;
    wire N__7143;
    wire N__7136;
    wire N__7131;
    wire N__7128;
    wire N__7125;
    wire N__7122;
    wire N__7119;
    wire N__7116;
    wire N__7113;
    wire N__7110;
    wire N__7107;
    wire N__7104;
    wire N__7101;
    wire N__7098;
    wire N__7095;
    wire N__7092;
    wire N__7091;
    wire N__7086;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7074;
    wire N__7071;
    wire N__7068;
    wire N__7065;
    wire N__7062;
    wire N__7061;
    wire N__7058;
    wire N__7053;
    wire N__7050;
    wire N__7049;
    wire N__7046;
    wire N__7043;
    wire N__7038;
    wire N__7035;
    wire N__7032;
    wire N__7029;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7017;
    wire N__7014;
    wire N__7011;
    wire N__7008;
    wire N__7005;
    wire N__7002;
    wire N__6999;
    wire N__6996;
    wire N__6993;
    wire N__6990;
    wire N__6987;
    wire N__6984;
    wire N__6981;
    wire N__6980;
    wire N__6979;
    wire N__6978;
    wire N__6973;
    wire N__6970;
    wire N__6967;
    wire N__6962;
    wire N__6959;
    wire N__6956;
    wire N__6953;
    wire N__6950;
    wire N__6945;
    wire N__6942;
    wire N__6941;
    wire N__6940;
    wire N__6939;
    wire N__6936;
    wire N__6929;
    wire N__6924;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6900;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6879;
    wire N__6876;
    wire N__6873;
    wire N__6870;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6852;
    wire N__6849;
    wire N__6846;
    wire N__6843;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6813;
    wire N__6810;
    wire N__6807;
    wire N__6804;
    wire N__6801;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6789;
    wire N__6786;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6762;
    wire N__6759;
    wire N__6756;
    wire N__6753;
    wire N__6750;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6732;
    wire N__6729;
    wire N__6726;
    wire N__6723;
    wire N__6722;
    wire N__6721;
    wire N__6718;
    wire N__6715;
    wire N__6712;
    wire N__6707;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6681;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6639;
    wire N__6638;
    wire N__6637;
    wire N__6636;
    wire N__6635;
    wire N__6632;
    wire N__6631;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6616;
    wire N__6615;
    wire N__6614;
    wire N__6609;
    wire N__6608;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6594;
    wire N__6593;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6575;
    wire N__6568;
    wire N__6555;
    wire N__6552;
    wire N__6551;
    wire N__6550;
    wire N__6549;
    wire N__6546;
    wire N__6543;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6535;
    wire N__6534;
    wire N__6529;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6515;
    wire N__6504;
    wire N__6503;
    wire N__6502;
    wire N__6499;
    wire N__6496;
    wire N__6491;
    wire N__6486;
    wire N__6485;
    wire N__6484;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6468;
    wire N__6465;
    wire N__6462;
    wire N__6459;
    wire N__6456;
    wire N__6447;
    wire N__6444;
    wire N__6443;
    wire N__6440;
    wire N__6439;
    wire N__6438;
    wire N__6435;
    wire N__6432;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6418;
    wire N__6415;
    wire N__6414;
    wire N__6413;
    wire N__6412;
    wire N__6409;
    wire N__6404;
    wire N__6397;
    wire N__6390;
    wire N__6387;
    wire N__6386;
    wire N__6385;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6373;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6357;
    wire N__6354;
    wire N__6351;
    wire N__6348;
    wire N__6345;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6333;
    wire N__6332;
    wire N__6327;
    wire N__6326;
    wire N__6325;
    wire N__6322;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6306;
    wire N__6305;
    wire N__6304;
    wire N__6301;
    wire N__6296;
    wire N__6293;
    wire N__6290;
    wire N__6285;
    wire N__6284;
    wire N__6283;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6251;
    wire N__6246;
    wire N__6243;
    wire N__6242;
    wire N__6241;
    wire N__6234;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6216;
    wire N__6213;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6200;
    wire N__6199;
    wire N__6194;
    wire N__6191;
    wire N__6186;
    wire N__6183;
    wire N__6180;
    wire N__6177;
    wire N__6174;
    wire N__6171;
    wire N__6168;
    wire N__6165;
    wire N__6162;
    wire N__6159;
    wire N__6156;
    wire N__6153;
    wire N__6150;
    wire N__6147;
    wire N__6144;
    wire N__6141;
    wire N__6138;
    wire N__6137;
    wire N__6136;
    wire N__6129;
    wire N__6126;
    wire N__6125;
    wire N__6124;
    wire N__6123;
    wire N__6120;
    wire N__6115;
    wire N__6112;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6084;
    wire N__6081;
    wire N__6080;
    wire N__6077;
    wire N__6074;
    wire N__6073;
    wire N__6070;
    wire N__6065;
    wire N__6060;
    wire N__6057;
    wire N__6054;
    wire N__6051;
    wire N__6048;
    wire N__6045;
    wire N__6044;
    wire N__6039;
    wire N__6036;
    wire N__6033;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5985;
    wire N__5982;
    wire N__5979;
    wire N__5976;
    wire N__5973;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5961;
    wire N__5958;
    wire N__5955;
    wire N__5954;
    wire N__5951;
    wire N__5948;
    wire N__5945;
    wire N__5942;
    wire N__5941;
    wire N__5940;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5919;
    wire N__5918;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5886;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5865;
    wire N__5864;
    wire N__5863;
    wire N__5860;
    wire N__5855;
    wire N__5850;
    wire N__5847;
    wire N__5846;
    wire N__5843;
    wire N__5842;
    wire N__5839;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5823;
    wire N__5822;
    wire N__5821;
    wire N__5818;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5800;
    wire N__5793;
    wire N__5790;
    wire N__5787;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5775;
    wire N__5772;
    wire N__5769;
    wire N__5766;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5754;
    wire N__5751;
    wire N__5748;
    wire N__5745;
    wire N__5742;
    wire N__5739;
    wire N__5736;
    wire N__5733;
    wire N__5730;
    wire N__5727;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5709;
    wire N__5706;
    wire N__5703;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5682;
    wire N__5679;
    wire N__5676;
    wire N__5673;
    wire N__5670;
    wire N__5667;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5634;
    wire N__5631;
    wire N__5628;
    wire N__5627;
    wire N__5626;
    wire N__5625;
    wire N__5624;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5616;
    wire N__5615;
    wire N__5610;
    wire N__5609;
    wire N__5608;
    wire N__5607;
    wire N__5606;
    wire N__5605;
    wire N__5604;
    wire N__5603;
    wire N__5602;
    wire N__5597;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5586;
    wire N__5585;
    wire N__5584;
    wire N__5583;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5563;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5543;
    wire N__5538;
    wire N__5531;
    wire N__5508;
    wire N__5507;
    wire N__5504;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5496;
    wire N__5495;
    wire N__5494;
    wire N__5493;
    wire N__5492;
    wire N__5491;
    wire N__5490;
    wire N__5487;
    wire N__5486;
    wire N__5485;
    wire N__5482;
    wire N__5481;
    wire N__5480;
    wire N__5479;
    wire N__5478;
    wire N__5477;
    wire N__5474;
    wire N__5469;
    wire N__5466;
    wire N__5459;
    wire N__5456;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5432;
    wire N__5423;
    wire N__5418;
    wire N__5403;
    wire N__5400;
    wire N__5399;
    wire N__5398;
    wire N__5397;
    wire N__5394;
    wire N__5391;
    wire N__5390;
    wire N__5387;
    wire N__5386;
    wire N__5385;
    wire N__5382;
    wire N__5379;
    wire N__5376;
    wire N__5373;
    wire N__5368;
    wire N__5365;
    wire N__5352;
    wire N__5349;
    wire N__5346;
    wire N__5343;
    wire N__5340;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5325;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5313;
    wire N__5312;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5295;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5280;
    wire N__5279;
    wire N__5278;
    wire N__5275;
    wire N__5270;
    wire N__5265;
    wire N__5262;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5210;
    wire N__5205;
    wire N__5202;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5190;
    wire N__5189;
    wire N__5188;
    wire N__5187;
    wire N__5180;
    wire N__5177;
    wire N__5172;
    wire N__5171;
    wire N__5170;
    wire N__5165;
    wire N__5162;
    wire N__5157;
    wire N__5156;
    wire N__5155;
    wire N__5152;
    wire N__5147;
    wire N__5142;
    wire N__5141;
    wire N__5136;
    wire N__5133;
    wire N__5130;
    wire N__5127;
    wire N__5124;
    wire N__5121;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5111;
    wire N__5106;
    wire N__5103;
    wire N__5102;
    wire N__5101;
    wire N__5100;
    wire N__5099;
    wire N__5096;
    wire N__5091;
    wire N__5088;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5072;
    wire N__5067;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5046;
    wire N__5043;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5028;
    wire N__5027;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5015;
    wire N__5010;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4963;
    wire N__4958;
    wire N__4955;
    wire N__4950;
    wire N__4949;
    wire N__4948;
    wire N__4943;
    wire N__4942;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4913;
    wire N__4912;
    wire N__4911;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4903;
    wire N__4900;
    wire N__4895;
    wire N__4890;
    wire N__4887;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4871;
    wire N__4870;
    wire N__4869;
    wire N__4868;
    wire N__4865;
    wire N__4864;
    wire N__4861;
    wire N__4860;
    wire N__4857;
    wire N__4856;
    wire N__4855;
    wire N__4854;
    wire N__4853;
    wire N__4852;
    wire N__4851;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4831;
    wire N__4826;
    wire N__4821;
    wire N__4816;
    wire N__4813;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4777;
    wire N__4776;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4749;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4737;
    wire N__4736;
    wire N__4733;
    wire N__4730;
    wire N__4725;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4710;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4698;
    wire N__4695;
    wire N__4692;
    wire N__4689;
    wire N__4688;
    wire N__4685;
    wire N__4682;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4670;
    wire N__4669;
    wire N__4666;
    wire N__4663;
    wire N__4662;
    wire N__4661;
    wire N__4660;
    wire N__4659;
    wire N__4658;
    wire N__4655;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4647;
    wire N__4644;
    wire N__4643;
    wire N__4642;
    wire N__4639;
    wire N__4636;
    wire N__4633;
    wire N__4630;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4614;
    wire N__4609;
    wire N__4604;
    wire N__4587;
    wire N__4584;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4544;
    wire N__4543;
    wire N__4538;
    wire N__4535;
    wire N__4530;
    wire N__4529;
    wire N__4524;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4494;
    wire N__4491;
    wire N__4488;
    wire N__4487;
    wire N__4482;
    wire N__4479;
    wire N__4476;
    wire N__4473;
    wire N__4470;
    wire N__4467;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4382;
    wire N__4381;
    wire N__4376;
    wire N__4373;
    wire N__4368;
    wire N__4365;
    wire N__4364;
    wire N__4361;
    wire N__4360;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4338;
    wire N__4337;
    wire N__4336;
    wire N__4335;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4317;
    wire N__4314;
    wire N__4313;
    wire N__4312;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4298;
    wire N__4295;
    wire N__4290;
    wire N__4287;
    wire N__4286;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4263;
    wire N__4260;
    wire N__4259;
    wire N__4258;
    wire N__4257;
    wire N__4256;
    wire N__4255;
    wire N__4254;
    wire N__4253;
    wire N__4250;
    wire N__4243;
    wire N__4236;
    wire N__4233;
    wire N__4224;
    wire N__4221;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4209;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4197;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4172;
    wire N__4171;
    wire N__4168;
    wire N__4163;
    wire N__4160;
    wire N__4155;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4147;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4129;
    wire N__4122;
    wire N__4119;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4107;
    wire N__4106;
    wire N__4105;
    wire N__4102;
    wire N__4101;
    wire N__4100;
    wire N__4095;
    wire N__4092;
    wire N__4089;
    wire N__4086;
    wire N__4077;
    wire N__4076;
    wire N__4075;
    wire N__4072;
    wire N__4067;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4038;
    wire N__4035;
    wire N__4032;
    wire N__4029;
    wire N__4026;
    wire N__4023;
    wire N__4020;
    wire N__4017;
    wire N__4014;
    wire N__4011;
    wire N__4008;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3987;
    wire N__3984;
    wire N__3981;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3963;
    wire N__3960;
    wire N__3957;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3900;
    wire N__3897;
    wire N__3894;
    wire N__3891;
    wire N__3888;
    wire N__3885;
    wire N__3882;
    wire N__3879;
    wire N__3876;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3845;
    wire N__3840;
    wire N__3837;
    wire N__3834;
    wire N__3831;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3819;
    wire N__3816;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3804;
    wire N__3801;
    wire N__3798;
    wire N__3795;
    wire N__3792;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3759;
    wire N__3756;
    wire N__3753;
    wire N__3750;
    wire N__3747;
    wire N__3744;
    wire N__3741;
    wire N__3738;
    wire N__3735;
    wire N__3732;
    wire N__3729;
    wire N__3726;
    wire N__3723;
    wire N__3722;
    wire N__3721;
    wire N__3716;
    wire N__3713;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3696;
    wire N__3693;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3681;
    wire N__3678;
    wire N__3675;
    wire N__3672;
    wire N__3669;
    wire N__3666;
    wire N__3663;
    wire N__3660;
    wire N__3657;
    wire N__3654;
    wire N__3651;
    wire N__3648;
    wire N__3645;
    wire N__3642;
    wire N__3639;
    wire N__3636;
    wire N__3633;
    wire N__3630;
    wire N__3627;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK40_PLL_i_i;
    wire N_897_i;
    wire CLK80_PLL_i_i;
    wire \U712_CHIP_RAM.N_193_cascade_ ;
    wire \U712_CHIP_RAM.N_176_cascade_ ;
    wire \U712_CHIP_RAM.N_253_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0 ;
    wire \U712_CHIP_RAM.N_298_cascade_ ;
    wire \U712_CHIP_RAM.N_323_cascade_ ;
    wire \U712_CHIP_RAM.N_304 ;
    wire \U712_CHIP_RAM.N_216 ;
    wire \U712_CHIP_RAM.N_216_cascade_ ;
    wire C3_c;
    wire \U712_CHIP_RAM.N_213 ;
    wire VBENn_c;
    wire A_c_12;
    wire A_c_5;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ;
    wire A_c_18;
    wire A_c_16;
    wire A_c_10;
    wire A_c_3;
    wire A_c_9;
    wire A_c_2;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_193 ;
    wire \U712_CHIP_RAM.N_177_cascade_ ;
    wire \U712_CHIP_RAM.N_223 ;
    wire \U712_CHIP_RAM.N_300 ;
    wire \U712_CHIP_RAM.N_223_cascade_ ;
    wire \U712_CHIP_RAM.N_187_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_1_cascade_ ;
    wire \U712_CHIP_RAM.N_264_cascade_ ;
    wire \U712_CHIP_RAM.N_262 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0 ;
    wire \U712_CHIP_RAM.N_220 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0_1 ;
    wire \U712_CHIP_RAM.N_323 ;
    wire \U712_CHIP_RAM.N_176 ;
    wire \U712_CHIP_RAM.N_242_cascade_ ;
    wire \U712_CHIP_RAM.N_319 ;
    wire \U712_CHIP_RAM.N_307 ;
    wire \U712_CHIP_RAM.N_177 ;
    wire \U712_CHIP_RAM.N_319_cascade_ ;
    wire \U712_CHIP_RAM.N_322 ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_311 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_i_i_a3_0 ;
    wire bfn_8_8_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.N_46 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.N_256_i ;
    wire \U712_CYCLE_TERM.N_207_i_0_en_cascade_ ;
    wire TACK_EN_i_ess;
    wire \U712_CYCLE_TERM.N_207_i_0_en_0 ;
    wire \U712_REG_SM.N_185_cascade_ ;
    wire C1_c;
    wire \U712_REG_SM.N_197_cascade_ ;
    wire \U712_REG_SM.C1_SYNCZ0Z_2 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.DS_EN_0_sqmuxa_0_a2_0_a3_1_cascade_ ;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.DS_EN_0_sqmuxa_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_6 ;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ;
    wire A_c_14;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ;
    wire A_c_15;
    wire A_c_8;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_42_1 ;
    wire \U712_CHIP_RAM.N_236 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_1 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_198_i ;
    wire \U712_CHIP_RAM.N_187 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.N_355_cascade_ ;
    wire \U712_CHIP_RAM.N_321 ;
    wire \U712_CHIP_RAM.N_235 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.N_217 ;
    wire \U712_CHIP_RAM.CPU_TACK_8_iv_i_i_2_cascade_ ;
    wire \U712_CHIP_RAM.N_219 ;
    wire \U712_CHIP_RAM.N_117_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_i_0_1 ;
    wire CPU_TACKm;
    wire \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861Z0Z_1 ;
    wire RAMSPACEn_c;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.N_197 ;
    wire \U712_REG_SM.N_215_cascade_ ;
    wire ASn_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_2 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_185 ;
    wire \U712_REG_SM.N_204_cascade_ ;
    wire \U712_REG_SM.N_215 ;
    wire \U712_REG_SM.N_204 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire TSn_c;
    wire REGSPACEn_c;
    wire \U712_REG_SM.REG_CYCLE_GOZ0 ;
    wire \U712_REG_SM.N_209 ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.DS_EN_0_sqmuxa ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire DBR_SYNCZ0Z_0;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire CMA_c_5;
    wire A_c_6;
    wire A_c_13;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ;
    wire A_c_4;
    wire A_c_11;
    wire A_c_7;
    wire \U712_CHIP_RAM.N_324_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_301 ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0 ;
    wire \U712_CHIP_RAM.N_242 ;
    wire \U712_CHIP_RAM.DBENn_7_0 ;
    wire \U712_CHIP_RAM.N_253 ;
    wire REG_TACK;
    wire \U712_CHIP_RAM.REFRESH_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_188 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire RAS1n_c;
    wire \U712_CHIP_RAM.REFRESH_SYNCZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.N_200 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_5 ;
    wire TACK_OUTn;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire A_c_1;
    wire SIZ_c_1;
    wire REG_CYCLEm;
    wire DRDENn_c;
    wire un1_LDSn_i_0;
    wire A_c_0;
    wire SIZ_c_0;
    wire DS_ENm;
    wire un1_UDSn_i_0;
    wire RnW_c;
    wire N_212;
    wire CONSTANT_ONE_NET;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire AWEn_c;
    wire DBDIR_c;
    wire \U712_CHIP_RAM.N_298 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_355 ;
    wire \U712_CHIP_RAM.BANK0_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_305 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ;
    wire \U712_CHIP_RAM.un5_DMA_CYCLE_START_0 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire CLK40_PLL_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_BYTE_ENABLE.N_275 ;
    wire N_148_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ;
    wire \U712_BYTE_ENABLE.N_271 ;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0_cascade_ ;
    wire N_171_i;
    wire DBENn_c;
    wire DMA_CYCLEm;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0 ;
    wire \U712_BYTE_ENABLE.N_277 ;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0_cascade_ ;
    wire N_150_i;
    wire \U712_BYTE_ENABLE.N_270 ;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0 ;
    wire \U712_BYTE_ENABLE.N_273 ;
    wire N_172_i;
    wire CASLn_c;
    wire CASUn_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire WEn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire A_c_17;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_12_8_0_;
    wire \U712_CHIP_RAM.REFRESH5lto1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH5lto2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire RESETn_c;
    wire RESETn_c_i;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire CASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire CMA_c_4;
    wire CPU_CYCLEm;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_ ;
    wire CMA_c_7;
    wire CLK80_PLL;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire RAS0n_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire C1_c_g;
    wire DBRn_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire _gnd_net_;
    wire C3_c_g;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ;
    wire RESETn_c_i_g;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__3645),
            .RESETB(N__6789),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__10288),
            .DIN(N__10287),
            .DOUT(N__10286),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__10288),
            .PADOUT(N__10287),
            .PADIN(N__10286),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7266),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__10279),
            .DIN(N__10278),
            .DOUT(N__10277),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__10279),
            .PADOUT(N__10278),
            .PADIN(N__10277),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__10270),
            .DIN(N__10269),
            .DOUT(N__10268),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__10270),
            .PADOUT(N__10269),
            .PADIN(N__10268),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8742),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__10261),
            .DIN(N__10260),
            .DOUT(N__10259),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__10261),
            .PADOUT(N__10260),
            .PADIN(N__10259),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6810),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__10252),
            .DIN(N__10251),
            .DOUT(N__10250),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__10252),
            .PADOUT(N__10251),
            .PADIN(N__10250),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__10243),
            .DIN(N__10242),
            .DOUT(N__10241),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__10243),
            .PADOUT(N__10242),
            .PADIN(N__10241),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__10234),
            .DIN(N__10233),
            .DOUT(N__10232),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__10234),
            .PADOUT(N__10233),
            .PADIN(N__10232),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__10225),
            .DIN(N__10224),
            .DOUT(N__10223),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__10225),
            .PADOUT(N__10224),
            .PADIN(N__10223),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__10216),
            .DIN(N__10215),
            .DOUT(N__10214),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__10216),
            .PADOUT(N__10215),
            .PADIN(N__10214),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__10207),
            .DIN(N__10206),
            .DOUT(N__10205),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__10207),
            .PADOUT(N__10206),
            .PADIN(N__10205),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__10198),
            .DIN(N__10197),
            .DOUT(N__10196),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__10198),
            .PADOUT(N__10197),
            .PADIN(N__10196),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8148),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__10189),
            .DIN(N__10188),
            .DOUT(N__10187),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__10189),
            .PADOUT(N__10188),
            .PADIN(N__10187),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__10180),
            .DIN(N__10179),
            .DOUT(N__10178),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__10180),
            .PADOUT(N__10179),
            .PADIN(N__10178),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__10171),
            .DIN(N__10170),
            .DOUT(N__10169),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__10171),
            .PADOUT(N__10170),
            .PADIN(N__10169),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__10162),
            .DIN(N__10161),
            .DOUT(N__10160),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__10162),
            .PADOUT(N__10161),
            .PADIN(N__10160),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3831),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__10153),
            .DIN(N__10152),
            .DOUT(N__10151),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__10153),
            .PADOUT(N__10152),
            .PADIN(N__10151),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__10144),
            .DIN(N__10143),
            .DOUT(N__10142),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__10144),
            .PADOUT(N__10143),
            .PADIN(N__10142),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__10135),
            .DIN(N__10134),
            .DOUT(N__10133),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__10135),
            .PADOUT(N__10134),
            .PADIN(N__10133),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8652),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__10126),
            .DIN(N__10125),
            .DOUT(N__10124),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__10126),
            .PADOUT(N__10125),
            .PADIN(N__10124),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__10117),
            .DIN(N__10116),
            .DOUT(N__10115),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__10117),
            .PADOUT(N__10116),
            .PADIN(N__10115),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8676),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__10108),
            .DIN(N__10107),
            .DOUT(N__10106),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__10108),
            .PADOUT(N__10107),
            .PADIN(N__10106),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__10099),
            .DIN(N__10098),
            .DOUT(N__10097),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__10099),
            .PADOUT(N__10098),
            .PADIN(N__10097),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__10090),
            .DIN(N__10089),
            .DOUT(N__10088),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__10090),
            .PADOUT(N__10089),
            .PADIN(N__10088),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__10081),
            .DIN(N__10080),
            .DOUT(N__10079),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__10081),
            .PADOUT(N__10080),
            .PADIN(N__10079),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__10072),
            .DIN(N__10071),
            .DOUT(N__10070),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__10072),
            .PADOUT(N__10071),
            .PADIN(N__10070),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__10063),
            .DIN(N__10062),
            .DOUT(N__10061),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__10063),
            .PADOUT(N__10062),
            .PADIN(N__10061),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5352),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__10054),
            .DIN(N__10053),
            .DOUT(N__10052),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__10054),
            .PADOUT(N__10053),
            .PADIN(N__10052),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__10045),
            .DIN(N__10044),
            .DOUT(N__10043),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__10045),
            .PADOUT(N__10044),
            .PADIN(N__10043),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__10036),
            .DIN(N__10035),
            .DOUT(N__10034),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__10036),
            .PADOUT(N__10035),
            .PADIN(N__10034),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__10027),
            .DIN(N__10026),
            .DOUT(N__10025),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__10027),
            .PADOUT(N__10026),
            .PADIN(N__10025),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__10018),
            .DIN(N__10017),
            .DOUT(N__10016),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__10018),
            .PADOUT(N__10017),
            .PADIN(N__10016),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__10009),
            .DIN(N__10008),
            .DOUT(N__10007),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__10009),
            .PADOUT(N__10008),
            .PADIN(N__10007),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7608),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__10000),
            .DIN(N__9999),
            .DOUT(N__9998),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__10000),
            .PADOUT(N__9999),
            .PADIN(N__9998),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__9991),
            .DIN(N__9990),
            .DOUT(N__9989),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__9991),
            .PADOUT(N__9990),
            .PADIN(N__9989),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__9982),
            .DIN(N__9981),
            .DOUT(N__9980),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__9982),
            .PADOUT(N__9981),
            .PADIN(N__9980),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__9973),
            .DIN(N__9972),
            .DOUT(N__9971),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__9973),
            .PADOUT(N__9972),
            .PADIN(N__9971),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__9964),
            .DIN(N__9963),
            .DOUT(N__9962),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__9964),
            .PADOUT(N__9963),
            .PADIN(N__9962),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6162),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__9955),
            .DIN(N__9954),
            .DOUT(N__9953),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__9955),
            .PADOUT(N__9954),
            .PADIN(N__9953),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__9946),
            .DIN(N__9945),
            .DOUT(N__9944),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__9946),
            .PADOUT(N__9945),
            .PADIN(N__9944),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7641),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__9937),
            .DIN(N__9936),
            .DOUT(N__9935),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__9937),
            .PADOUT(N__9936),
            .PADIN(N__9935),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__9928),
            .DIN(N__9927),
            .DOUT(N__9926),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__9928),
            .PADOUT(N__9927),
            .PADIN(N__9926),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__9919),
            .DIN(N__9918),
            .DOUT(N__9917),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__9919),
            .PADOUT(N__9918),
            .PADIN(N__9917),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3663),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__9910),
            .DIN(N__9909),
            .DOUT(N__9908),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__9910),
            .PADOUT(N__9909),
            .PADIN(N__9908),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4998),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__9901),
            .DIN(N__9900),
            .DOUT(N__9899),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__9901),
            .PADOUT(N__9900),
            .PADIN(N__9899),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7575),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__9892),
            .DIN(N__9891),
            .DOUT(N__9890),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__9892),
            .PADOUT(N__9891),
            .PADIN(N__9890),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__9883),
            .DIN(N__9882),
            .DOUT(N__9881),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__9883),
            .PADOUT(N__9882),
            .PADIN(N__9881),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_0_iopad (
            .OE(N__9874),
            .DIN(N__9873),
            .DOUT(N__9872),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__9874),
            .PADOUT(N__9873),
            .PADIN(N__9872),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__9865),
            .DIN(N__9864),
            .DOUT(N__9863),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__9865),
            .PADOUT(N__9864),
            .PADIN(N__9863),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5130),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__9856),
            .DIN(N__9855),
            .DOUT(N__9854),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__9856),
            .PADOUT(N__9855),
            .PADIN(N__9854),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__9847),
            .DIN(N__9846),
            .DOUT(N__9845),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__9847),
            .PADOUT(N__9846),
            .PADIN(N__9845),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8610),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__9838),
            .DIN(N__9837),
            .DOUT(N__9836),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__9838),
            .PADOUT(N__9837),
            .PADIN(N__9836),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6186),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__9829),
            .DIN(N__9828),
            .DOUT(N__9827),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__9829),
            .PADOUT(N__9828),
            .PADIN(N__9827),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7170),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__9820),
            .DIN(N__9819),
            .DOUT(N__9818),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__9820),
            .PADOUT(N__9819),
            .PADIN(N__9818),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7392),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__9811),
            .DIN(N__9810),
            .DOUT(N__9809),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__9811),
            .PADOUT(N__9810),
            .PADIN(N__9809),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4994),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__9802),
            .DIN(N__9801),
            .DOUT(N__9800),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__9802),
            .PADOUT(N__9801),
            .PADIN(N__9800),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__9793),
            .DIN(N__9792),
            .DOUT(N__9791),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__9793),
            .PADOUT(N__9792),
            .PADIN(N__9791),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__9784),
            .DIN(N__9783),
            .DOUT(N__9782),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__9784),
            .PADOUT(N__9783),
            .PADIN(N__9782),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6870),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__9775),
            .DIN(N__9774),
            .DOUT(N__9773),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__9775),
            .PADOUT(N__9774),
            .PADIN(N__9773),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7014),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__9766),
            .DIN(N__9765),
            .DOUT(N__9764),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__9766),
            .PADOUT(N__9765),
            .PADIN(N__9764),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6681),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_OUT_obuf_iopad (
            .OE(N__9757),
            .DIN(N__9756),
            .DOUT(N__9755),
            .PACKAGEPIN(CLK40_OUT));
    defparam CLK40_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40_OUT_obuf_preio (
            .PADOEN(N__9757),
            .PADOUT(N__9756),
            .PADIN(N__9755),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3693),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__9748),
            .DIN(N__9747),
            .DOUT(N__9746),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__9748),
            .PADOUT(N__9747),
            .PADIN(N__9746),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7116),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__9739),
            .DIN(N__9738),
            .DOUT(N__9737),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__9739),
            .PADOUT(N__9738),
            .PADIN(N__9737),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__9730),
            .DIN(N__9729),
            .DOUT(N__9728),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__9730),
            .PADOUT(N__9729),
            .PADIN(N__9728),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__9721),
            .DIN(N__9720),
            .DOUT(N__9719),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__9721),
            .PADOUT(N__9720),
            .PADIN(N__9719),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__9712),
            .DIN(N__9711),
            .DOUT(N__9710),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__9712),
            .PADOUT(N__9711),
            .PADIN(N__9710),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__9703),
            .DIN(N__9702),
            .DOUT(N__9701),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__9703),
            .PADOUT(N__9702),
            .PADIN(N__9701),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5772),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__9694),
            .DIN(N__9693),
            .DOUT(N__9692),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__9694),
            .PADOUT(N__9693),
            .PADIN(N__9692),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__9685),
            .DIN(N__9684),
            .DOUT(N__9683),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__9685),
            .PADOUT(N__9684),
            .PADIN(N__9683),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7287),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__9676),
            .DIN(N__9675),
            .DOUT(N__9674),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__9676),
            .PADOUT(N__9675),
            .PADIN(N__9674),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3678),
            .DIN0(),
            .DOUT0(N__6357),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__9667),
            .DIN(N__9666),
            .DOUT(N__9665),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__9667),
            .PADOUT(N__9666),
            .PADIN(N__9665),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6762),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__9658),
            .DIN(N__9657),
            .DOUT(N__9656),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__9658),
            .PADOUT(N__9657),
            .PADIN(N__9656),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__9649),
            .DIN(N__9648),
            .DOUT(N__9647),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__9649),
            .PADOUT(N__9648),
            .PADIN(N__9647),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__9640),
            .DIN(N__9639),
            .DOUT(N__9638),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__9640),
            .PADOUT(N__9639),
            .PADIN(N__9638),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7536),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__9631),
            .DIN(N__9630),
            .DOUT(N__9629),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__9631),
            .PADOUT(N__9630),
            .PADIN(N__9629),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__9622),
            .DIN(N__9621),
            .DOUT(N__9620),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__9622),
            .PADOUT(N__9621),
            .PADIN(N__9620),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__9613),
            .DIN(N__9612),
            .DOUT(N__9611),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__9613),
            .PADOUT(N__9612),
            .PADIN(N__9611),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__9604),
            .DIN(N__9603),
            .DOUT(N__9602),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__9604),
            .PADOUT(N__9603),
            .PADIN(N__9602),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__9595),
            .DIN(N__9594),
            .DOUT(N__9593),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__9595),
            .PADOUT(N__9594),
            .PADIN(N__9593),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5742),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__9586),
            .DIN(N__9585),
            .DOUT(N__9584),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__9586),
            .PADOUT(N__9585),
            .PADIN(N__9584),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6021),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2291 (
            .O(N__9567),
            .I(N__9564));
    LocalMux I__2290 (
            .O(N__9564),
            .I(N__9561));
    Span4Mux_v I__2289 (
            .O(N__9561),
            .I(N__9558));
    Odrv4 I__2288 (
            .O(N__9558),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2287 (
            .O(N__9555),
            .I(N__9552));
    LocalMux I__2286 (
            .O(N__9552),
            .I(N__9548));
    InMux I__2285 (
            .O(N__9551),
            .I(N__9545));
    Span4Mux_v I__2284 (
            .O(N__9548),
            .I(N__9542));
    LocalMux I__2283 (
            .O(N__9545),
            .I(N__9539));
    Span4Mux_v I__2282 (
            .O(N__9542),
            .I(N__9536));
    Sp12to4 I__2281 (
            .O(N__9539),
            .I(N__9533));
    Sp12to4 I__2280 (
            .O(N__9536),
            .I(N__9528));
    Span12Mux_v I__2279 (
            .O(N__9533),
            .I(N__9528));
    Span12Mux_h I__2278 (
            .O(N__9528),
            .I(N__9525));
    Odrv12 I__2277 (
            .O(N__9525),
            .I(DRA_c_7));
    CascadeMux I__2276 (
            .O(N__9522),
            .I(N__9519));
    InMux I__2275 (
            .O(N__9519),
            .I(N__9516));
    LocalMux I__2274 (
            .O(N__9516),
            .I(N__9513));
    Span4Mux_h I__2273 (
            .O(N__9513),
            .I(N__9510));
    Odrv4 I__2272 (
            .O(N__9510),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2271 (
            .O(N__9507),
            .I(N__9504));
    LocalMux I__2270 (
            .O(N__9504),
            .I(N__9495));
    ClkMux I__2269 (
            .O(N__9503),
            .I(N__9480));
    ClkMux I__2268 (
            .O(N__9502),
            .I(N__9480));
    ClkMux I__2267 (
            .O(N__9501),
            .I(N__9480));
    ClkMux I__2266 (
            .O(N__9500),
            .I(N__9480));
    ClkMux I__2265 (
            .O(N__9499),
            .I(N__9480));
    ClkMux I__2264 (
            .O(N__9498),
            .I(N__9480));
    Glb2LocalMux I__2263 (
            .O(N__9495),
            .I(N__9480));
    GlobalMux I__2262 (
            .O(N__9480),
            .I(N__9477));
    gio2CtrlBuf I__2261 (
            .O(N__9477),
            .I(C3_c_g));
    CEMux I__2260 (
            .O(N__9474),
            .I(N__9471));
    LocalMux I__2259 (
            .O(N__9471),
            .I(N__9464));
    CEMux I__2258 (
            .O(N__9470),
            .I(N__9461));
    CEMux I__2257 (
            .O(N__9469),
            .I(N__9458));
    CEMux I__2256 (
            .O(N__9468),
            .I(N__9455));
    CEMux I__2255 (
            .O(N__9467),
            .I(N__9452));
    Span4Mux_v I__2254 (
            .O(N__9464),
            .I(N__9446));
    LocalMux I__2253 (
            .O(N__9461),
            .I(N__9446));
    LocalMux I__2252 (
            .O(N__9458),
            .I(N__9443));
    LocalMux I__2251 (
            .O(N__9455),
            .I(N__9438));
    LocalMux I__2250 (
            .O(N__9452),
            .I(N__9438));
    CEMux I__2249 (
            .O(N__9451),
            .I(N__9435));
    Span4Mux_h I__2248 (
            .O(N__9446),
            .I(N__9430));
    Span4Mux_v I__2247 (
            .O(N__9443),
            .I(N__9430));
    Span4Mux_v I__2246 (
            .O(N__9438),
            .I(N__9427));
    LocalMux I__2245 (
            .O(N__9435),
            .I(N__9424));
    Odrv4 I__2244 (
            .O(N__9430),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ));
    Odrv4 I__2243 (
            .O(N__9427),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ));
    Odrv12 I__2242 (
            .O(N__9424),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ));
    InMux I__2241 (
            .O(N__9417),
            .I(N__9409));
    InMux I__2240 (
            .O(N__9416),
            .I(N__9406));
    InMux I__2239 (
            .O(N__9415),
            .I(N__9403));
    InMux I__2238 (
            .O(N__9414),
            .I(N__9400));
    InMux I__2237 (
            .O(N__9413),
            .I(N__9397));
    InMux I__2236 (
            .O(N__9412),
            .I(N__9394));
    LocalMux I__2235 (
            .O(N__9409),
            .I(N__9388));
    LocalMux I__2234 (
            .O(N__9406),
            .I(N__9382));
    LocalMux I__2233 (
            .O(N__9403),
            .I(N__9372));
    LocalMux I__2232 (
            .O(N__9400),
            .I(N__9360));
    LocalMux I__2231 (
            .O(N__9397),
            .I(N__9351));
    LocalMux I__2230 (
            .O(N__9394),
            .I(N__9342));
    SRMux I__2229 (
            .O(N__9393),
            .I(N__9246));
    SRMux I__2228 (
            .O(N__9392),
            .I(N__9246));
    SRMux I__2227 (
            .O(N__9391),
            .I(N__9246));
    Glb2LocalMux I__2226 (
            .O(N__9388),
            .I(N__9246));
    SRMux I__2225 (
            .O(N__9387),
            .I(N__9246));
    SRMux I__2224 (
            .O(N__9386),
            .I(N__9246));
    SRMux I__2223 (
            .O(N__9385),
            .I(N__9246));
    Glb2LocalMux I__2222 (
            .O(N__9382),
            .I(N__9246));
    SRMux I__2221 (
            .O(N__9381),
            .I(N__9246));
    SRMux I__2220 (
            .O(N__9380),
            .I(N__9246));
    SRMux I__2219 (
            .O(N__9379),
            .I(N__9246));
    SRMux I__2218 (
            .O(N__9378),
            .I(N__9246));
    SRMux I__2217 (
            .O(N__9377),
            .I(N__9246));
    SRMux I__2216 (
            .O(N__9376),
            .I(N__9246));
    SRMux I__2215 (
            .O(N__9375),
            .I(N__9246));
    Glb2LocalMux I__2214 (
            .O(N__9372),
            .I(N__9246));
    SRMux I__2213 (
            .O(N__9371),
            .I(N__9246));
    SRMux I__2212 (
            .O(N__9370),
            .I(N__9246));
    SRMux I__2211 (
            .O(N__9369),
            .I(N__9246));
    SRMux I__2210 (
            .O(N__9368),
            .I(N__9246));
    SRMux I__2209 (
            .O(N__9367),
            .I(N__9246));
    SRMux I__2208 (
            .O(N__9366),
            .I(N__9246));
    SRMux I__2207 (
            .O(N__9365),
            .I(N__9246));
    SRMux I__2206 (
            .O(N__9364),
            .I(N__9246));
    SRMux I__2205 (
            .O(N__9363),
            .I(N__9246));
    Glb2LocalMux I__2204 (
            .O(N__9360),
            .I(N__9246));
    SRMux I__2203 (
            .O(N__9359),
            .I(N__9246));
    SRMux I__2202 (
            .O(N__9358),
            .I(N__9246));
    SRMux I__2201 (
            .O(N__9357),
            .I(N__9246));
    SRMux I__2200 (
            .O(N__9356),
            .I(N__9246));
    SRMux I__2199 (
            .O(N__9355),
            .I(N__9246));
    SRMux I__2198 (
            .O(N__9354),
            .I(N__9246));
    Glb2LocalMux I__2197 (
            .O(N__9351),
            .I(N__9246));
    SRMux I__2196 (
            .O(N__9350),
            .I(N__9246));
    SRMux I__2195 (
            .O(N__9349),
            .I(N__9246));
    SRMux I__2194 (
            .O(N__9348),
            .I(N__9246));
    SRMux I__2193 (
            .O(N__9347),
            .I(N__9246));
    SRMux I__2192 (
            .O(N__9346),
            .I(N__9246));
    SRMux I__2191 (
            .O(N__9345),
            .I(N__9246));
    Glb2LocalMux I__2190 (
            .O(N__9342),
            .I(N__9246));
    SRMux I__2189 (
            .O(N__9341),
            .I(N__9246));
    SRMux I__2188 (
            .O(N__9340),
            .I(N__9246));
    SRMux I__2187 (
            .O(N__9339),
            .I(N__9246));
    SRMux I__2186 (
            .O(N__9338),
            .I(N__9246));
    SRMux I__2185 (
            .O(N__9337),
            .I(N__9246));
    GlobalMux I__2184 (
            .O(N__9246),
            .I(N__9243));
    gio2CtrlBuf I__2183 (
            .O(N__9243),
            .I(RESETn_c_i_g));
    InMux I__2182 (
            .O(N__9240),
            .I(N__9237));
    LocalMux I__2181 (
            .O(N__9237),
            .I(N__9234));
    Odrv12 I__2180 (
            .O(N__9234),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__2179 (
            .O(N__9231),
            .I(N__9228));
    LocalMux I__2178 (
            .O(N__9228),
            .I(N__9225));
    Odrv12 I__2177 (
            .O(N__9225),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2176 (
            .O(N__9222),
            .I(N__9219));
    LocalMux I__2175 (
            .O(N__9219),
            .I(N__9216));
    Odrv4 I__2174 (
            .O(N__9216),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2173 (
            .O(N__9213),
            .I(N__9209));
    InMux I__2172 (
            .O(N__9212),
            .I(N__9206));
    LocalMux I__2171 (
            .O(N__9209),
            .I(N__9203));
    LocalMux I__2170 (
            .O(N__9206),
            .I(N__9200));
    Span4Mux_h I__2169 (
            .O(N__9203),
            .I(N__9197));
    Span4Mux_v I__2168 (
            .O(N__9200),
            .I(N__9194));
    Sp12to4 I__2167 (
            .O(N__9197),
            .I(N__9191));
    Sp12to4 I__2166 (
            .O(N__9194),
            .I(N__9188));
    Span12Mux_v I__2165 (
            .O(N__9191),
            .I(N__9185));
    Span12Mux_h I__2164 (
            .O(N__9188),
            .I(N__9182));
    Span12Mux_h I__2163 (
            .O(N__9185),
            .I(N__9177));
    Span12Mux_v I__2162 (
            .O(N__9182),
            .I(N__9177));
    Odrv12 I__2161 (
            .O(N__9177),
            .I(DRA_c_4));
    InMux I__2160 (
            .O(N__9174),
            .I(N__9171));
    LocalMux I__2159 (
            .O(N__9171),
            .I(N__9168));
    Span4Mux_h I__2158 (
            .O(N__9168),
            .I(N__9165));
    Odrv4 I__2157 (
            .O(N__9165),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2156 (
            .O(N__9162),
            .I(N__9159));
    LocalMux I__2155 (
            .O(N__9159),
            .I(N__9156));
    Span4Mux_h I__2154 (
            .O(N__9156),
            .I(N__9153));
    Odrv4 I__2153 (
            .O(N__9153),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2152 (
            .O(N__9150),
            .I(N__9146));
    InMux I__2151 (
            .O(N__9149),
            .I(N__9143));
    LocalMux I__2150 (
            .O(N__9146),
            .I(N__9138));
    LocalMux I__2149 (
            .O(N__9143),
            .I(N__9138));
    Span12Mux_v I__2148 (
            .O(N__9138),
            .I(N__9135));
    Span12Mux_h I__2147 (
            .O(N__9135),
            .I(N__9132));
    Span12Mux_v I__2146 (
            .O(N__9132),
            .I(N__9129));
    Odrv12 I__2145 (
            .O(N__9129),
            .I(DRA_c_9));
    InMux I__2144 (
            .O(N__9126),
            .I(N__9123));
    LocalMux I__2143 (
            .O(N__9123),
            .I(N__9120));
    Odrv4 I__2142 (
            .O(N__9120),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__2141 (
            .O(N__9117),
            .I(N__9113));
    InMux I__2140 (
            .O(N__9116),
            .I(N__9110));
    LocalMux I__2139 (
            .O(N__9113),
            .I(N__9105));
    LocalMux I__2138 (
            .O(N__9110),
            .I(N__9105));
    Span12Mux_v I__2137 (
            .O(N__9105),
            .I(N__9102));
    Span12Mux_h I__2136 (
            .O(N__9102),
            .I(N__9099));
    Span12Mux_v I__2135 (
            .O(N__9099),
            .I(N__9096));
    Odrv12 I__2134 (
            .O(N__9096),
            .I(DRA_c_1));
    InMux I__2133 (
            .O(N__9093),
            .I(N__9090));
    LocalMux I__2132 (
            .O(N__9090),
            .I(N__9087));
    Odrv12 I__2131 (
            .O(N__9087),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    CEMux I__2130 (
            .O(N__9084),
            .I(N__9078));
    CEMux I__2129 (
            .O(N__9083),
            .I(N__9075));
    CEMux I__2128 (
            .O(N__9082),
            .I(N__9072));
    CEMux I__2127 (
            .O(N__9081),
            .I(N__9069));
    LocalMux I__2126 (
            .O(N__9078),
            .I(N__9066));
    LocalMux I__2125 (
            .O(N__9075),
            .I(N__9062));
    LocalMux I__2124 (
            .O(N__9072),
            .I(N__9059));
    LocalMux I__2123 (
            .O(N__9069),
            .I(N__9056));
    Span4Mux_v I__2122 (
            .O(N__9066),
            .I(N__9053));
    CEMux I__2121 (
            .O(N__9065),
            .I(N__9050));
    Span4Mux_h I__2120 (
            .O(N__9062),
            .I(N__9047));
    Span4Mux_v I__2119 (
            .O(N__9059),
            .I(N__9038));
    Span4Mux_v I__2118 (
            .O(N__9056),
            .I(N__9038));
    Span4Mux_v I__2117 (
            .O(N__9053),
            .I(N__9038));
    LocalMux I__2116 (
            .O(N__9050),
            .I(N__9038));
    Odrv4 I__2115 (
            .O(N__9047),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ));
    Odrv4 I__2114 (
            .O(N__9038),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ));
    InMux I__2113 (
            .O(N__9033),
            .I(N__9029));
    InMux I__2112 (
            .O(N__9032),
            .I(N__9026));
    LocalMux I__2111 (
            .O(N__9029),
            .I(N__9021));
    LocalMux I__2110 (
            .O(N__9026),
            .I(N__9021));
    Span4Mux_h I__2109 (
            .O(N__9021),
            .I(N__9018));
    Sp12to4 I__2108 (
            .O(N__9018),
            .I(N__9015));
    Span12Mux_v I__2107 (
            .O(N__9015),
            .I(N__9012));
    Odrv12 I__2106 (
            .O(N__9012),
            .I(DRA_c_5));
    InMux I__2105 (
            .O(N__9009),
            .I(N__9006));
    LocalMux I__2104 (
            .O(N__9006),
            .I(N__9003));
    Odrv4 I__2103 (
            .O(N__9003),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2102 (
            .O(N__9000),
            .I(N__8997));
    LocalMux I__2101 (
            .O(N__8997),
            .I(N__8993));
    InMux I__2100 (
            .O(N__8996),
            .I(N__8990));
    Span4Mux_h I__2099 (
            .O(N__8993),
            .I(N__8985));
    LocalMux I__2098 (
            .O(N__8990),
            .I(N__8985));
    Span4Mux_h I__2097 (
            .O(N__8985),
            .I(N__8982));
    Span4Mux_v I__2096 (
            .O(N__8982),
            .I(N__8979));
    Sp12to4 I__2095 (
            .O(N__8979),
            .I(N__8976));
    Odrv12 I__2094 (
            .O(N__8976),
            .I(DRA_c_8));
    InMux I__2093 (
            .O(N__8973),
            .I(N__8970));
    LocalMux I__2092 (
            .O(N__8970),
            .I(N__8967));
    Odrv4 I__2091 (
            .O(N__8967),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2090 (
            .O(N__8964),
            .I(N__8961));
    LocalMux I__2089 (
            .O(N__8961),
            .I(N__8958));
    Span4Mux_h I__2088 (
            .O(N__8958),
            .I(N__8955));
    Odrv4 I__2087 (
            .O(N__8955),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2086 (
            .O(N__8952),
            .I(N__8949));
    LocalMux I__2085 (
            .O(N__8949),
            .I(N__8945));
    InMux I__2084 (
            .O(N__8948),
            .I(N__8942));
    Span4Mux_v I__2083 (
            .O(N__8945),
            .I(N__8939));
    LocalMux I__2082 (
            .O(N__8942),
            .I(N__8936));
    Sp12to4 I__2081 (
            .O(N__8939),
            .I(N__8933));
    Span12Mux_h I__2080 (
            .O(N__8936),
            .I(N__8930));
    Span12Mux_h I__2079 (
            .O(N__8933),
            .I(N__8927));
    Odrv12 I__2078 (
            .O(N__8930),
            .I(RAS0n_c));
    Odrv12 I__2077 (
            .O(N__8927),
            .I(RAS0n_c));
    InMux I__2076 (
            .O(N__8922),
            .I(N__8919));
    LocalMux I__2075 (
            .O(N__8919),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    InMux I__2074 (
            .O(N__8916),
            .I(N__8913));
    LocalMux I__2073 (
            .O(N__8913),
            .I(N__8909));
    InMux I__2072 (
            .O(N__8912),
            .I(N__8906));
    Span4Mux_h I__2071 (
            .O(N__8909),
            .I(N__8901));
    LocalMux I__2070 (
            .O(N__8906),
            .I(N__8901));
    Sp12to4 I__2069 (
            .O(N__8901),
            .I(N__8898));
    Span12Mux_v I__2068 (
            .O(N__8898),
            .I(N__8895));
    Span12Mux_h I__2067 (
            .O(N__8895),
            .I(N__8892));
    Odrv12 I__2066 (
            .O(N__8892),
            .I(DRA_c_6));
    InMux I__2065 (
            .O(N__8889),
            .I(N__8883));
    InMux I__2064 (
            .O(N__8888),
            .I(N__8883));
    LocalMux I__2063 (
            .O(N__8883),
            .I(N__8880));
    Span4Mux_h I__2062 (
            .O(N__8880),
            .I(N__8877));
    Odrv4 I__2061 (
            .O(N__8877),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__2060 (
            .O(N__8874),
            .I(N__8871));
    LocalMux I__2059 (
            .O(N__8871),
            .I(N__8862));
    ClkMux I__2058 (
            .O(N__8870),
            .I(N__8847));
    ClkMux I__2057 (
            .O(N__8869),
            .I(N__8847));
    ClkMux I__2056 (
            .O(N__8868),
            .I(N__8847));
    ClkMux I__2055 (
            .O(N__8867),
            .I(N__8847));
    ClkMux I__2054 (
            .O(N__8866),
            .I(N__8847));
    ClkMux I__2053 (
            .O(N__8865),
            .I(N__8847));
    Glb2LocalMux I__2052 (
            .O(N__8862),
            .I(N__8847));
    GlobalMux I__2051 (
            .O(N__8847),
            .I(N__8844));
    gio2CtrlBuf I__2050 (
            .O(N__8844),
            .I(C1_c_g));
    InMux I__2049 (
            .O(N__8841),
            .I(N__8837));
    InMux I__2048 (
            .O(N__8840),
            .I(N__8833));
    LocalMux I__2047 (
            .O(N__8837),
            .I(N__8830));
    InMux I__2046 (
            .O(N__8836),
            .I(N__8827));
    LocalMux I__2045 (
            .O(N__8833),
            .I(N__8824));
    Span4Mux_h I__2044 (
            .O(N__8830),
            .I(N__8819));
    LocalMux I__2043 (
            .O(N__8827),
            .I(N__8819));
    Span4Mux_v I__2042 (
            .O(N__8824),
            .I(N__8816));
    Sp12to4 I__2041 (
            .O(N__8819),
            .I(N__8813));
    Sp12to4 I__2040 (
            .O(N__8816),
            .I(N__8810));
    Span12Mux_v I__2039 (
            .O(N__8813),
            .I(N__8807));
    Span12Mux_h I__2038 (
            .O(N__8810),
            .I(N__8804));
    Span12Mux_h I__2037 (
            .O(N__8807),
            .I(N__8801));
    Span12Mux_v I__2036 (
            .O(N__8804),
            .I(N__8798));
    Odrv12 I__2035 (
            .O(N__8801),
            .I(DBRn_c));
    Odrv12 I__2034 (
            .O(N__8798),
            .I(DBRn_c));
    InMux I__2033 (
            .O(N__8793),
            .I(N__8790));
    LocalMux I__2032 (
            .O(N__8790),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__2031 (
            .O(N__8787),
            .I(N__8784));
    LocalMux I__2030 (
            .O(N__8784),
            .I(N__8781));
    Odrv4 I__2029 (
            .O(N__8781),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__2028 (
            .O(N__8778),
            .I(N__8774));
    InMux I__2027 (
            .O(N__8777),
            .I(N__8771));
    LocalMux I__2026 (
            .O(N__8774),
            .I(N__8768));
    LocalMux I__2025 (
            .O(N__8771),
            .I(N__8765));
    Span12Mux_h I__2024 (
            .O(N__8768),
            .I(N__8762));
    Span12Mux_v I__2023 (
            .O(N__8765),
            .I(N__8759));
    Span12Mux_v I__2022 (
            .O(N__8762),
            .I(N__8754));
    Span12Mux_h I__2021 (
            .O(N__8759),
            .I(N__8754));
    Odrv12 I__2020 (
            .O(N__8754),
            .I(DRA_c_3));
    InMux I__2019 (
            .O(N__8751),
            .I(N__8748));
    LocalMux I__2018 (
            .O(N__8748),
            .I(N__8745));
    Odrv12 I__2017 (
            .O(N__8745),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    IoInMux I__2016 (
            .O(N__8742),
            .I(N__8739));
    LocalMux I__2015 (
            .O(N__8739),
            .I(N__8736));
    Span4Mux_s2_v I__2014 (
            .O(N__8736),
            .I(N__8733));
    Span4Mux_v I__2013 (
            .O(N__8733),
            .I(N__8730));
    Span4Mux_h I__2012 (
            .O(N__8730),
            .I(N__8727));
    Span4Mux_h I__2011 (
            .O(N__8727),
            .I(N__8724));
    Odrv4 I__2010 (
            .O(N__8724),
            .I(CASn_c));
    InMux I__2009 (
            .O(N__8721),
            .I(N__8715));
    CascadeMux I__2008 (
            .O(N__8720),
            .I(N__8712));
    CascadeMux I__2007 (
            .O(N__8719),
            .I(N__8709));
    InMux I__2006 (
            .O(N__8718),
            .I(N__8706));
    LocalMux I__2005 (
            .O(N__8715),
            .I(N__8703));
    InMux I__2004 (
            .O(N__8712),
            .I(N__8699));
    InMux I__2003 (
            .O(N__8709),
            .I(N__8696));
    LocalMux I__2002 (
            .O(N__8706),
            .I(N__8691));
    Span4Mux_h I__2001 (
            .O(N__8703),
            .I(N__8691));
    InMux I__2000 (
            .O(N__8702),
            .I(N__8688));
    LocalMux I__1999 (
            .O(N__8699),
            .I(N__8685));
    LocalMux I__1998 (
            .O(N__8696),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1997 (
            .O(N__8691),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1996 (
            .O(N__8688),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1995 (
            .O(N__8685),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1994 (
            .O(N__8676),
            .I(N__8673));
    LocalMux I__1993 (
            .O(N__8673),
            .I(N__8670));
    Span4Mux_s2_v I__1992 (
            .O(N__8670),
            .I(N__8667));
    Span4Mux_v I__1991 (
            .O(N__8667),
            .I(N__8664));
    Span4Mux_h I__1990 (
            .O(N__8664),
            .I(N__8661));
    Odrv4 I__1989 (
            .O(N__8661),
            .I(CRCSn_c));
    InMux I__1988 (
            .O(N__8658),
            .I(N__8655));
    LocalMux I__1987 (
            .O(N__8655),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__1986 (
            .O(N__8652),
            .I(N__8649));
    LocalMux I__1985 (
            .O(N__8649),
            .I(N__8646));
    Span4Mux_s3_v I__1984 (
            .O(N__8646),
            .I(N__8643));
    Span4Mux_h I__1983 (
            .O(N__8643),
            .I(N__8640));
    Odrv4 I__1982 (
            .O(N__8640),
            .I(CMA_c_0));
    InMux I__1981 (
            .O(N__8637),
            .I(N__8631));
    InMux I__1980 (
            .O(N__8636),
            .I(N__8631));
    LocalMux I__1979 (
            .O(N__8631),
            .I(N__8628));
    Span4Mux_h I__1978 (
            .O(N__8628),
            .I(N__8625));
    Odrv4 I__1977 (
            .O(N__8625),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__1976 (
            .O(N__8622),
            .I(N__8619));
    LocalMux I__1975 (
            .O(N__8619),
            .I(N__8616));
    Span4Mux_h I__1974 (
            .O(N__8616),
            .I(N__8613));
    Odrv4 I__1973 (
            .O(N__8613),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    IoInMux I__1972 (
            .O(N__8610),
            .I(N__8607));
    LocalMux I__1971 (
            .O(N__8607),
            .I(N__8604));
    IoSpan4Mux I__1970 (
            .O(N__8604),
            .I(N__8601));
    Sp12to4 I__1969 (
            .O(N__8601),
            .I(N__8598));
    Span12Mux_s7_v I__1968 (
            .O(N__8598),
            .I(N__8595));
    Span12Mux_h I__1967 (
            .O(N__8595),
            .I(N__8592));
    Odrv12 I__1966 (
            .O(N__8592),
            .I(CMA_c_4));
    CascadeMux I__1965 (
            .O(N__8589),
            .I(N__8585));
    CascadeMux I__1964 (
            .O(N__8588),
            .I(N__8580));
    InMux I__1963 (
            .O(N__8585),
            .I(N__8573));
    CascadeMux I__1962 (
            .O(N__8584),
            .I(N__8566));
    CascadeMux I__1961 (
            .O(N__8583),
            .I(N__8563));
    InMux I__1960 (
            .O(N__8580),
            .I(N__8559));
    InMux I__1959 (
            .O(N__8579),
            .I(N__8556));
    CascadeMux I__1958 (
            .O(N__8578),
            .I(N__8553));
    CascadeMux I__1957 (
            .O(N__8577),
            .I(N__8549));
    CascadeMux I__1956 (
            .O(N__8576),
            .I(N__8545));
    LocalMux I__1955 (
            .O(N__8573),
            .I(N__8540));
    InMux I__1954 (
            .O(N__8572),
            .I(N__8535));
    InMux I__1953 (
            .O(N__8571),
            .I(N__8532));
    InMux I__1952 (
            .O(N__8570),
            .I(N__8521));
    InMux I__1951 (
            .O(N__8569),
            .I(N__8521));
    InMux I__1950 (
            .O(N__8566),
            .I(N__8521));
    InMux I__1949 (
            .O(N__8563),
            .I(N__8521));
    InMux I__1948 (
            .O(N__8562),
            .I(N__8518));
    LocalMux I__1947 (
            .O(N__8559),
            .I(N__8512));
    LocalMux I__1946 (
            .O(N__8556),
            .I(N__8512));
    InMux I__1945 (
            .O(N__8553),
            .I(N__8509));
    InMux I__1944 (
            .O(N__8552),
            .I(N__8506));
    InMux I__1943 (
            .O(N__8549),
            .I(N__8497));
    InMux I__1942 (
            .O(N__8548),
            .I(N__8497));
    InMux I__1941 (
            .O(N__8545),
            .I(N__8497));
    InMux I__1940 (
            .O(N__8544),
            .I(N__8497));
    InMux I__1939 (
            .O(N__8543),
            .I(N__8493));
    Span4Mux_v I__1938 (
            .O(N__8540),
            .I(N__8490));
    InMux I__1937 (
            .O(N__8539),
            .I(N__8487));
    InMux I__1936 (
            .O(N__8538),
            .I(N__8484));
    LocalMux I__1935 (
            .O(N__8535),
            .I(N__8481));
    LocalMux I__1934 (
            .O(N__8532),
            .I(N__8478));
    InMux I__1933 (
            .O(N__8531),
            .I(N__8473));
    InMux I__1932 (
            .O(N__8530),
            .I(N__8473));
    LocalMux I__1931 (
            .O(N__8521),
            .I(N__8468));
    LocalMux I__1930 (
            .O(N__8518),
            .I(N__8468));
    InMux I__1929 (
            .O(N__8517),
            .I(N__8465));
    Span4Mux_h I__1928 (
            .O(N__8512),
            .I(N__8456));
    LocalMux I__1927 (
            .O(N__8509),
            .I(N__8456));
    LocalMux I__1926 (
            .O(N__8506),
            .I(N__8456));
    LocalMux I__1925 (
            .O(N__8497),
            .I(N__8456));
    InMux I__1924 (
            .O(N__8496),
            .I(N__8453));
    LocalMux I__1923 (
            .O(N__8493),
            .I(N__8444));
    Sp12to4 I__1922 (
            .O(N__8490),
            .I(N__8444));
    LocalMux I__1921 (
            .O(N__8487),
            .I(N__8444));
    LocalMux I__1920 (
            .O(N__8484),
            .I(N__8444));
    Span4Mux_v I__1919 (
            .O(N__8481),
            .I(N__8437));
    Span4Mux_h I__1918 (
            .O(N__8478),
            .I(N__8437));
    LocalMux I__1917 (
            .O(N__8473),
            .I(N__8437));
    Span4Mux_v I__1916 (
            .O(N__8468),
            .I(N__8432));
    LocalMux I__1915 (
            .O(N__8465),
            .I(N__8432));
    Span4Mux_h I__1914 (
            .O(N__8456),
            .I(N__8429));
    LocalMux I__1913 (
            .O(N__8453),
            .I(N__8424));
    Span12Mux_h I__1912 (
            .O(N__8444),
            .I(N__8424));
    Span4Mux_h I__1911 (
            .O(N__8437),
            .I(N__8421));
    Odrv4 I__1910 (
            .O(N__8432),
            .I(CPU_CYCLEm));
    Odrv4 I__1909 (
            .O(N__8429),
            .I(CPU_CYCLEm));
    Odrv12 I__1908 (
            .O(N__8424),
            .I(CPU_CYCLEm));
    Odrv4 I__1907 (
            .O(N__8421),
            .I(CPU_CYCLEm));
    InMux I__1906 (
            .O(N__8412),
            .I(N__8409));
    LocalMux I__1905 (
            .O(N__8409),
            .I(N__8406));
    Span4Mux_h I__1904 (
            .O(N__8406),
            .I(N__8403));
    Odrv4 I__1903 (
            .O(N__8403),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    CascadeMux I__1902 (
            .O(N__8400),
            .I(N__8395));
    InMux I__1901 (
            .O(N__8399),
            .I(N__8390));
    CascadeMux I__1900 (
            .O(N__8398),
            .I(N__8387));
    InMux I__1899 (
            .O(N__8395),
            .I(N__8382));
    InMux I__1898 (
            .O(N__8394),
            .I(N__8379));
    CascadeMux I__1897 (
            .O(N__8393),
            .I(N__8376));
    LocalMux I__1896 (
            .O(N__8390),
            .I(N__8373));
    InMux I__1895 (
            .O(N__8387),
            .I(N__8370));
    InMux I__1894 (
            .O(N__8386),
            .I(N__8365));
    InMux I__1893 (
            .O(N__8385),
            .I(N__8365));
    LocalMux I__1892 (
            .O(N__8382),
            .I(N__8361));
    LocalMux I__1891 (
            .O(N__8379),
            .I(N__8353));
    InMux I__1890 (
            .O(N__8376),
            .I(N__8350));
    Span4Mux_h I__1889 (
            .O(N__8373),
            .I(N__8343));
    LocalMux I__1888 (
            .O(N__8370),
            .I(N__8343));
    LocalMux I__1887 (
            .O(N__8365),
            .I(N__8343));
    CascadeMux I__1886 (
            .O(N__8364),
            .I(N__8331));
    Span4Mux_v I__1885 (
            .O(N__8361),
            .I(N__8327));
    InMux I__1884 (
            .O(N__8360),
            .I(N__8318));
    InMux I__1883 (
            .O(N__8359),
            .I(N__8318));
    InMux I__1882 (
            .O(N__8358),
            .I(N__8318));
    InMux I__1881 (
            .O(N__8357),
            .I(N__8318));
    InMux I__1880 (
            .O(N__8356),
            .I(N__8315));
    Span4Mux_h I__1879 (
            .O(N__8353),
            .I(N__8312));
    LocalMux I__1878 (
            .O(N__8350),
            .I(N__8307));
    Span4Mux_v I__1877 (
            .O(N__8343),
            .I(N__8307));
    InMux I__1876 (
            .O(N__8342),
            .I(N__8302));
    InMux I__1875 (
            .O(N__8341),
            .I(N__8302));
    InMux I__1874 (
            .O(N__8340),
            .I(N__8291));
    InMux I__1873 (
            .O(N__8339),
            .I(N__8291));
    InMux I__1872 (
            .O(N__8338),
            .I(N__8291));
    InMux I__1871 (
            .O(N__8337),
            .I(N__8291));
    InMux I__1870 (
            .O(N__8336),
            .I(N__8291));
    InMux I__1869 (
            .O(N__8335),
            .I(N__8282));
    InMux I__1868 (
            .O(N__8334),
            .I(N__8282));
    InMux I__1867 (
            .O(N__8331),
            .I(N__8282));
    InMux I__1866 (
            .O(N__8330),
            .I(N__8282));
    Sp12to4 I__1865 (
            .O(N__8327),
            .I(N__8275));
    LocalMux I__1864 (
            .O(N__8318),
            .I(N__8275));
    LocalMux I__1863 (
            .O(N__8315),
            .I(N__8275));
    Odrv4 I__1862 (
            .O(N__8312),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1861 (
            .O(N__8307),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1860 (
            .O(N__8302),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1859 (
            .O(N__8291),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1858 (
            .O(N__8282),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__1857 (
            .O(N__8275),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    CascadeMux I__1856 (
            .O(N__8262),
            .I(N__8259));
    InMux I__1855 (
            .O(N__8259),
            .I(N__8253));
    CascadeMux I__1854 (
            .O(N__8258),
            .I(N__8249));
    CascadeMux I__1853 (
            .O(N__8257),
            .I(N__8246));
    CascadeMux I__1852 (
            .O(N__8256),
            .I(N__8242));
    LocalMux I__1851 (
            .O(N__8253),
            .I(N__8239));
    InMux I__1850 (
            .O(N__8252),
            .I(N__8234));
    InMux I__1849 (
            .O(N__8249),
            .I(N__8234));
    InMux I__1848 (
            .O(N__8246),
            .I(N__8231));
    InMux I__1847 (
            .O(N__8245),
            .I(N__8226));
    InMux I__1846 (
            .O(N__8242),
            .I(N__8226));
    Span4Mux_v I__1845 (
            .O(N__8239),
            .I(N__8219));
    LocalMux I__1844 (
            .O(N__8234),
            .I(N__8219));
    LocalMux I__1843 (
            .O(N__8231),
            .I(N__8214));
    LocalMux I__1842 (
            .O(N__8226),
            .I(N__8214));
    CascadeMux I__1841 (
            .O(N__8225),
            .I(N__8211));
    InMux I__1840 (
            .O(N__8224),
            .I(N__8207));
    Span4Mux_h I__1839 (
            .O(N__8219),
            .I(N__8204));
    Span4Mux_v I__1838 (
            .O(N__8214),
            .I(N__8201));
    InMux I__1837 (
            .O(N__8211),
            .I(N__8196));
    InMux I__1836 (
            .O(N__8210),
            .I(N__8196));
    LocalMux I__1835 (
            .O(N__8207),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__1834 (
            .O(N__8204),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__1833 (
            .O(N__8201),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1832 (
            .O(N__8196),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    InMux I__1831 (
            .O(N__8187),
            .I(N__8179));
    InMux I__1830 (
            .O(N__8186),
            .I(N__8176));
    InMux I__1829 (
            .O(N__8185),
            .I(N__8173));
    InMux I__1828 (
            .O(N__8184),
            .I(N__8170));
    InMux I__1827 (
            .O(N__8183),
            .I(N__8167));
    InMux I__1826 (
            .O(N__8182),
            .I(N__8164));
    LocalMux I__1825 (
            .O(N__8179),
            .I(\U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1 ));
    LocalMux I__1824 (
            .O(N__8176),
            .I(\U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1 ));
    LocalMux I__1823 (
            .O(N__8173),
            .I(\U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1 ));
    LocalMux I__1822 (
            .O(N__8170),
            .I(\U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1 ));
    LocalMux I__1821 (
            .O(N__8167),
            .I(\U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1 ));
    LocalMux I__1820 (
            .O(N__8164),
            .I(\U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1 ));
    CascadeMux I__1819 (
            .O(N__8151),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_ ));
    IoInMux I__1818 (
            .O(N__8148),
            .I(N__8145));
    LocalMux I__1817 (
            .O(N__8145),
            .I(N__8142));
    IoSpan4Mux I__1816 (
            .O(N__8142),
            .I(N__8139));
    Span4Mux_s2_h I__1815 (
            .O(N__8139),
            .I(N__8136));
    Sp12to4 I__1814 (
            .O(N__8136),
            .I(N__8133));
    Span12Mux_h I__1813 (
            .O(N__8133),
            .I(N__8130));
    Odrv12 I__1812 (
            .O(N__8130),
            .I(CMA_c_7));
    InMux I__1811 (
            .O(N__8127),
            .I(N__8124));
    LocalMux I__1810 (
            .O(N__8124),
            .I(N__8096));
    ClkMux I__1809 (
            .O(N__8123),
            .I(N__8019));
    ClkMux I__1808 (
            .O(N__8122),
            .I(N__8019));
    ClkMux I__1807 (
            .O(N__8121),
            .I(N__8019));
    ClkMux I__1806 (
            .O(N__8120),
            .I(N__8019));
    ClkMux I__1805 (
            .O(N__8119),
            .I(N__8019));
    ClkMux I__1804 (
            .O(N__8118),
            .I(N__8019));
    ClkMux I__1803 (
            .O(N__8117),
            .I(N__8019));
    ClkMux I__1802 (
            .O(N__8116),
            .I(N__8019));
    ClkMux I__1801 (
            .O(N__8115),
            .I(N__8019));
    ClkMux I__1800 (
            .O(N__8114),
            .I(N__8019));
    ClkMux I__1799 (
            .O(N__8113),
            .I(N__8019));
    ClkMux I__1798 (
            .O(N__8112),
            .I(N__8019));
    ClkMux I__1797 (
            .O(N__8111),
            .I(N__8019));
    ClkMux I__1796 (
            .O(N__8110),
            .I(N__8019));
    ClkMux I__1795 (
            .O(N__8109),
            .I(N__8019));
    ClkMux I__1794 (
            .O(N__8108),
            .I(N__8019));
    ClkMux I__1793 (
            .O(N__8107),
            .I(N__8019));
    ClkMux I__1792 (
            .O(N__8106),
            .I(N__8019));
    ClkMux I__1791 (
            .O(N__8105),
            .I(N__8019));
    ClkMux I__1790 (
            .O(N__8104),
            .I(N__8019));
    ClkMux I__1789 (
            .O(N__8103),
            .I(N__8019));
    ClkMux I__1788 (
            .O(N__8102),
            .I(N__8019));
    ClkMux I__1787 (
            .O(N__8101),
            .I(N__8019));
    ClkMux I__1786 (
            .O(N__8100),
            .I(N__8019));
    ClkMux I__1785 (
            .O(N__8099),
            .I(N__8019));
    Glb2LocalMux I__1784 (
            .O(N__8096),
            .I(N__8019));
    ClkMux I__1783 (
            .O(N__8095),
            .I(N__8019));
    ClkMux I__1782 (
            .O(N__8094),
            .I(N__8019));
    ClkMux I__1781 (
            .O(N__8093),
            .I(N__8019));
    ClkMux I__1780 (
            .O(N__8092),
            .I(N__8019));
    ClkMux I__1779 (
            .O(N__8091),
            .I(N__8019));
    ClkMux I__1778 (
            .O(N__8090),
            .I(N__8019));
    ClkMux I__1777 (
            .O(N__8089),
            .I(N__8019));
    ClkMux I__1776 (
            .O(N__8088),
            .I(N__8019));
    GlobalMux I__1775 (
            .O(N__8019),
            .I(CLK80_PLL));
    CEMux I__1774 (
            .O(N__8016),
            .I(N__8012));
    CEMux I__1773 (
            .O(N__8015),
            .I(N__8009));
    LocalMux I__1772 (
            .O(N__8012),
            .I(N__8004));
    LocalMux I__1771 (
            .O(N__8009),
            .I(N__8001));
    CEMux I__1770 (
            .O(N__8008),
            .I(N__7997));
    CEMux I__1769 (
            .O(N__8007),
            .I(N__7994));
    Span4Mux_v I__1768 (
            .O(N__8004),
            .I(N__7989));
    Span4Mux_v I__1767 (
            .O(N__8001),
            .I(N__7989));
    CEMux I__1766 (
            .O(N__8000),
            .I(N__7986));
    LocalMux I__1765 (
            .O(N__7997),
            .I(N__7981));
    LocalMux I__1764 (
            .O(N__7994),
            .I(N__7978));
    Span4Mux_h I__1763 (
            .O(N__7989),
            .I(N__7973));
    LocalMux I__1762 (
            .O(N__7986),
            .I(N__7973));
    CEMux I__1761 (
            .O(N__7985),
            .I(N__7970));
    CEMux I__1760 (
            .O(N__7984),
            .I(N__7967));
    Span4Mux_v I__1759 (
            .O(N__7981),
            .I(N__7964));
    Span4Mux_h I__1758 (
            .O(N__7978),
            .I(N__7959));
    Span4Mux_h I__1757 (
            .O(N__7973),
            .I(N__7959));
    LocalMux I__1756 (
            .O(N__7970),
            .I(N__7954));
    LocalMux I__1755 (
            .O(N__7967),
            .I(N__7954));
    Odrv4 I__1754 (
            .O(N__7964),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__1753 (
            .O(N__7959),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__1752 (
            .O(N__7954),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    InMux I__1751 (
            .O(N__7947),
            .I(N__7944));
    LocalMux I__1750 (
            .O(N__7944),
            .I(N__7941));
    Span4Mux_v I__1749 (
            .O(N__7941),
            .I(N__7937));
    InMux I__1748 (
            .O(N__7940),
            .I(N__7934));
    Sp12to4 I__1747 (
            .O(N__7937),
            .I(N__7931));
    LocalMux I__1746 (
            .O(N__7934),
            .I(N__7928));
    Span12Mux_h I__1745 (
            .O(N__7931),
            .I(N__7925));
    Span12Mux_h I__1744 (
            .O(N__7928),
            .I(N__7922));
    Span12Mux_v I__1743 (
            .O(N__7925),
            .I(N__7919));
    Span12Mux_v I__1742 (
            .O(N__7922),
            .I(N__7916));
    Odrv12 I__1741 (
            .O(N__7919),
            .I(DRA_c_2));
    Odrv12 I__1740 (
            .O(N__7916),
            .I(DRA_c_2));
    InMux I__1739 (
            .O(N__7911),
            .I(N__7908));
    LocalMux I__1738 (
            .O(N__7908),
            .I(N__7905));
    Odrv4 I__1737 (
            .O(N__7905),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1736 (
            .O(N__7902),
            .I(N__7898));
    InMux I__1735 (
            .O(N__7901),
            .I(N__7895));
    LocalMux I__1734 (
            .O(N__7898),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    LocalMux I__1733 (
            .O(N__7895),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    InMux I__1732 (
            .O(N__7890),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__1731 (
            .O(N__7887),
            .I(N__7883));
    InMux I__1730 (
            .O(N__7886),
            .I(N__7880));
    LocalMux I__1729 (
            .O(N__7883),
            .I(N__7877));
    LocalMux I__1728 (
            .O(N__7880),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    Odrv4 I__1727 (
            .O(N__7877),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__1726 (
            .O(N__7872),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    CascadeMux I__1725 (
            .O(N__7869),
            .I(N__7865));
    InMux I__1724 (
            .O(N__7868),
            .I(N__7862));
    InMux I__1723 (
            .O(N__7865),
            .I(N__7859));
    LocalMux I__1722 (
            .O(N__7862),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__1721 (
            .O(N__7859),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__1720 (
            .O(N__7854),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__1719 (
            .O(N__7851),
            .I(N__7847));
    InMux I__1718 (
            .O(N__7850),
            .I(N__7844));
    LocalMux I__1717 (
            .O(N__7847),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__1716 (
            .O(N__7844),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__1715 (
            .O(N__7839),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__1714 (
            .O(N__7836),
            .I(N__7832));
    InMux I__1713 (
            .O(N__7835),
            .I(N__7829));
    LocalMux I__1712 (
            .O(N__7832),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__1711 (
            .O(N__7829),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__1710 (
            .O(N__7824),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__1709 (
            .O(N__7821),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    CascadeMux I__1708 (
            .O(N__7818),
            .I(N__7815));
    InMux I__1707 (
            .O(N__7815),
            .I(N__7811));
    InMux I__1706 (
            .O(N__7814),
            .I(N__7808));
    LocalMux I__1705 (
            .O(N__7811),
            .I(N__7805));
    LocalMux I__1704 (
            .O(N__7808),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv12 I__1703 (
            .O(N__7805),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    SRMux I__1702 (
            .O(N__7800),
            .I(N__7797));
    LocalMux I__1701 (
            .O(N__7797),
            .I(N__7794));
    Span4Mux_h I__1700 (
            .O(N__7794),
            .I(N__7791));
    Odrv4 I__1699 (
            .O(N__7791),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    CascadeMux I__1698 (
            .O(N__7788),
            .I(N__7785));
    InMux I__1697 (
            .O(N__7785),
            .I(N__7774));
    InMux I__1696 (
            .O(N__7784),
            .I(N__7774));
    InMux I__1695 (
            .O(N__7783),
            .I(N__7766));
    InMux I__1694 (
            .O(N__7782),
            .I(N__7766));
    InMux I__1693 (
            .O(N__7781),
            .I(N__7766));
    InMux I__1692 (
            .O(N__7780),
            .I(N__7761));
    InMux I__1691 (
            .O(N__7779),
            .I(N__7761));
    LocalMux I__1690 (
            .O(N__7774),
            .I(N__7756));
    InMux I__1689 (
            .O(N__7773),
            .I(N__7753));
    LocalMux I__1688 (
            .O(N__7766),
            .I(N__7750));
    LocalMux I__1687 (
            .O(N__7761),
            .I(N__7747));
    InMux I__1686 (
            .O(N__7760),
            .I(N__7742));
    InMux I__1685 (
            .O(N__7759),
            .I(N__7742));
    Span4Mux_v I__1684 (
            .O(N__7756),
            .I(N__7737));
    LocalMux I__1683 (
            .O(N__7753),
            .I(N__7737));
    Span4Mux_v I__1682 (
            .O(N__7750),
            .I(N__7734));
    Span4Mux_h I__1681 (
            .O(N__7747),
            .I(N__7729));
    LocalMux I__1680 (
            .O(N__7742),
            .I(N__7729));
    Span4Mux_v I__1679 (
            .O(N__7737),
            .I(N__7725));
    Span4Mux_v I__1678 (
            .O(N__7734),
            .I(N__7720));
    Span4Mux_v I__1677 (
            .O(N__7729),
            .I(N__7720));
    InMux I__1676 (
            .O(N__7728),
            .I(N__7717));
    Sp12to4 I__1675 (
            .O(N__7725),
            .I(N__7712));
    Sp12to4 I__1674 (
            .O(N__7720),
            .I(N__7712));
    LocalMux I__1673 (
            .O(N__7717),
            .I(N__7709));
    Span12Mux_h I__1672 (
            .O(N__7712),
            .I(N__7706));
    Span12Mux_h I__1671 (
            .O(N__7709),
            .I(N__7703));
    Odrv12 I__1670 (
            .O(N__7706),
            .I(RESETn_c));
    Odrv12 I__1669 (
            .O(N__7703),
            .I(RESETn_c));
    IoInMux I__1668 (
            .O(N__7698),
            .I(N__7695));
    LocalMux I__1667 (
            .O(N__7695),
            .I(N__7692));
    Span12Mux_s7_v I__1666 (
            .O(N__7692),
            .I(N__7689));
    Odrv12 I__1665 (
            .O(N__7689),
            .I(RESETn_c_i));
    InMux I__1664 (
            .O(N__7686),
            .I(N__7683));
    LocalMux I__1663 (
            .O(N__7683),
            .I(N__7678));
    InMux I__1662 (
            .O(N__7682),
            .I(N__7675));
    InMux I__1661 (
            .O(N__7681),
            .I(N__7668));
    Span4Mux_h I__1660 (
            .O(N__7678),
            .I(N__7663));
    LocalMux I__1659 (
            .O(N__7675),
            .I(N__7663));
    InMux I__1658 (
            .O(N__7674),
            .I(N__7660));
    InMux I__1657 (
            .O(N__7673),
            .I(N__7653));
    InMux I__1656 (
            .O(N__7672),
            .I(N__7653));
    InMux I__1655 (
            .O(N__7671),
            .I(N__7653));
    LocalMux I__1654 (
            .O(N__7668),
            .I(N__7650));
    Odrv4 I__1653 (
            .O(N__7663),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1652 (
            .O(N__7660),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1651 (
            .O(N__7653),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1650 (
            .O(N__7650),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__1649 (
            .O(N__7641),
            .I(N__7638));
    LocalMux I__1648 (
            .O(N__7638),
            .I(N__7635));
    Span12Mux_s6_v I__1647 (
            .O(N__7635),
            .I(N__7632));
    Odrv12 I__1646 (
            .O(N__7632),
            .I(RASn_c));
    CascadeMux I__1645 (
            .O(N__7629),
            .I(N__7626));
    InMux I__1644 (
            .O(N__7626),
            .I(N__7623));
    LocalMux I__1643 (
            .O(N__7623),
            .I(N__7620));
    Span4Mux_h I__1642 (
            .O(N__7620),
            .I(N__7617));
    Odrv4 I__1641 (
            .O(N__7617),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    InMux I__1640 (
            .O(N__7614),
            .I(N__7611));
    LocalMux I__1639 (
            .O(N__7611),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__1638 (
            .O(N__7608),
            .I(N__7605));
    LocalMux I__1637 (
            .O(N__7605),
            .I(N__7602));
    Span4Mux_s3_h I__1636 (
            .O(N__7602),
            .I(N__7599));
    Span4Mux_v I__1635 (
            .O(N__7599),
            .I(N__7596));
    Span4Mux_h I__1634 (
            .O(N__7596),
            .I(N__7593));
    Span4Mux_h I__1633 (
            .O(N__7593),
            .I(N__7590));
    Span4Mux_h I__1632 (
            .O(N__7590),
            .I(N__7587));
    Odrv4 I__1631 (
            .O(N__7587),
            .I(CMA_c_6));
    InMux I__1630 (
            .O(N__7584),
            .I(N__7581));
    LocalMux I__1629 (
            .O(N__7581),
            .I(N__7578));
    Odrv12 I__1628 (
            .O(N__7578),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__1627 (
            .O(N__7575),
            .I(N__7572));
    LocalMux I__1626 (
            .O(N__7572),
            .I(N__7569));
    IoSpan4Mux I__1625 (
            .O(N__7569),
            .I(N__7566));
    IoSpan4Mux I__1624 (
            .O(N__7566),
            .I(N__7563));
    Span4Mux_s2_h I__1623 (
            .O(N__7563),
            .I(N__7560));
    Sp12to4 I__1622 (
            .O(N__7560),
            .I(N__7557));
    Span12Mux_h I__1621 (
            .O(N__7557),
            .I(N__7554));
    Odrv12 I__1620 (
            .O(N__7554),
            .I(CMA_c_3));
    InMux I__1619 (
            .O(N__7551),
            .I(N__7548));
    LocalMux I__1618 (
            .O(N__7548),
            .I(N__7545));
    Span12Mux_v I__1617 (
            .O(N__7545),
            .I(N__7542));
    Span12Mux_h I__1616 (
            .O(N__7542),
            .I(N__7539));
    Odrv12 I__1615 (
            .O(N__7539),
            .I(A_c_17));
    IoInMux I__1614 (
            .O(N__7536),
            .I(N__7533));
    LocalMux I__1613 (
            .O(N__7533),
            .I(N__7530));
    Span4Mux_s3_h I__1612 (
            .O(N__7530),
            .I(N__7527));
    Span4Mux_v I__1611 (
            .O(N__7527),
            .I(N__7524));
    Span4Mux_h I__1610 (
            .O(N__7524),
            .I(N__7521));
    Span4Mux_h I__1609 (
            .O(N__7521),
            .I(N__7518));
    Span4Mux_h I__1608 (
            .O(N__7518),
            .I(N__7515));
    Odrv4 I__1607 (
            .O(N__7515),
            .I(CMA_c_8));
    CascadeMux I__1606 (
            .O(N__7512),
            .I(N__7509));
    InMux I__1605 (
            .O(N__7509),
            .I(N__7505));
    InMux I__1604 (
            .O(N__7508),
            .I(N__7501));
    LocalMux I__1603 (
            .O(N__7505),
            .I(N__7496));
    CascadeMux I__1602 (
            .O(N__7504),
            .I(N__7492));
    LocalMux I__1601 (
            .O(N__7501),
            .I(N__7489));
    InMux I__1600 (
            .O(N__7500),
            .I(N__7486));
    CascadeMux I__1599 (
            .O(N__7499),
            .I(N__7483));
    Span4Mux_h I__1598 (
            .O(N__7496),
            .I(N__7480));
    CascadeMux I__1597 (
            .O(N__7495),
            .I(N__7477));
    InMux I__1596 (
            .O(N__7492),
            .I(N__7473));
    Span4Mux_v I__1595 (
            .O(N__7489),
            .I(N__7468));
    LocalMux I__1594 (
            .O(N__7486),
            .I(N__7468));
    InMux I__1593 (
            .O(N__7483),
            .I(N__7465));
    Span4Mux_v I__1592 (
            .O(N__7480),
            .I(N__7462));
    InMux I__1591 (
            .O(N__7477),
            .I(N__7457));
    InMux I__1590 (
            .O(N__7476),
            .I(N__7457));
    LocalMux I__1589 (
            .O(N__7473),
            .I(N__7454));
    Span4Mux_h I__1588 (
            .O(N__7468),
            .I(N__7451));
    LocalMux I__1587 (
            .O(N__7465),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1586 (
            .O(N__7462),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1585 (
            .O(N__7457),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1584 (
            .O(N__7454),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1583 (
            .O(N__7451),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    InMux I__1582 (
            .O(N__7440),
            .I(N__7436));
    InMux I__1581 (
            .O(N__7439),
            .I(N__7433));
    LocalMux I__1580 (
            .O(N__7436),
            .I(N__7430));
    LocalMux I__1579 (
            .O(N__7433),
            .I(N__7427));
    Span4Mux_v I__1578 (
            .O(N__7430),
            .I(N__7422));
    Span4Mux_h I__1577 (
            .O(N__7427),
            .I(N__7419));
    InMux I__1576 (
            .O(N__7426),
            .I(N__7414));
    InMux I__1575 (
            .O(N__7425),
            .I(N__7414));
    Odrv4 I__1574 (
            .O(N__7422),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    Odrv4 I__1573 (
            .O(N__7419),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1572 (
            .O(N__7414),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    InMux I__1571 (
            .O(N__7407),
            .I(N__7404));
    LocalMux I__1570 (
            .O(N__7404),
            .I(N__7401));
    Span12Mux_v I__1569 (
            .O(N__7401),
            .I(N__7398));
    Span12Mux_h I__1568 (
            .O(N__7398),
            .I(N__7395));
    Odrv12 I__1567 (
            .O(N__7395),
            .I(A_c_19));
    IoInMux I__1566 (
            .O(N__7392),
            .I(N__7389));
    LocalMux I__1565 (
            .O(N__7389),
            .I(N__7386));
    Span4Mux_s3_h I__1564 (
            .O(N__7386),
            .I(N__7383));
    Span4Mux_v I__1563 (
            .O(N__7383),
            .I(N__7380));
    Span4Mux_h I__1562 (
            .O(N__7380),
            .I(N__7377));
    Span4Mux_h I__1561 (
            .O(N__7377),
            .I(N__7374));
    Span4Mux_h I__1560 (
            .O(N__7374),
            .I(N__7371));
    Odrv4 I__1559 (
            .O(N__7371),
            .I(CMA_c_9));
    InMux I__1558 (
            .O(N__7368),
            .I(N__7364));
    InMux I__1557 (
            .O(N__7367),
            .I(N__7361));
    LocalMux I__1556 (
            .O(N__7364),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    LocalMux I__1555 (
            .O(N__7361),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__1554 (
            .O(N__7356),
            .I(bfn_12_8_0_));
    InMux I__1553 (
            .O(N__7353),
            .I(N__7349));
    InMux I__1552 (
            .O(N__7352),
            .I(N__7346));
    LocalMux I__1551 (
            .O(N__7349),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    LocalMux I__1550 (
            .O(N__7346),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    InMux I__1549 (
            .O(N__7341),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    CascadeMux I__1548 (
            .O(N__7338),
            .I(N__7335));
    InMux I__1547 (
            .O(N__7335),
            .I(N__7330));
    InMux I__1546 (
            .O(N__7334),
            .I(N__7327));
    InMux I__1545 (
            .O(N__7333),
            .I(N__7324));
    LocalMux I__1544 (
            .O(N__7330),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__1543 (
            .O(N__7327),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__1542 (
            .O(N__7324),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__1541 (
            .O(N__7317),
            .I(N__7313));
    InMux I__1540 (
            .O(N__7316),
            .I(N__7310));
    LocalMux I__1539 (
            .O(N__7313),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    LocalMux I__1538 (
            .O(N__7310),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__1537 (
            .O(N__7305),
            .I(N__7302));
    LocalMux I__1536 (
            .O(N__7302),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ));
    InMux I__1535 (
            .O(N__7299),
            .I(N__7296));
    LocalMux I__1534 (
            .O(N__7296),
            .I(N__7293));
    Odrv4 I__1533 (
            .O(N__7293),
            .I(\U712_BYTE_ENABLE.N_271 ));
    CascadeMux I__1532 (
            .O(N__7290),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0_cascade_ ));
    IoInMux I__1531 (
            .O(N__7287),
            .I(N__7284));
    LocalMux I__1530 (
            .O(N__7284),
            .I(N__7281));
    IoSpan4Mux I__1529 (
            .O(N__7281),
            .I(N__7278));
    Span4Mux_s3_h I__1528 (
            .O(N__7278),
            .I(N__7275));
    Sp12to4 I__1527 (
            .O(N__7275),
            .I(N__7272));
    Span12Mux_h I__1526 (
            .O(N__7272),
            .I(N__7269));
    Odrv12 I__1525 (
            .O(N__7269),
            .I(N_171_i));
    IoInMux I__1524 (
            .O(N__7266),
            .I(N__7263));
    LocalMux I__1523 (
            .O(N__7263),
            .I(N__7260));
    Span4Mux_s1_v I__1522 (
            .O(N__7260),
            .I(N__7255));
    InMux I__1521 (
            .O(N__7259),
            .I(N__7250));
    InMux I__1520 (
            .O(N__7258),
            .I(N__7250));
    Sp12to4 I__1519 (
            .O(N__7255),
            .I(N__7247));
    LocalMux I__1518 (
            .O(N__7250),
            .I(N__7244));
    Span12Mux_h I__1517 (
            .O(N__7247),
            .I(N__7240));
    Span4Mux_v I__1516 (
            .O(N__7244),
            .I(N__7237));
    InMux I__1515 (
            .O(N__7243),
            .I(N__7234));
    Odrv12 I__1514 (
            .O(N__7240),
            .I(DBENn_c));
    Odrv4 I__1513 (
            .O(N__7237),
            .I(DBENn_c));
    LocalMux I__1512 (
            .O(N__7234),
            .I(DBENn_c));
    InMux I__1511 (
            .O(N__7227),
            .I(N__7223));
    InMux I__1510 (
            .O(N__7226),
            .I(N__7220));
    LocalMux I__1509 (
            .O(N__7223),
            .I(N__7213));
    LocalMux I__1508 (
            .O(N__7220),
            .I(N__7213));
    InMux I__1507 (
            .O(N__7219),
            .I(N__7208));
    InMux I__1506 (
            .O(N__7218),
            .I(N__7208));
    Span12Mux_v I__1505 (
            .O(N__7213),
            .I(N__7203));
    LocalMux I__1504 (
            .O(N__7208),
            .I(N__7200));
    InMux I__1503 (
            .O(N__7207),
            .I(N__7197));
    InMux I__1502 (
            .O(N__7206),
            .I(N__7194));
    Odrv12 I__1501 (
            .O(N__7203),
            .I(DMA_CYCLEm));
    Odrv4 I__1500 (
            .O(N__7200),
            .I(DMA_CYCLEm));
    LocalMux I__1499 (
            .O(N__7197),
            .I(DMA_CYCLEm));
    LocalMux I__1498 (
            .O(N__7194),
            .I(DMA_CYCLEm));
    InMux I__1497 (
            .O(N__7185),
            .I(N__7182));
    LocalMux I__1496 (
            .O(N__7182),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0 ));
    InMux I__1495 (
            .O(N__7179),
            .I(N__7176));
    LocalMux I__1494 (
            .O(N__7176),
            .I(\U712_BYTE_ENABLE.N_277 ));
    CascadeMux I__1493 (
            .O(N__7173),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0_cascade_ ));
    IoInMux I__1492 (
            .O(N__7170),
            .I(N__7167));
    LocalMux I__1491 (
            .O(N__7167),
            .I(N__7164));
    Span4Mux_s3_v I__1490 (
            .O(N__7164),
            .I(N__7161));
    Span4Mux_v I__1489 (
            .O(N__7161),
            .I(N__7158));
    Span4Mux_v I__1488 (
            .O(N__7158),
            .I(N__7155));
    Span4Mux_v I__1487 (
            .O(N__7155),
            .I(N__7152));
    Odrv4 I__1486 (
            .O(N__7152),
            .I(N_150_i));
    InMux I__1485 (
            .O(N__7149),
            .I(N__7143));
    InMux I__1484 (
            .O(N__7148),
            .I(N__7136));
    InMux I__1483 (
            .O(N__7147),
            .I(N__7136));
    InMux I__1482 (
            .O(N__7146),
            .I(N__7136));
    LocalMux I__1481 (
            .O(N__7143),
            .I(\U712_BYTE_ENABLE.N_270 ));
    LocalMux I__1480 (
            .O(N__7136),
            .I(\U712_BYTE_ENABLE.N_270 ));
    InMux I__1479 (
            .O(N__7131),
            .I(N__7128));
    LocalMux I__1478 (
            .O(N__7128),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0 ));
    CascadeMux I__1477 (
            .O(N__7125),
            .I(N__7122));
    InMux I__1476 (
            .O(N__7122),
            .I(N__7119));
    LocalMux I__1475 (
            .O(N__7119),
            .I(\U712_BYTE_ENABLE.N_273 ));
    IoInMux I__1474 (
            .O(N__7116),
            .I(N__7113));
    LocalMux I__1473 (
            .O(N__7113),
            .I(N__7110));
    IoSpan4Mux I__1472 (
            .O(N__7110),
            .I(N__7107));
    Span4Mux_s2_h I__1471 (
            .O(N__7107),
            .I(N__7104));
    Sp12to4 I__1470 (
            .O(N__7104),
            .I(N__7101));
    Span12Mux_h I__1469 (
            .O(N__7101),
            .I(N__7098));
    Span12Mux_v I__1468 (
            .O(N__7098),
            .I(N__7095));
    Odrv12 I__1467 (
            .O(N__7095),
            .I(N_172_i));
    InMux I__1466 (
            .O(N__7092),
            .I(N__7086));
    InMux I__1465 (
            .O(N__7091),
            .I(N__7086));
    LocalMux I__1464 (
            .O(N__7086),
            .I(N__7082));
    InMux I__1463 (
            .O(N__7085),
            .I(N__7079));
    Span4Mux_h I__1462 (
            .O(N__7082),
            .I(N__7074));
    LocalMux I__1461 (
            .O(N__7079),
            .I(N__7074));
    Sp12to4 I__1460 (
            .O(N__7074),
            .I(N__7071));
    Span12Mux_v I__1459 (
            .O(N__7071),
            .I(N__7068));
    Span12Mux_h I__1458 (
            .O(N__7068),
            .I(N__7065));
    Odrv12 I__1457 (
            .O(N__7065),
            .I(CASLn_c));
    CascadeMux I__1456 (
            .O(N__7062),
            .I(N__7058));
    InMux I__1455 (
            .O(N__7061),
            .I(N__7053));
    InMux I__1454 (
            .O(N__7058),
            .I(N__7053));
    LocalMux I__1453 (
            .O(N__7053),
            .I(N__7050));
    Span4Mux_v I__1452 (
            .O(N__7050),
            .I(N__7046));
    InMux I__1451 (
            .O(N__7049),
            .I(N__7043));
    Sp12to4 I__1450 (
            .O(N__7046),
            .I(N__7038));
    LocalMux I__1449 (
            .O(N__7043),
            .I(N__7038));
    Span12Mux_h I__1448 (
            .O(N__7038),
            .I(N__7035));
    Span12Mux_v I__1447 (
            .O(N__7035),
            .I(N__7032));
    Odrv12 I__1446 (
            .O(N__7032),
            .I(CASUn_c));
    InMux I__1445 (
            .O(N__7029),
            .I(N__7025));
    InMux I__1444 (
            .O(N__7028),
            .I(N__7022));
    LocalMux I__1443 (
            .O(N__7025),
            .I(N__7017));
    LocalMux I__1442 (
            .O(N__7022),
            .I(N__7017));
    Odrv4 I__1441 (
            .O(N__7017),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    IoInMux I__1440 (
            .O(N__7014),
            .I(N__7011));
    LocalMux I__1439 (
            .O(N__7011),
            .I(N__7008));
    Span12Mux_s4_h I__1438 (
            .O(N__7008),
            .I(N__7005));
    Span12Mux_h I__1437 (
            .O(N__7005),
            .I(N__7002));
    Odrv12 I__1436 (
            .O(N__7002),
            .I(WEn_c));
    InMux I__1435 (
            .O(N__6999),
            .I(N__6996));
    LocalMux I__1434 (
            .O(N__6996),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ));
    InMux I__1433 (
            .O(N__6993),
            .I(N__6990));
    LocalMux I__1432 (
            .O(N__6990),
            .I(\U712_CHIP_RAM.un5_DMA_CYCLE_START_0 ));
    InMux I__1431 (
            .O(N__6987),
            .I(N__6984));
    LocalMux I__1430 (
            .O(N__6984),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    InMux I__1429 (
            .O(N__6981),
            .I(N__6973));
    InMux I__1428 (
            .O(N__6980),
            .I(N__6973));
    InMux I__1427 (
            .O(N__6979),
            .I(N__6970));
    InMux I__1426 (
            .O(N__6978),
            .I(N__6967));
    LocalMux I__1425 (
            .O(N__6973),
            .I(N__6962));
    LocalMux I__1424 (
            .O(N__6970),
            .I(N__6962));
    LocalMux I__1423 (
            .O(N__6967),
            .I(N__6959));
    Span4Mux_h I__1422 (
            .O(N__6962),
            .I(N__6956));
    Span12Mux_v I__1421 (
            .O(N__6959),
            .I(N__6953));
    Sp12to4 I__1420 (
            .O(N__6956),
            .I(N__6950));
    Span12Mux_h I__1419 (
            .O(N__6953),
            .I(N__6945));
    Span12Mux_v I__1418 (
            .O(N__6950),
            .I(N__6945));
    Odrv12 I__1417 (
            .O(N__6945),
            .I(CLK40_PLL_i));
    InMux I__1416 (
            .O(N__6942),
            .I(N__6936));
    InMux I__1415 (
            .O(N__6941),
            .I(N__6929));
    InMux I__1414 (
            .O(N__6940),
            .I(N__6929));
    InMux I__1413 (
            .O(N__6939),
            .I(N__6929));
    LocalMux I__1412 (
            .O(N__6936),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1411 (
            .O(N__6929),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__1410 (
            .O(N__6924),
            .I(N__6920));
    InMux I__1409 (
            .O(N__6923),
            .I(N__6917));
    LocalMux I__1408 (
            .O(N__6920),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__1407 (
            .O(N__6917),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    CascadeMux I__1406 (
            .O(N__6912),
            .I(N__6909));
    InMux I__1405 (
            .O(N__6909),
            .I(N__6906));
    LocalMux I__1404 (
            .O(N__6906),
            .I(N__6903));
    Odrv4 I__1403 (
            .O(N__6903),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_2 ));
    CascadeMux I__1402 (
            .O(N__6900),
            .I(N__6896));
    CascadeMux I__1401 (
            .O(N__6899),
            .I(N__6893));
    InMux I__1400 (
            .O(N__6896),
            .I(N__6890));
    InMux I__1399 (
            .O(N__6893),
            .I(N__6887));
    LocalMux I__1398 (
            .O(N__6890),
            .I(N__6884));
    LocalMux I__1397 (
            .O(N__6887),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    Odrv12 I__1396 (
            .O(N__6884),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    InMux I__1395 (
            .O(N__6879),
            .I(N__6876));
    LocalMux I__1394 (
            .O(N__6876),
            .I(N__6873));
    Odrv12 I__1393 (
            .O(N__6873),
            .I(\U712_BYTE_ENABLE.N_275 ));
    IoInMux I__1392 (
            .O(N__6870),
            .I(N__6867));
    LocalMux I__1391 (
            .O(N__6867),
            .I(N__6864));
    Span4Mux_s1_h I__1390 (
            .O(N__6864),
            .I(N__6861));
    Span4Mux_h I__1389 (
            .O(N__6861),
            .I(N__6858));
    Sp12to4 I__1388 (
            .O(N__6858),
            .I(N__6855));
    Span12Mux_s11_v I__1387 (
            .O(N__6855),
            .I(N__6852));
    Span12Mux_h I__1386 (
            .O(N__6852),
            .I(N__6849));
    Odrv12 I__1385 (
            .O(N__6849),
            .I(N_148_i));
    InMux I__1384 (
            .O(N__6846),
            .I(N__6843));
    LocalMux I__1383 (
            .O(N__6843),
            .I(N__6839));
    InMux I__1382 (
            .O(N__6842),
            .I(N__6836));
    Span4Mux_v I__1381 (
            .O(N__6839),
            .I(N__6833));
    LocalMux I__1380 (
            .O(N__6836),
            .I(N__6830));
    Sp12to4 I__1379 (
            .O(N__6833),
            .I(N__6827));
    Sp12to4 I__1378 (
            .O(N__6830),
            .I(N__6824));
    Span12Mux_h I__1377 (
            .O(N__6827),
            .I(N__6821));
    Span12Mux_v I__1376 (
            .O(N__6824),
            .I(N__6818));
    Span12Mux_v I__1375 (
            .O(N__6821),
            .I(N__6813));
    Span12Mux_h I__1374 (
            .O(N__6818),
            .I(N__6813));
    Odrv12 I__1373 (
            .O(N__6813),
            .I(RnW_c));
    IoInMux I__1372 (
            .O(N__6810),
            .I(N__6807));
    LocalMux I__1371 (
            .O(N__6807),
            .I(N__6804));
    Span4Mux_s1_h I__1370 (
            .O(N__6804),
            .I(N__6801));
    Sp12to4 I__1369 (
            .O(N__6801),
            .I(N__6798));
    Span12Mux_s8_v I__1368 (
            .O(N__6798),
            .I(N__6795));
    Span12Mux_h I__1367 (
            .O(N__6795),
            .I(N__6792));
    Odrv12 I__1366 (
            .O(N__6792),
            .I(N_212));
    IoInMux I__1365 (
            .O(N__6789),
            .I(N__6786));
    LocalMux I__1364 (
            .O(N__6786),
            .I(N__6782));
    InMux I__1363 (
            .O(N__6785),
            .I(N__6779));
    Span4Mux_s3_v I__1362 (
            .O(N__6782),
            .I(N__6776));
    LocalMux I__1361 (
            .O(N__6779),
            .I(N__6773));
    Span4Mux_h I__1360 (
            .O(N__6776),
            .I(N__6770));
    Span4Mux_v I__1359 (
            .O(N__6773),
            .I(N__6767));
    Odrv4 I__1358 (
            .O(N__6770),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1357 (
            .O(N__6767),
            .I(CONSTANT_ONE_NET));
    IoInMux I__1356 (
            .O(N__6762),
            .I(N__6759));
    LocalMux I__1355 (
            .O(N__6759),
            .I(N__6756));
    Span12Mux_s2_v I__1354 (
            .O(N__6756),
            .I(N__6753));
    Odrv12 I__1353 (
            .O(N__6753),
            .I(CMA_c_2));
    InMux I__1352 (
            .O(N__6750),
            .I(N__6747));
    LocalMux I__1351 (
            .O(N__6747),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    InMux I__1350 (
            .O(N__6744),
            .I(N__6741));
    LocalMux I__1349 (
            .O(N__6741),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    InMux I__1348 (
            .O(N__6738),
            .I(N__6735));
    LocalMux I__1347 (
            .O(N__6735),
            .I(N__6732));
    Odrv4 I__1346 (
            .O(N__6732),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    InMux I__1345 (
            .O(N__6729),
            .I(N__6726));
    LocalMux I__1344 (
            .O(N__6726),
            .I(N__6723));
    Span4Mux_v I__1343 (
            .O(N__6723),
            .I(N__6718));
    InMux I__1342 (
            .O(N__6722),
            .I(N__6715));
    InMux I__1341 (
            .O(N__6721),
            .I(N__6712));
    Span4Mux_h I__1340 (
            .O(N__6718),
            .I(N__6707));
    LocalMux I__1339 (
            .O(N__6715),
            .I(N__6707));
    LocalMux I__1338 (
            .O(N__6712),
            .I(N__6704));
    Span4Mux_v I__1337 (
            .O(N__6707),
            .I(N__6701));
    Span4Mux_v I__1336 (
            .O(N__6704),
            .I(N__6698));
    Span4Mux_h I__1335 (
            .O(N__6701),
            .I(N__6695));
    Sp12to4 I__1334 (
            .O(N__6698),
            .I(N__6692));
    Sp12to4 I__1333 (
            .O(N__6695),
            .I(N__6689));
    Span12Mux_h I__1332 (
            .O(N__6692),
            .I(N__6686));
    Odrv12 I__1331 (
            .O(N__6689),
            .I(AWEn_c));
    Odrv12 I__1330 (
            .O(N__6686),
            .I(AWEn_c));
    IoInMux I__1329 (
            .O(N__6681),
            .I(N__6678));
    LocalMux I__1328 (
            .O(N__6678),
            .I(N__6675));
    Span4Mux_s3_v I__1327 (
            .O(N__6675),
            .I(N__6672));
    Span4Mux_v I__1326 (
            .O(N__6672),
            .I(N__6669));
    Span4Mux_h I__1325 (
            .O(N__6669),
            .I(N__6665));
    InMux I__1324 (
            .O(N__6668),
            .I(N__6662));
    Odrv4 I__1323 (
            .O(N__6665),
            .I(DBDIR_c));
    LocalMux I__1322 (
            .O(N__6662),
            .I(DBDIR_c));
    InMux I__1321 (
            .O(N__6657),
            .I(N__6654));
    LocalMux I__1320 (
            .O(N__6654),
            .I(N__6651));
    Span4Mux_h I__1319 (
            .O(N__6651),
            .I(N__6647));
    InMux I__1318 (
            .O(N__6650),
            .I(N__6644));
    Odrv4 I__1317 (
            .O(N__6647),
            .I(\U712_CHIP_RAM.N_298 ));
    LocalMux I__1316 (
            .O(N__6644),
            .I(\U712_CHIP_RAM.N_298 ));
    CascadeMux I__1315 (
            .O(N__6639),
            .I(N__6632));
    CascadeMux I__1314 (
            .O(N__6638),
            .I(N__6628));
    InMux I__1313 (
            .O(N__6637),
            .I(N__6625));
    InMux I__1312 (
            .O(N__6636),
            .I(N__6622));
    InMux I__1311 (
            .O(N__6635),
            .I(N__6619));
    InMux I__1310 (
            .O(N__6632),
            .I(N__6616));
    InMux I__1309 (
            .O(N__6631),
            .I(N__6609));
    InMux I__1308 (
            .O(N__6628),
            .I(N__6609));
    LocalMux I__1307 (
            .O(N__6625),
            .I(N__6601));
    LocalMux I__1306 (
            .O(N__6622),
            .I(N__6601));
    LocalMux I__1305 (
            .O(N__6619),
            .I(N__6601));
    LocalMux I__1304 (
            .O(N__6616),
            .I(N__6598));
    InMux I__1303 (
            .O(N__6615),
            .I(N__6595));
    InMux I__1302 (
            .O(N__6614),
            .I(N__6589));
    LocalMux I__1301 (
            .O(N__6609),
            .I(N__6586));
    InMux I__1300 (
            .O(N__6608),
            .I(N__6583));
    Span4Mux_v I__1299 (
            .O(N__6601),
            .I(N__6580));
    Span4Mux_h I__1298 (
            .O(N__6598),
            .I(N__6575));
    LocalMux I__1297 (
            .O(N__6595),
            .I(N__6575));
    InMux I__1296 (
            .O(N__6594),
            .I(N__6568));
    InMux I__1295 (
            .O(N__6593),
            .I(N__6568));
    InMux I__1294 (
            .O(N__6592),
            .I(N__6568));
    LocalMux I__1293 (
            .O(N__6589),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv12 I__1292 (
            .O(N__6586),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1291 (
            .O(N__6583),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1290 (
            .O(N__6580),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1289 (
            .O(N__6575),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1288 (
            .O(N__6568),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__1287 (
            .O(N__6555),
            .I(N__6552));
    LocalMux I__1286 (
            .O(N__6552),
            .I(N__6546));
    InMux I__1285 (
            .O(N__6551),
            .I(N__6543));
    InMux I__1284 (
            .O(N__6550),
            .I(N__6539));
    InMux I__1283 (
            .O(N__6549),
            .I(N__6536));
    Span4Mux_v I__1282 (
            .O(N__6546),
            .I(N__6529));
    LocalMux I__1281 (
            .O(N__6543),
            .I(N__6529));
    InMux I__1280 (
            .O(N__6542),
            .I(N__6526));
    LocalMux I__1279 (
            .O(N__6539),
            .I(N__6523));
    LocalMux I__1278 (
            .O(N__6536),
            .I(N__6520));
    InMux I__1277 (
            .O(N__6535),
            .I(N__6515));
    InMux I__1276 (
            .O(N__6534),
            .I(N__6515));
    Odrv4 I__1275 (
            .O(N__6529),
            .I(\U712_CHIP_RAM.N_355 ));
    LocalMux I__1274 (
            .O(N__6526),
            .I(\U712_CHIP_RAM.N_355 ));
    Odrv4 I__1273 (
            .O(N__6523),
            .I(\U712_CHIP_RAM.N_355 ));
    Odrv4 I__1272 (
            .O(N__6520),
            .I(\U712_CHIP_RAM.N_355 ));
    LocalMux I__1271 (
            .O(N__6515),
            .I(\U712_CHIP_RAM.N_355 ));
    CascadeMux I__1270 (
            .O(N__6504),
            .I(N__6499));
    InMux I__1269 (
            .O(N__6503),
            .I(N__6496));
    InMux I__1268 (
            .O(N__6502),
            .I(N__6491));
    InMux I__1267 (
            .O(N__6499),
            .I(N__6491));
    LocalMux I__1266 (
            .O(N__6496),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    LocalMux I__1265 (
            .O(N__6491),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    InMux I__1264 (
            .O(N__6486),
            .I(N__6481));
    InMux I__1263 (
            .O(N__6485),
            .I(N__6478));
    InMux I__1262 (
            .O(N__6484),
            .I(N__6475));
    LocalMux I__1261 (
            .O(N__6481),
            .I(N__6472));
    LocalMux I__1260 (
            .O(N__6478),
            .I(N__6469));
    LocalMux I__1259 (
            .O(N__6475),
            .I(N__6465));
    Span4Mux_h I__1258 (
            .O(N__6472),
            .I(N__6462));
    Span4Mux_h I__1257 (
            .O(N__6469),
            .I(N__6459));
    InMux I__1256 (
            .O(N__6468),
            .I(N__6456));
    Odrv12 I__1255 (
            .O(N__6465),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__1254 (
            .O(N__6462),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__1253 (
            .O(N__6459),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1252 (
            .O(N__6456),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    CascadeMux I__1251 (
            .O(N__6447),
            .I(N__6444));
    InMux I__1250 (
            .O(N__6444),
            .I(N__6440));
    InMux I__1249 (
            .O(N__6443),
            .I(N__6435));
    LocalMux I__1248 (
            .O(N__6440),
            .I(N__6432));
    InMux I__1247 (
            .O(N__6439),
            .I(N__6429));
    InMux I__1246 (
            .O(N__6438),
            .I(N__6426));
    LocalMux I__1245 (
            .O(N__6435),
            .I(N__6423));
    Span4Mux_v I__1244 (
            .O(N__6432),
            .I(N__6418));
    LocalMux I__1243 (
            .O(N__6429),
            .I(N__6418));
    LocalMux I__1242 (
            .O(N__6426),
            .I(N__6415));
    Span4Mux_h I__1241 (
            .O(N__6423),
            .I(N__6409));
    Span4Mux_h I__1240 (
            .O(N__6418),
            .I(N__6404));
    Span4Mux_h I__1239 (
            .O(N__6415),
            .I(N__6404));
    InMux I__1238 (
            .O(N__6414),
            .I(N__6397));
    InMux I__1237 (
            .O(N__6413),
            .I(N__6397));
    InMux I__1236 (
            .O(N__6412),
            .I(N__6397));
    Odrv4 I__1235 (
            .O(N__6409),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1234 (
            .O(N__6404),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1233 (
            .O(N__6397),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1232 (
            .O(N__6390),
            .I(N__6387));
    LocalMux I__1231 (
            .O(N__6387),
            .I(N__6381));
    InMux I__1230 (
            .O(N__6386),
            .I(N__6378));
    InMux I__1229 (
            .O(N__6385),
            .I(N__6373));
    InMux I__1228 (
            .O(N__6384),
            .I(N__6373));
    Span4Mux_v I__1227 (
            .O(N__6381),
            .I(N__6368));
    LocalMux I__1226 (
            .O(N__6378),
            .I(N__6368));
    LocalMux I__1225 (
            .O(N__6373),
            .I(N__6365));
    Span4Mux_h I__1224 (
            .O(N__6368),
            .I(N__6362));
    Odrv12 I__1223 (
            .O(N__6365),
            .I(\U712_CHIP_RAM.N_305 ));
    Odrv4 I__1222 (
            .O(N__6362),
            .I(\U712_CHIP_RAM.N_305 ));
    IoInMux I__1221 (
            .O(N__6357),
            .I(N__6354));
    LocalMux I__1220 (
            .O(N__6354),
            .I(N__6351));
    Span12Mux_s1_h I__1219 (
            .O(N__6351),
            .I(N__6348));
    Span12Mux_v I__1218 (
            .O(N__6348),
            .I(N__6345));
    Span12Mux_h I__1217 (
            .O(N__6345),
            .I(N__6341));
    InMux I__1216 (
            .O(N__6344),
            .I(N__6338));
    Odrv12 I__1215 (
            .O(N__6341),
            .I(TACK_OUTn));
    LocalMux I__1214 (
            .O(N__6338),
            .I(TACK_OUTn));
    InMux I__1213 (
            .O(N__6333),
            .I(N__6327));
    InMux I__1212 (
            .O(N__6332),
            .I(N__6327));
    LocalMux I__1211 (
            .O(N__6327),
            .I(N__6322));
    InMux I__1210 (
            .O(N__6326),
            .I(N__6317));
    InMux I__1209 (
            .O(N__6325),
            .I(N__6317));
    Span4Mux_v I__1208 (
            .O(N__6322),
            .I(N__6314));
    LocalMux I__1207 (
            .O(N__6317),
            .I(N__6311));
    Odrv4 I__1206 (
            .O(N__6314),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    Odrv4 I__1205 (
            .O(N__6311),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CascadeMux I__1204 (
            .O(N__6306),
            .I(N__6301));
    InMux I__1203 (
            .O(N__6305),
            .I(N__6296));
    InMux I__1202 (
            .O(N__6304),
            .I(N__6296));
    InMux I__1201 (
            .O(N__6301),
            .I(N__6293));
    LocalMux I__1200 (
            .O(N__6296),
            .I(N__6290));
    LocalMux I__1199 (
            .O(N__6293),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    Odrv12 I__1198 (
            .O(N__6290),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__1197 (
            .O(N__6285),
            .I(N__6276));
    InMux I__1196 (
            .O(N__6284),
            .I(N__6276));
    InMux I__1195 (
            .O(N__6283),
            .I(N__6276));
    LocalMux I__1194 (
            .O(N__6276),
            .I(N__6273));
    Span4Mux_v I__1193 (
            .O(N__6273),
            .I(N__6270));
    Span4Mux_v I__1192 (
            .O(N__6270),
            .I(N__6266));
    InMux I__1191 (
            .O(N__6269),
            .I(N__6263));
    Span4Mux_v I__1190 (
            .O(N__6266),
            .I(N__6260));
    LocalMux I__1189 (
            .O(N__6263),
            .I(N__6257));
    Span4Mux_h I__1188 (
            .O(N__6260),
            .I(N__6254));
    Sp12to4 I__1187 (
            .O(N__6257),
            .I(N__6251));
    Sp12to4 I__1186 (
            .O(N__6254),
            .I(N__6246));
    Span12Mux_v I__1185 (
            .O(N__6251),
            .I(N__6246));
    Odrv12 I__1184 (
            .O(N__6246),
            .I(A_c_1));
    InMux I__1183 (
            .O(N__6243),
            .I(N__6234));
    InMux I__1182 (
            .O(N__6242),
            .I(N__6234));
    InMux I__1181 (
            .O(N__6241),
            .I(N__6234));
    LocalMux I__1180 (
            .O(N__6234),
            .I(N__6231));
    Span4Mux_v I__1179 (
            .O(N__6231),
            .I(N__6228));
    Sp12to4 I__1178 (
            .O(N__6228),
            .I(N__6225));
    Span12Mux_v I__1177 (
            .O(N__6225),
            .I(N__6222));
    Span12Mux_h I__1176 (
            .O(N__6222),
            .I(N__6219));
    Odrv12 I__1175 (
            .O(N__6219),
            .I(SIZ_c_1));
    InMux I__1174 (
            .O(N__6216),
            .I(N__6213));
    LocalMux I__1173 (
            .O(N__6213),
            .I(N__6209));
    InMux I__1172 (
            .O(N__6212),
            .I(N__6206));
    Span4Mux_h I__1171 (
            .O(N__6209),
            .I(N__6203));
    LocalMux I__1170 (
            .O(N__6206),
            .I(N__6200));
    Span4Mux_v I__1169 (
            .O(N__6203),
            .I(N__6194));
    Span4Mux_v I__1168 (
            .O(N__6200),
            .I(N__6194));
    InMux I__1167 (
            .O(N__6199),
            .I(N__6191));
    Odrv4 I__1166 (
            .O(N__6194),
            .I(REG_CYCLEm));
    LocalMux I__1165 (
            .O(N__6191),
            .I(REG_CYCLEm));
    IoInMux I__1164 (
            .O(N__6186),
            .I(N__6183));
    LocalMux I__1163 (
            .O(N__6183),
            .I(N__6180));
    Span4Mux_s2_v I__1162 (
            .O(N__6180),
            .I(N__6177));
    Span4Mux_h I__1161 (
            .O(N__6177),
            .I(N__6174));
    Span4Mux_h I__1160 (
            .O(N__6174),
            .I(N__6171));
    Sp12to4 I__1159 (
            .O(N__6171),
            .I(N__6168));
    Span12Mux_s11_v I__1158 (
            .O(N__6168),
            .I(N__6165));
    Odrv12 I__1157 (
            .O(N__6165),
            .I(DRDENn_c));
    IoInMux I__1156 (
            .O(N__6162),
            .I(N__6159));
    LocalMux I__1155 (
            .O(N__6159),
            .I(N__6156));
    IoSpan4Mux I__1154 (
            .O(N__6156),
            .I(N__6153));
    IoSpan4Mux I__1153 (
            .O(N__6153),
            .I(N__6150));
    Span4Mux_s1_v I__1152 (
            .O(N__6150),
            .I(N__6147));
    Sp12to4 I__1151 (
            .O(N__6147),
            .I(N__6144));
    Span12Mux_s9_v I__1150 (
            .O(N__6144),
            .I(N__6141));
    Odrv12 I__1149 (
            .O(N__6141),
            .I(un1_LDSn_i_0));
    InMux I__1148 (
            .O(N__6138),
            .I(N__6129));
    InMux I__1147 (
            .O(N__6137),
            .I(N__6129));
    InMux I__1146 (
            .O(N__6136),
            .I(N__6129));
    LocalMux I__1145 (
            .O(N__6129),
            .I(N__6126));
    Span4Mux_v I__1144 (
            .O(N__6126),
            .I(N__6120));
    InMux I__1143 (
            .O(N__6125),
            .I(N__6115));
    InMux I__1142 (
            .O(N__6124),
            .I(N__6115));
    InMux I__1141 (
            .O(N__6123),
            .I(N__6112));
    Span4Mux_v I__1140 (
            .O(N__6120),
            .I(N__6107));
    LocalMux I__1139 (
            .O(N__6115),
            .I(N__6107));
    LocalMux I__1138 (
            .O(N__6112),
            .I(N__6104));
    Span4Mux_v I__1137 (
            .O(N__6107),
            .I(N__6101));
    Sp12to4 I__1136 (
            .O(N__6104),
            .I(N__6098));
    Sp12to4 I__1135 (
            .O(N__6101),
            .I(N__6095));
    Span12Mux_v I__1134 (
            .O(N__6098),
            .I(N__6092));
    Span12Mux_h I__1133 (
            .O(N__6095),
            .I(N__6089));
    Odrv12 I__1132 (
            .O(N__6092),
            .I(A_c_0));
    Odrv12 I__1131 (
            .O(N__6089),
            .I(A_c_0));
    InMux I__1130 (
            .O(N__6084),
            .I(N__6081));
    LocalMux I__1129 (
            .O(N__6081),
            .I(N__6077));
    CascadeMux I__1128 (
            .O(N__6080),
            .I(N__6074));
    Span4Mux_v I__1127 (
            .O(N__6077),
            .I(N__6070));
    InMux I__1126 (
            .O(N__6074),
            .I(N__6065));
    InMux I__1125 (
            .O(N__6073),
            .I(N__6065));
    Span4Mux_v I__1124 (
            .O(N__6070),
            .I(N__6060));
    LocalMux I__1123 (
            .O(N__6065),
            .I(N__6060));
    Span4Mux_v I__1122 (
            .O(N__6060),
            .I(N__6057));
    Span4Mux_v I__1121 (
            .O(N__6057),
            .I(N__6054));
    Sp12to4 I__1120 (
            .O(N__6054),
            .I(N__6051));
    Span12Mux_h I__1119 (
            .O(N__6051),
            .I(N__6048));
    Odrv12 I__1118 (
            .O(N__6048),
            .I(SIZ_c_0));
    InMux I__1117 (
            .O(N__6045),
            .I(N__6039));
    InMux I__1116 (
            .O(N__6044),
            .I(N__6039));
    LocalMux I__1115 (
            .O(N__6039),
            .I(N__6036));
    Span4Mux_v I__1114 (
            .O(N__6036),
            .I(N__6033));
    Span4Mux_v I__1113 (
            .O(N__6033),
            .I(N__6029));
    InMux I__1112 (
            .O(N__6032),
            .I(N__6026));
    Odrv4 I__1111 (
            .O(N__6029),
            .I(DS_ENm));
    LocalMux I__1110 (
            .O(N__6026),
            .I(DS_ENm));
    IoInMux I__1109 (
            .O(N__6021),
            .I(N__6018));
    LocalMux I__1108 (
            .O(N__6018),
            .I(N__6015));
    Span12Mux_s9_v I__1107 (
            .O(N__6015),
            .I(N__6012));
    Span12Mux_h I__1106 (
            .O(N__6012),
            .I(N__6009));
    Odrv12 I__1105 (
            .O(N__6009),
            .I(un1_UDSn_i_0));
    InMux I__1104 (
            .O(N__6006),
            .I(N__6003));
    LocalMux I__1103 (
            .O(N__6003),
            .I(N__6000));
    Odrv4 I__1102 (
            .O(N__6000),
            .I(\U712_CHIP_RAM.N_242 ));
    InMux I__1101 (
            .O(N__5997),
            .I(N__5994));
    LocalMux I__1100 (
            .O(N__5994),
            .I(N__5991));
    Span4Mux_v I__1099 (
            .O(N__5991),
            .I(N__5988));
    Odrv4 I__1098 (
            .O(N__5988),
            .I(\U712_CHIP_RAM.DBENn_7_0 ));
    InMux I__1097 (
            .O(N__5985),
            .I(N__5982));
    LocalMux I__1096 (
            .O(N__5982),
            .I(N__5979));
    Odrv4 I__1095 (
            .O(N__5979),
            .I(\U712_CHIP_RAM.N_253 ));
    CascadeMux I__1094 (
            .O(N__5976),
            .I(N__5973));
    InMux I__1093 (
            .O(N__5973),
            .I(N__5969));
    InMux I__1092 (
            .O(N__5972),
            .I(N__5966));
    LocalMux I__1091 (
            .O(N__5969),
            .I(REG_TACK));
    LocalMux I__1090 (
            .O(N__5966),
            .I(REG_TACK));
    InMux I__1089 (
            .O(N__5961),
            .I(N__5958));
    LocalMux I__1088 (
            .O(N__5958),
            .I(\U712_CHIP_RAM.REFRESH_SYNCZ0Z_1 ));
    InMux I__1087 (
            .O(N__5955),
            .I(N__5951));
    InMux I__1086 (
            .O(N__5954),
            .I(N__5948));
    LocalMux I__1085 (
            .O(N__5951),
            .I(N__5945));
    LocalMux I__1084 (
            .O(N__5948),
            .I(N__5942));
    Span4Mux_h I__1083 (
            .O(N__5945),
            .I(N__5937));
    Span4Mux_h I__1082 (
            .O(N__5942),
            .I(N__5934));
    InMux I__1081 (
            .O(N__5941),
            .I(N__5931));
    InMux I__1080 (
            .O(N__5940),
            .I(N__5928));
    Odrv4 I__1079 (
            .O(N__5937),
            .I(\U712_REG_SM.N_188 ));
    Odrv4 I__1078 (
            .O(N__5934),
            .I(\U712_REG_SM.N_188 ));
    LocalMux I__1077 (
            .O(N__5931),
            .I(\U712_REG_SM.N_188 ));
    LocalMux I__1076 (
            .O(N__5928),
            .I(\U712_REG_SM.N_188 ));
    CascadeMux I__1075 (
            .O(N__5919),
            .I(N__5914));
    InMux I__1074 (
            .O(N__5918),
            .I(N__5911));
    InMux I__1073 (
            .O(N__5917),
            .I(N__5908));
    InMux I__1072 (
            .O(N__5914),
            .I(N__5905));
    LocalMux I__1071 (
            .O(N__5911),
            .I(N__5902));
    LocalMux I__1070 (
            .O(N__5908),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1069 (
            .O(N__5905),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    Odrv4 I__1068 (
            .O(N__5902),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    InMux I__1067 (
            .O(N__5895),
            .I(N__5892));
    LocalMux I__1066 (
            .O(N__5892),
            .I(N__5889));
    Span4Mux_v I__1065 (
            .O(N__5889),
            .I(N__5886));
    Sp12to4 I__1064 (
            .O(N__5886),
            .I(N__5883));
    Span12Mux_h I__1063 (
            .O(N__5883),
            .I(N__5880));
    Odrv12 I__1062 (
            .O(N__5880),
            .I(RAS1n_c));
    InMux I__1061 (
            .O(N__5877),
            .I(N__5873));
    InMux I__1060 (
            .O(N__5876),
            .I(N__5870));
    LocalMux I__1059 (
            .O(N__5873),
            .I(\U712_CHIP_RAM.REFRESH_SYNCZ0Z_0 ));
    LocalMux I__1058 (
            .O(N__5870),
            .I(\U712_CHIP_RAM.REFRESH_SYNCZ0Z_0 ));
    InMux I__1057 (
            .O(N__5865),
            .I(N__5860));
    InMux I__1056 (
            .O(N__5864),
            .I(N__5855));
    InMux I__1055 (
            .O(N__5863),
            .I(N__5855));
    LocalMux I__1054 (
            .O(N__5860),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1053 (
            .O(N__5855),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    CascadeMux I__1052 (
            .O(N__5850),
            .I(N__5847));
    InMux I__1051 (
            .O(N__5847),
            .I(N__5843));
    InMux I__1050 (
            .O(N__5846),
            .I(N__5839));
    LocalMux I__1049 (
            .O(N__5843),
            .I(N__5836));
    InMux I__1048 (
            .O(N__5842),
            .I(N__5833));
    LocalMux I__1047 (
            .O(N__5839),
            .I(N__5830));
    Odrv4 I__1046 (
            .O(N__5836),
            .I(\U712_REG_SM.N_200 ));
    LocalMux I__1045 (
            .O(N__5833),
            .I(\U712_REG_SM.N_200 ));
    Odrv4 I__1044 (
            .O(N__5830),
            .I(\U712_REG_SM.N_200 ));
    CascadeMux I__1043 (
            .O(N__5823),
            .I(N__5818));
    InMux I__1042 (
            .O(N__5822),
            .I(N__5814));
    InMux I__1041 (
            .O(N__5821),
            .I(N__5811));
    InMux I__1040 (
            .O(N__5818),
            .I(N__5808));
    InMux I__1039 (
            .O(N__5817),
            .I(N__5805));
    LocalMux I__1038 (
            .O(N__5814),
            .I(N__5800));
    LocalMux I__1037 (
            .O(N__5811),
            .I(N__5800));
    LocalMux I__1036 (
            .O(N__5808),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    LocalMux I__1035 (
            .O(N__5805),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    Odrv4 I__1034 (
            .O(N__5800),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    InMux I__1033 (
            .O(N__5793),
            .I(N__5790));
    LocalMux I__1032 (
            .O(N__5790),
            .I(N__5787));
    Odrv4 I__1031 (
            .O(N__5787),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    InMux I__1030 (
            .O(N__5784),
            .I(N__5781));
    LocalMux I__1029 (
            .O(N__5781),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    InMux I__1028 (
            .O(N__5778),
            .I(N__5775));
    LocalMux I__1027 (
            .O(N__5775),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    IoInMux I__1026 (
            .O(N__5772),
            .I(N__5769));
    LocalMux I__1025 (
            .O(N__5769),
            .I(N__5766));
    IoSpan4Mux I__1024 (
            .O(N__5766),
            .I(N__5763));
    Sp12to4 I__1023 (
            .O(N__5763),
            .I(N__5760));
    Span12Mux_s9_v I__1022 (
            .O(N__5760),
            .I(N__5757));
    Odrv12 I__1021 (
            .O(N__5757),
            .I(CMA_c_1));
    InMux I__1020 (
            .O(N__5754),
            .I(N__5751));
    LocalMux I__1019 (
            .O(N__5751),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__1018 (
            .O(N__5748),
            .I(N__5745));
    LocalMux I__1017 (
            .O(N__5745),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    IoInMux I__1016 (
            .O(N__5742),
            .I(N__5739));
    LocalMux I__1015 (
            .O(N__5739),
            .I(N__5736));
    IoSpan4Mux I__1014 (
            .O(N__5736),
            .I(N__5733));
    IoSpan4Mux I__1013 (
            .O(N__5733),
            .I(N__5730));
    Sp12to4 I__1012 (
            .O(N__5730),
            .I(N__5727));
    Span12Mux_s9_h I__1011 (
            .O(N__5727),
            .I(N__5724));
    Odrv12 I__1010 (
            .O(N__5724),
            .I(CMA_c_5));
    InMux I__1009 (
            .O(N__5721),
            .I(N__5718));
    LocalMux I__1008 (
            .O(N__5718),
            .I(N__5715));
    Span12Mux_v I__1007 (
            .O(N__5715),
            .I(N__5712));
    Span12Mux_h I__1006 (
            .O(N__5712),
            .I(N__5709));
    Odrv12 I__1005 (
            .O(N__5709),
            .I(A_c_6));
    InMux I__1004 (
            .O(N__5706),
            .I(N__5703));
    LocalMux I__1003 (
            .O(N__5703),
            .I(N__5700));
    Span12Mux_h I__1002 (
            .O(N__5700),
            .I(N__5697));
    Odrv12 I__1001 (
            .O(N__5697),
            .I(A_c_13));
    CascadeMux I__1000 (
            .O(N__5694),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ));
    InMux I__999 (
            .O(N__5691),
            .I(N__5688));
    LocalMux I__998 (
            .O(N__5688),
            .I(N__5685));
    Span12Mux_v I__997 (
            .O(N__5685),
            .I(N__5682));
    Span12Mux_h I__996 (
            .O(N__5682),
            .I(N__5679));
    Odrv12 I__995 (
            .O(N__5679),
            .I(A_c_4));
    InMux I__994 (
            .O(N__5676),
            .I(N__5673));
    LocalMux I__993 (
            .O(N__5673),
            .I(N__5670));
    Span4Mux_v I__992 (
            .O(N__5670),
            .I(N__5667));
    Sp12to4 I__991 (
            .O(N__5667),
            .I(N__5664));
    Span12Mux_h I__990 (
            .O(N__5664),
            .I(N__5661));
    Odrv12 I__989 (
            .O(N__5661),
            .I(A_c_11));
    InMux I__988 (
            .O(N__5658),
            .I(N__5655));
    LocalMux I__987 (
            .O(N__5655),
            .I(N__5652));
    Span4Mux_v I__986 (
            .O(N__5652),
            .I(N__5649));
    Span4Mux_v I__985 (
            .O(N__5649),
            .I(N__5646));
    Sp12to4 I__984 (
            .O(N__5646),
            .I(N__5643));
    Span12Mux_h I__983 (
            .O(N__5643),
            .I(N__5640));
    Odrv12 I__982 (
            .O(N__5640),
            .I(A_c_7));
    CascadeMux I__981 (
            .O(N__5637),
            .I(\U712_CHIP_RAM.N_324_cascade_ ));
    InMux I__980 (
            .O(N__5634),
            .I(N__5631));
    LocalMux I__979 (
            .O(N__5631),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    InMux I__978 (
            .O(N__5628),
            .I(N__5620));
    CascadeMux I__977 (
            .O(N__5627),
            .I(N__5617));
    InMux I__976 (
            .O(N__5626),
            .I(N__5610));
    InMux I__975 (
            .O(N__5625),
            .I(N__5610));
    InMux I__974 (
            .O(N__5624),
            .I(N__5597));
    InMux I__973 (
            .O(N__5623),
            .I(N__5597));
    LocalMux I__972 (
            .O(N__5620),
            .I(N__5593));
    InMux I__971 (
            .O(N__5617),
            .I(N__5590));
    InMux I__970 (
            .O(N__5616),
            .I(N__5587));
    InMux I__969 (
            .O(N__5615),
            .I(N__5579));
    LocalMux I__968 (
            .O(N__5610),
            .I(N__5576));
    InMux I__967 (
            .O(N__5609),
            .I(N__5573));
    InMux I__966 (
            .O(N__5608),
            .I(N__5570));
    InMux I__965 (
            .O(N__5607),
            .I(N__5563));
    InMux I__964 (
            .O(N__5606),
            .I(N__5563));
    InMux I__963 (
            .O(N__5605),
            .I(N__5563));
    InMux I__962 (
            .O(N__5604),
            .I(N__5556));
    InMux I__961 (
            .O(N__5603),
            .I(N__5556));
    InMux I__960 (
            .O(N__5602),
            .I(N__5556));
    LocalMux I__959 (
            .O(N__5597),
            .I(N__5553));
    InMux I__958 (
            .O(N__5596),
            .I(N__5550));
    Span4Mux_h I__957 (
            .O(N__5593),
            .I(N__5543));
    LocalMux I__956 (
            .O(N__5590),
            .I(N__5543));
    LocalMux I__955 (
            .O(N__5587),
            .I(N__5543));
    InMux I__954 (
            .O(N__5586),
            .I(N__5538));
    InMux I__953 (
            .O(N__5585),
            .I(N__5538));
    InMux I__952 (
            .O(N__5584),
            .I(N__5531));
    InMux I__951 (
            .O(N__5583),
            .I(N__5531));
    InMux I__950 (
            .O(N__5582),
            .I(N__5531));
    LocalMux I__949 (
            .O(N__5579),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__948 (
            .O(N__5576),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__947 (
            .O(N__5573),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__946 (
            .O(N__5570),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__945 (
            .O(N__5563),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__944 (
            .O(N__5556),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__943 (
            .O(N__5553),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__942 (
            .O(N__5550),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__941 (
            .O(N__5543),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__940 (
            .O(N__5538),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__939 (
            .O(N__5531),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    CascadeMux I__938 (
            .O(N__5508),
            .I(N__5504));
    InMux I__937 (
            .O(N__5507),
            .I(N__5500));
    InMux I__936 (
            .O(N__5504),
            .I(N__5497));
    CascadeMux I__935 (
            .O(N__5503),
            .I(N__5487));
    LocalMux I__934 (
            .O(N__5500),
            .I(N__5482));
    LocalMux I__933 (
            .O(N__5497),
            .I(N__5474));
    InMux I__932 (
            .O(N__5496),
            .I(N__5469));
    InMux I__931 (
            .O(N__5495),
            .I(N__5469));
    InMux I__930 (
            .O(N__5494),
            .I(N__5466));
    InMux I__929 (
            .O(N__5493),
            .I(N__5459));
    InMux I__928 (
            .O(N__5492),
            .I(N__5459));
    InMux I__927 (
            .O(N__5491),
            .I(N__5459));
    InMux I__926 (
            .O(N__5490),
            .I(N__5456));
    InMux I__925 (
            .O(N__5487),
            .I(N__5449));
    InMux I__924 (
            .O(N__5486),
            .I(N__5449));
    InMux I__923 (
            .O(N__5485),
            .I(N__5449));
    Span4Mux_h I__922 (
            .O(N__5482),
            .I(N__5446));
    InMux I__921 (
            .O(N__5481),
            .I(N__5443));
    InMux I__920 (
            .O(N__5480),
            .I(N__5440));
    InMux I__919 (
            .O(N__5479),
            .I(N__5437));
    InMux I__918 (
            .O(N__5478),
            .I(N__5432));
    InMux I__917 (
            .O(N__5477),
            .I(N__5432));
    Span4Mux_v I__916 (
            .O(N__5474),
            .I(N__5423));
    LocalMux I__915 (
            .O(N__5469),
            .I(N__5423));
    LocalMux I__914 (
            .O(N__5466),
            .I(N__5423));
    LocalMux I__913 (
            .O(N__5459),
            .I(N__5423));
    LocalMux I__912 (
            .O(N__5456),
            .I(N__5418));
    LocalMux I__911 (
            .O(N__5449),
            .I(N__5418));
    Odrv4 I__910 (
            .O(N__5446),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__909 (
            .O(N__5443),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__908 (
            .O(N__5440),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__907 (
            .O(N__5437),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__906 (
            .O(N__5432),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__905 (
            .O(N__5423),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__904 (
            .O(N__5418),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__903 (
            .O(N__5403),
            .I(N__5400));
    LocalMux I__902 (
            .O(N__5400),
            .I(N__5394));
    InMux I__901 (
            .O(N__5399),
            .I(N__5391));
    CascadeMux I__900 (
            .O(N__5398),
            .I(N__5387));
    InMux I__899 (
            .O(N__5397),
            .I(N__5382));
    Span4Mux_h I__898 (
            .O(N__5394),
            .I(N__5379));
    LocalMux I__897 (
            .O(N__5391),
            .I(N__5376));
    InMux I__896 (
            .O(N__5390),
            .I(N__5373));
    InMux I__895 (
            .O(N__5387),
            .I(N__5368));
    InMux I__894 (
            .O(N__5386),
            .I(N__5368));
    InMux I__893 (
            .O(N__5385),
            .I(N__5365));
    LocalMux I__892 (
            .O(N__5382),
            .I(\U712_CHIP_RAM.N_301 ));
    Odrv4 I__891 (
            .O(N__5379),
            .I(\U712_CHIP_RAM.N_301 ));
    Odrv4 I__890 (
            .O(N__5376),
            .I(\U712_CHIP_RAM.N_301 ));
    LocalMux I__889 (
            .O(N__5373),
            .I(\U712_CHIP_RAM.N_301 ));
    LocalMux I__888 (
            .O(N__5368),
            .I(\U712_CHIP_RAM.N_301 ));
    LocalMux I__887 (
            .O(N__5365),
            .I(\U712_CHIP_RAM.N_301 ));
    IoInMux I__886 (
            .O(N__5352),
            .I(N__5349));
    LocalMux I__885 (
            .O(N__5349),
            .I(N__5346));
    IoSpan4Mux I__884 (
            .O(N__5346),
            .I(N__5343));
    Span4Mux_s1_h I__883 (
            .O(N__5343),
            .I(N__5340));
    Span4Mux_v I__882 (
            .O(N__5340),
            .I(N__5337));
    Sp12to4 I__881 (
            .O(N__5337),
            .I(N__5334));
    Span12Mux_s10_h I__880 (
            .O(N__5334),
            .I(N__5331));
    Odrv12 I__879 (
            .O(N__5331),
            .I(CLK_EN_c));
    CEMux I__878 (
            .O(N__5328),
            .I(N__5325));
    LocalMux I__877 (
            .O(N__5325),
            .I(N__5322));
    Odrv12 I__876 (
            .O(N__5322),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0 ));
    CascadeMux I__875 (
            .O(N__5319),
            .I(\U712_REG_SM.N_204_cascade_ ));
    CascadeMux I__874 (
            .O(N__5316),
            .I(N__5313));
    InMux I__873 (
            .O(N__5313),
            .I(N__5308));
    InMux I__872 (
            .O(N__5312),
            .I(N__5305));
    InMux I__871 (
            .O(N__5311),
            .I(N__5302));
    LocalMux I__870 (
            .O(N__5308),
            .I(\U712_REG_SM.N_215 ));
    LocalMux I__869 (
            .O(N__5305),
            .I(\U712_REG_SM.N_215 ));
    LocalMux I__868 (
            .O(N__5302),
            .I(\U712_REG_SM.N_215 ));
    CascadeMux I__867 (
            .O(N__5295),
            .I(N__5291));
    InMux I__866 (
            .O(N__5294),
            .I(N__5288));
    InMux I__865 (
            .O(N__5291),
            .I(N__5285));
    LocalMux I__864 (
            .O(N__5288),
            .I(\U712_REG_SM.N_204 ));
    LocalMux I__863 (
            .O(N__5285),
            .I(\U712_REG_SM.N_204 ));
    InMux I__862 (
            .O(N__5280),
            .I(N__5275));
    InMux I__861 (
            .O(N__5279),
            .I(N__5270));
    InMux I__860 (
            .O(N__5278),
            .I(N__5270));
    LocalMux I__859 (
            .O(N__5275),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__858 (
            .O(N__5270),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    InMux I__857 (
            .O(N__5265),
            .I(N__5262));
    LocalMux I__856 (
            .O(N__5262),
            .I(N__5258));
    InMux I__855 (
            .O(N__5261),
            .I(N__5255));
    Span4Mux_v I__854 (
            .O(N__5258),
            .I(N__5250));
    LocalMux I__853 (
            .O(N__5255),
            .I(N__5250));
    Span4Mux_v I__852 (
            .O(N__5250),
            .I(N__5247));
    Span4Mux_v I__851 (
            .O(N__5247),
            .I(N__5244));
    Sp12to4 I__850 (
            .O(N__5244),
            .I(N__5241));
    Span12Mux_h I__849 (
            .O(N__5241),
            .I(N__5238));
    Odrv12 I__848 (
            .O(N__5238),
            .I(TSn_c));
    CascadeMux I__847 (
            .O(N__5235),
            .I(N__5232));
    InMux I__846 (
            .O(N__5232),
            .I(N__5229));
    LocalMux I__845 (
            .O(N__5229),
            .I(N__5226));
    Span4Mux_v I__844 (
            .O(N__5226),
            .I(N__5223));
    Span4Mux_v I__843 (
            .O(N__5223),
            .I(N__5220));
    Sp12to4 I__842 (
            .O(N__5220),
            .I(N__5217));
    Span12Mux_h I__841 (
            .O(N__5217),
            .I(N__5214));
    Odrv12 I__840 (
            .O(N__5214),
            .I(REGSPACEn_c));
    InMux I__839 (
            .O(N__5211),
            .I(N__5205));
    InMux I__838 (
            .O(N__5210),
            .I(N__5205));
    LocalMux I__837 (
            .O(N__5205),
            .I(\U712_REG_SM.REG_CYCLE_GOZ0 ));
    InMux I__836 (
            .O(N__5202),
            .I(N__5198));
    InMux I__835 (
            .O(N__5201),
            .I(N__5195));
    LocalMux I__834 (
            .O(N__5198),
            .I(\U712_REG_SM.N_209 ));
    LocalMux I__833 (
            .O(N__5195),
            .I(\U712_REG_SM.N_209 ));
    InMux I__832 (
            .O(N__5190),
            .I(N__5180));
    InMux I__831 (
            .O(N__5189),
            .I(N__5180));
    InMux I__830 (
            .O(N__5188),
            .I(N__5180));
    InMux I__829 (
            .O(N__5187),
            .I(N__5177));
    LocalMux I__828 (
            .O(N__5180),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__827 (
            .O(N__5177),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__826 (
            .O(N__5172),
            .I(N__5165));
    InMux I__825 (
            .O(N__5171),
            .I(N__5165));
    InMux I__824 (
            .O(N__5170),
            .I(N__5162));
    LocalMux I__823 (
            .O(N__5165),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa ));
    LocalMux I__822 (
            .O(N__5162),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa ));
    InMux I__821 (
            .O(N__5157),
            .I(N__5152));
    InMux I__820 (
            .O(N__5156),
            .I(N__5147));
    InMux I__819 (
            .O(N__5155),
            .I(N__5147));
    LocalMux I__818 (
            .O(N__5152),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__817 (
            .O(N__5147),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    InMux I__816 (
            .O(N__5142),
            .I(N__5136));
    InMux I__815 (
            .O(N__5141),
            .I(N__5136));
    LocalMux I__814 (
            .O(N__5136),
            .I(N__5133));
    Odrv4 I__813 (
            .O(N__5133),
            .I(DBR_SYNCZ0Z_0));
    IoInMux I__812 (
            .O(N__5130),
            .I(N__5127));
    LocalMux I__811 (
            .O(N__5127),
            .I(N__5124));
    Span4Mux_s0_v I__810 (
            .O(N__5124),
            .I(N__5121));
    Sp12to4 I__809 (
            .O(N__5121),
            .I(N__5118));
    Span12Mux_h I__808 (
            .O(N__5118),
            .I(N__5115));
    Odrv12 I__807 (
            .O(N__5115),
            .I(CMA_c_10));
    InMux I__806 (
            .O(N__5112),
            .I(N__5106));
    InMux I__805 (
            .O(N__5111),
            .I(N__5106));
    LocalMux I__804 (
            .O(N__5106),
            .I(CPU_TACKm));
    CascadeMux I__803 (
            .O(N__5103),
            .I(N__5096));
    InMux I__802 (
            .O(N__5102),
            .I(N__5091));
    InMux I__801 (
            .O(N__5101),
            .I(N__5091));
    InMux I__800 (
            .O(N__5100),
            .I(N__5088));
    InMux I__799 (
            .O(N__5099),
            .I(N__5083));
    InMux I__798 (
            .O(N__5096),
            .I(N__5083));
    LocalMux I__797 (
            .O(N__5091),
            .I(N__5080));
    LocalMux I__796 (
            .O(N__5088),
            .I(N__5077));
    LocalMux I__795 (
            .O(N__5083),
            .I(N__5072));
    Span4Mux_v I__794 (
            .O(N__5080),
            .I(N__5072));
    Odrv4 I__793 (
            .O(N__5077),
            .I(\U712_CHIP_RAM.REFRESH_SYNC_RNI5J861Z0Z_1 ));
    Odrv4 I__792 (
            .O(N__5072),
            .I(\U712_CHIP_RAM.REFRESH_SYNC_RNI5J861Z0Z_1 ));
    CascadeMux I__791 (
            .O(N__5067),
            .I(N__5064));
    InMux I__790 (
            .O(N__5064),
            .I(N__5061));
    LocalMux I__789 (
            .O(N__5061),
            .I(N__5058));
    Span4Mux_v I__788 (
            .O(N__5058),
            .I(N__5055));
    Sp12to4 I__787 (
            .O(N__5055),
            .I(N__5052));
    Span12Mux_h I__786 (
            .O(N__5052),
            .I(N__5049));
    Span12Mux_v I__785 (
            .O(N__5049),
            .I(N__5046));
    Odrv12 I__784 (
            .O(N__5046),
            .I(RAMSPACEn_c));
    CascadeMux I__783 (
            .O(N__5043),
            .I(N__5039));
    InMux I__782 (
            .O(N__5042),
            .I(N__5036));
    InMux I__781 (
            .O(N__5039),
            .I(N__5033));
    LocalMux I__780 (
            .O(N__5036),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__779 (
            .O(N__5033),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__778 (
            .O(N__5028),
            .I(N__5022));
    InMux I__777 (
            .O(N__5027),
            .I(N__5022));
    LocalMux I__776 (
            .O(N__5022),
            .I(DBR_SYNCZ0Z_1));
    CascadeMux I__775 (
            .O(N__5019),
            .I(N__5016));
    InMux I__774 (
            .O(N__5016),
            .I(N__5010));
    InMux I__773 (
            .O(N__5015),
            .I(N__5010));
    LocalMux I__772 (
            .O(N__5010),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    InMux I__771 (
            .O(N__5007),
            .I(N__5004));
    LocalMux I__770 (
            .O(N__5004),
            .I(\U712_REG_SM.N_197 ));
    CascadeMux I__769 (
            .O(N__5001),
            .I(\U712_REG_SM.N_215_cascade_ ));
    IoInMux I__768 (
            .O(N__4998),
            .I(N__4995));
    LocalMux I__767 (
            .O(N__4995),
            .I(N__4991));
    IoInMux I__766 (
            .O(N__4994),
            .I(N__4988));
    Span4Mux_s2_v I__765 (
            .O(N__4991),
            .I(N__4985));
    LocalMux I__764 (
            .O(N__4988),
            .I(N__4982));
    Span4Mux_h I__763 (
            .O(N__4985),
            .I(N__4979));
    IoSpan4Mux I__762 (
            .O(N__4982),
            .I(N__4976));
    Span4Mux_v I__761 (
            .O(N__4979),
            .I(N__4973));
    IoSpan4Mux I__760 (
            .O(N__4976),
            .I(N__4970));
    Sp12to4 I__759 (
            .O(N__4973),
            .I(N__4967));
    Sp12to4 I__758 (
            .O(N__4970),
            .I(N__4964));
    Span12Mux_h I__757 (
            .O(N__4967),
            .I(N__4958));
    Span12Mux_s6_v I__756 (
            .O(N__4964),
            .I(N__4958));
    InMux I__755 (
            .O(N__4963),
            .I(N__4955));
    Odrv12 I__754 (
            .O(N__4958),
            .I(ASn_c));
    LocalMux I__753 (
            .O(N__4955),
            .I(ASn_c));
    InMux I__752 (
            .O(N__4950),
            .I(N__4943));
    InMux I__751 (
            .O(N__4949),
            .I(N__4943));
    InMux I__750 (
            .O(N__4948),
            .I(N__4938));
    LocalMux I__749 (
            .O(N__4943),
            .I(N__4935));
    InMux I__748 (
            .O(N__4942),
            .I(N__4932));
    InMux I__747 (
            .O(N__4941),
            .I(N__4929));
    LocalMux I__746 (
            .O(N__4938),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    Odrv4 I__745 (
            .O(N__4935),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__744 (
            .O(N__4932),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__743 (
            .O(N__4929),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    CascadeMux I__742 (
            .O(N__4920),
            .I(N__4917));
    InMux I__741 (
            .O(N__4917),
            .I(N__4914));
    LocalMux I__740 (
            .O(N__4914),
            .I(N__4907));
    InMux I__739 (
            .O(N__4913),
            .I(N__4904));
    InMux I__738 (
            .O(N__4912),
            .I(N__4900));
    InMux I__737 (
            .O(N__4911),
            .I(N__4895));
    InMux I__736 (
            .O(N__4910),
            .I(N__4895));
    Span4Mux_v I__735 (
            .O(N__4907),
            .I(N__4890));
    LocalMux I__734 (
            .O(N__4904),
            .I(N__4890));
    InMux I__733 (
            .O(N__4903),
            .I(N__4887));
    LocalMux I__732 (
            .O(N__4900),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__731 (
            .O(N__4895),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__730 (
            .O(N__4890),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__729 (
            .O(N__4887),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__728 (
            .O(N__4878),
            .I(N__4875));
    LocalMux I__727 (
            .O(N__4875),
            .I(\U712_REG_SM.N_185 ));
    InMux I__726 (
            .O(N__4872),
            .I(N__4865));
    CascadeMux I__725 (
            .O(N__4871),
            .I(N__4861));
    CascadeMux I__724 (
            .O(N__4870),
            .I(N__4857));
    InMux I__723 (
            .O(N__4869),
            .I(N__4846));
    InMux I__722 (
            .O(N__4868),
            .I(N__4846));
    LocalMux I__721 (
            .O(N__4865),
            .I(N__4843));
    InMux I__720 (
            .O(N__4864),
            .I(N__4840));
    InMux I__719 (
            .O(N__4861),
            .I(N__4837));
    InMux I__718 (
            .O(N__4860),
            .I(N__4834));
    InMux I__717 (
            .O(N__4857),
            .I(N__4831));
    InMux I__716 (
            .O(N__4856),
            .I(N__4826));
    InMux I__715 (
            .O(N__4855),
            .I(N__4826));
    InMux I__714 (
            .O(N__4854),
            .I(N__4821));
    InMux I__713 (
            .O(N__4853),
            .I(N__4821));
    InMux I__712 (
            .O(N__4852),
            .I(N__4816));
    InMux I__711 (
            .O(N__4851),
            .I(N__4816));
    LocalMux I__710 (
            .O(N__4846),
            .I(N__4813));
    Odrv4 I__709 (
            .O(N__4843),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__708 (
            .O(N__4840),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__707 (
            .O(N__4837),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__706 (
            .O(N__4834),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__705 (
            .O(N__4831),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__704 (
            .O(N__4826),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__703 (
            .O(N__4821),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__702 (
            .O(N__4816),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__701 (
            .O(N__4813),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__700 (
            .O(N__4794),
            .I(N__4791));
    LocalMux I__699 (
            .O(N__4791),
            .I(\U712_CHIP_RAM.N_198_i ));
    CascadeMux I__698 (
            .O(N__4788),
            .I(N__4784));
    CascadeMux I__697 (
            .O(N__4787),
            .I(N__4781));
    InMux I__696 (
            .O(N__4784),
            .I(N__4778));
    InMux I__695 (
            .O(N__4781),
            .I(N__4772));
    LocalMux I__694 (
            .O(N__4778),
            .I(N__4769));
    InMux I__693 (
            .O(N__4777),
            .I(N__4766));
    InMux I__692 (
            .O(N__4776),
            .I(N__4763));
    InMux I__691 (
            .O(N__4775),
            .I(N__4760));
    LocalMux I__690 (
            .O(N__4772),
            .I(\U712_CHIP_RAM.N_187 ));
    Odrv4 I__689 (
            .O(N__4769),
            .I(\U712_CHIP_RAM.N_187 ));
    LocalMux I__688 (
            .O(N__4766),
            .I(\U712_CHIP_RAM.N_187 ));
    LocalMux I__687 (
            .O(N__4763),
            .I(\U712_CHIP_RAM.N_187 ));
    LocalMux I__686 (
            .O(N__4760),
            .I(\U712_CHIP_RAM.N_187 ));
    InMux I__685 (
            .O(N__4749),
            .I(N__4745));
    InMux I__684 (
            .O(N__4748),
            .I(N__4742));
    LocalMux I__683 (
            .O(N__4745),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__682 (
            .O(N__4742),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__681 (
            .O(N__4737),
            .I(N__4733));
    InMux I__680 (
            .O(N__4736),
            .I(N__4730));
    LocalMux I__679 (
            .O(N__4733),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__678 (
            .O(N__4730),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__677 (
            .O(N__4725),
            .I(N__4721));
    InMux I__676 (
            .O(N__4724),
            .I(N__4718));
    InMux I__675 (
            .O(N__4721),
            .I(N__4715));
    LocalMux I__674 (
            .O(N__4718),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__673 (
            .O(N__4715),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__672 (
            .O(N__4710),
            .I(N__4706));
    InMux I__671 (
            .O(N__4709),
            .I(N__4703));
    LocalMux I__670 (
            .O(N__4706),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__669 (
            .O(N__4703),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    CascadeMux I__668 (
            .O(N__4698),
            .I(\U712_CHIP_RAM.N_355_cascade_ ));
    InMux I__667 (
            .O(N__4695),
            .I(N__4692));
    LocalMux I__666 (
            .O(N__4692),
            .I(N__4689));
    Span4Mux_v I__665 (
            .O(N__4689),
            .I(N__4685));
    InMux I__664 (
            .O(N__4688),
            .I(N__4682));
    Odrv4 I__663 (
            .O(N__4685),
            .I(\U712_CHIP_RAM.N_321 ));
    LocalMux I__662 (
            .O(N__4682),
            .I(\U712_CHIP_RAM.N_321 ));
    InMux I__661 (
            .O(N__4677),
            .I(N__4674));
    LocalMux I__660 (
            .O(N__4674),
            .I(\U712_CHIP_RAM.N_235 ));
    InMux I__659 (
            .O(N__4671),
            .I(N__4666));
    InMux I__658 (
            .O(N__4670),
            .I(N__4663));
    CascadeMux I__657 (
            .O(N__4669),
            .I(N__4655));
    LocalMux I__656 (
            .O(N__4666),
            .I(N__4651));
    LocalMux I__655 (
            .O(N__4663),
            .I(N__4648));
    CascadeMux I__654 (
            .O(N__4662),
            .I(N__4644));
    InMux I__653 (
            .O(N__4661),
            .I(N__4639));
    InMux I__652 (
            .O(N__4660),
            .I(N__4636));
    InMux I__651 (
            .O(N__4659),
            .I(N__4633));
    InMux I__650 (
            .O(N__4658),
            .I(N__4630));
    InMux I__649 (
            .O(N__4655),
            .I(N__4625));
    InMux I__648 (
            .O(N__4654),
            .I(N__4625));
    Span4Mux_v I__647 (
            .O(N__4651),
            .I(N__4622));
    Span4Mux_v I__646 (
            .O(N__4648),
            .I(N__4619));
    InMux I__645 (
            .O(N__4647),
            .I(N__4614));
    InMux I__644 (
            .O(N__4644),
            .I(N__4614));
    InMux I__643 (
            .O(N__4643),
            .I(N__4609));
    InMux I__642 (
            .O(N__4642),
            .I(N__4609));
    LocalMux I__641 (
            .O(N__4639),
            .I(N__4604));
    LocalMux I__640 (
            .O(N__4636),
            .I(N__4604));
    LocalMux I__639 (
            .O(N__4633),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__638 (
            .O(N__4630),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__637 (
            .O(N__4625),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__636 (
            .O(N__4622),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__635 (
            .O(N__4619),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__634 (
            .O(N__4614),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__633 (
            .O(N__4609),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__632 (
            .O(N__4604),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__631 (
            .O(N__4587),
            .I(N__4584));
    LocalMux I__630 (
            .O(N__4584),
            .I(N__4580));
    InMux I__629 (
            .O(N__4583),
            .I(N__4577));
    Span4Mux_h I__628 (
            .O(N__4580),
            .I(N__4574));
    LocalMux I__627 (
            .O(N__4577),
            .I(\U712_CHIP_RAM.N_217 ));
    Odrv4 I__626 (
            .O(N__4574),
            .I(\U712_CHIP_RAM.N_217 ));
    CascadeMux I__625 (
            .O(N__4569),
            .I(\U712_CHIP_RAM.CPU_TACK_8_iv_i_i_2_cascade_ ));
    InMux I__624 (
            .O(N__4566),
            .I(N__4563));
    LocalMux I__623 (
            .O(N__4563),
            .I(N__4560));
    Span4Mux_h I__622 (
            .O(N__4560),
            .I(N__4557));
    Odrv4 I__621 (
            .O(N__4557),
            .I(\U712_CHIP_RAM.N_219 ));
    CascadeMux I__620 (
            .O(N__4554),
            .I(\U712_CHIP_RAM.N_117_cascade_ ));
    InMux I__619 (
            .O(N__4551),
            .I(N__4548));
    LocalMux I__618 (
            .O(N__4548),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_i_0_1 ));
    InMux I__617 (
            .O(N__4545),
            .I(N__4538));
    InMux I__616 (
            .O(N__4544),
            .I(N__4538));
    InMux I__615 (
            .O(N__4543),
            .I(N__4535));
    LocalMux I__614 (
            .O(N__4538),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ));
    LocalMux I__613 (
            .O(N__4535),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ));
    InMux I__612 (
            .O(N__4530),
            .I(N__4524));
    InMux I__611 (
            .O(N__4529),
            .I(N__4524));
    LocalMux I__610 (
            .O(N__4524),
            .I(\U712_CHIP_RAM.N_42_1 ));
    InMux I__609 (
            .O(N__4521),
            .I(N__4518));
    LocalMux I__608 (
            .O(N__4518),
            .I(\U712_CHIP_RAM.N_236 ));
    InMux I__607 (
            .O(N__4515),
            .I(N__4512));
    LocalMux I__606 (
            .O(N__4512),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    InMux I__605 (
            .O(N__4509),
            .I(N__4506));
    LocalMux I__604 (
            .O(N__4506),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_0 ));
    InMux I__603 (
            .O(N__4503),
            .I(N__4500));
    LocalMux I__602 (
            .O(N__4500),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_1 ));
    CascadeMux I__601 (
            .O(N__4497),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_cascade_ ));
    CascadeMux I__600 (
            .O(N__4494),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_cascade_ ));
    CascadeMux I__599 (
            .O(N__4491),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ));
    InMux I__598 (
            .O(N__4488),
            .I(N__4482));
    InMux I__597 (
            .O(N__4487),
            .I(N__4482));
    LocalMux I__596 (
            .O(N__4482),
            .I(N__4479));
    Span4Mux_v I__595 (
            .O(N__4479),
            .I(N__4476));
    Span4Mux_h I__594 (
            .O(N__4476),
            .I(N__4473));
    Sp12to4 I__593 (
            .O(N__4473),
            .I(N__4470));
    Odrv12 I__592 (
            .O(N__4470),
            .I(A_c_14));
    InMux I__591 (
            .O(N__4467),
            .I(N__4464));
    LocalMux I__590 (
            .O(N__4464),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ));
    InMux I__589 (
            .O(N__4461),
            .I(N__4458));
    LocalMux I__588 (
            .O(N__4458),
            .I(N__4455));
    Span4Mux_v I__587 (
            .O(N__4455),
            .I(N__4452));
    Span4Mux_v I__586 (
            .O(N__4452),
            .I(N__4449));
    Sp12to4 I__585 (
            .O(N__4449),
            .I(N__4446));
    Odrv12 I__584 (
            .O(N__4446),
            .I(A_c_15));
    InMux I__583 (
            .O(N__4443),
            .I(N__4440));
    LocalMux I__582 (
            .O(N__4440),
            .I(N__4437));
    Sp12to4 I__581 (
            .O(N__4437),
            .I(N__4434));
    Span12Mux_v I__580 (
            .O(N__4434),
            .I(N__4431));
    Span12Mux_h I__579 (
            .O(N__4431),
            .I(N__4428));
    Odrv12 I__578 (
            .O(N__4428),
            .I(A_c_8));
    CascadeMux I__577 (
            .O(N__4425),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_0_cascade_ ));
    CascadeMux I__576 (
            .O(N__4422),
            .I(\U712_REG_SM.N_185_cascade_ ));
    InMux I__575 (
            .O(N__4419),
            .I(N__4416));
    LocalMux I__574 (
            .O(N__4416),
            .I(N__4412));
    IoInMux I__573 (
            .O(N__4415),
            .I(N__4409));
    Span4Mux_v I__572 (
            .O(N__4412),
            .I(N__4406));
    LocalMux I__571 (
            .O(N__4409),
            .I(N__4403));
    Sp12to4 I__570 (
            .O(N__4406),
            .I(N__4400));
    Span4Mux_s3_h I__569 (
            .O(N__4403),
            .I(N__4397));
    Span12Mux_h I__568 (
            .O(N__4400),
            .I(N__4392));
    Sp12to4 I__567 (
            .O(N__4397),
            .I(N__4392));
    Span12Mux_v I__566 (
            .O(N__4392),
            .I(N__4389));
    Odrv12 I__565 (
            .O(N__4389),
            .I(C1_c));
    CascadeMux I__564 (
            .O(N__4386),
            .I(\U712_REG_SM.N_197_cascade_ ));
    InMux I__563 (
            .O(N__4383),
            .I(N__4376));
    InMux I__562 (
            .O(N__4382),
            .I(N__4376));
    InMux I__561 (
            .O(N__4381),
            .I(N__4373));
    LocalMux I__560 (
            .O(N__4376),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    LocalMux I__559 (
            .O(N__4373),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    CascadeMux I__558 (
            .O(N__4368),
            .I(N__4365));
    InMux I__557 (
            .O(N__4365),
            .I(N__4361));
    InMux I__556 (
            .O(N__4364),
            .I(N__4356));
    LocalMux I__555 (
            .O(N__4361),
            .I(N__4353));
    InMux I__554 (
            .O(N__4360),
            .I(N__4350));
    InMux I__553 (
            .O(N__4359),
            .I(N__4347));
    LocalMux I__552 (
            .O(N__4356),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    Odrv4 I__551 (
            .O(N__4353),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__550 (
            .O(N__4350),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__549 (
            .O(N__4347),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__548 (
            .O(N__4338),
            .I(N__4330));
    InMux I__547 (
            .O(N__4337),
            .I(N__4330));
    InMux I__546 (
            .O(N__4336),
            .I(N__4327));
    InMux I__545 (
            .O(N__4335),
            .I(N__4324));
    LocalMux I__544 (
            .O(N__4330),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__543 (
            .O(N__4327),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__542 (
            .O(N__4324),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    CascadeMux I__541 (
            .O(N__4317),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa_0_a2_0_a3_1_cascade_ ));
    CascadeMux I__540 (
            .O(N__4314),
            .I(N__4308));
    CascadeMux I__539 (
            .O(N__4313),
            .I(N__4305));
    InMux I__538 (
            .O(N__4312),
            .I(N__4298));
    InMux I__537 (
            .O(N__4311),
            .I(N__4298));
    InMux I__536 (
            .O(N__4308),
            .I(N__4298));
    InMux I__535 (
            .O(N__4305),
            .I(N__4295));
    LocalMux I__534 (
            .O(N__4298),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__533 (
            .O(N__4295),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    CascadeMux I__532 (
            .O(N__4290),
            .I(\U712_REG_SM.DS_EN_0_sqmuxa_cascade_ ));
    InMux I__531 (
            .O(N__4287),
            .I(N__4281));
    InMux I__530 (
            .O(N__4286),
            .I(N__4281));
    LocalMux I__529 (
            .O(N__4281),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    InMux I__528 (
            .O(N__4278),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__527 (
            .O(N__4275),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__526 (
            .O(N__4272),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__525 (
            .O(N__4269),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    CascadeMux I__524 (
            .O(N__4266),
            .I(N__4263));
    InMux I__523 (
            .O(N__4263),
            .I(N__4260));
    LocalMux I__522 (
            .O(N__4260),
            .I(N__4250));
    InMux I__521 (
            .O(N__4259),
            .I(N__4243));
    InMux I__520 (
            .O(N__4258),
            .I(N__4243));
    InMux I__519 (
            .O(N__4257),
            .I(N__4243));
    InMux I__518 (
            .O(N__4256),
            .I(N__4236));
    InMux I__517 (
            .O(N__4255),
            .I(N__4236));
    InMux I__516 (
            .O(N__4254),
            .I(N__4236));
    InMux I__515 (
            .O(N__4253),
            .I(N__4233));
    Odrv4 I__514 (
            .O(N__4250),
            .I(\U712_CHIP_RAM.N_46 ));
    LocalMux I__513 (
            .O(N__4243),
            .I(\U712_CHIP_RAM.N_46 ));
    LocalMux I__512 (
            .O(N__4236),
            .I(\U712_CHIP_RAM.N_46 ));
    LocalMux I__511 (
            .O(N__4233),
            .I(\U712_CHIP_RAM.N_46 ));
    InMux I__510 (
            .O(N__4224),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    CEMux I__509 (
            .O(N__4221),
            .I(N__4217));
    CEMux I__508 (
            .O(N__4220),
            .I(N__4214));
    LocalMux I__507 (
            .O(N__4217),
            .I(\U712_CHIP_RAM.N_256_i ));
    LocalMux I__506 (
            .O(N__4214),
            .I(\U712_CHIP_RAM.N_256_i ));
    CascadeMux I__505 (
            .O(N__4209),
            .I(\U712_CYCLE_TERM.N_207_i_0_en_cascade_ ));
    InMux I__504 (
            .O(N__4206),
            .I(N__4203));
    LocalMux I__503 (
            .O(N__4203),
            .I(N__4200));
    Span12Mux_v I__502 (
            .O(N__4200),
            .I(N__4197));
    Odrv12 I__501 (
            .O(N__4197),
            .I(TACK_EN_i_ess));
    CEMux I__500 (
            .O(N__4194),
            .I(N__4191));
    LocalMux I__499 (
            .O(N__4191),
            .I(N__4188));
    Odrv4 I__498 (
            .O(N__4188),
            .I(\U712_CYCLE_TERM.N_207_i_0_en_0 ));
    CascadeMux I__497 (
            .O(N__4185),
            .I(\U712_CHIP_RAM.N_242_cascade_ ));
    InMux I__496 (
            .O(N__4182),
            .I(N__4179));
    LocalMux I__495 (
            .O(N__4179),
            .I(N__4176));
    Odrv4 I__494 (
            .O(N__4176),
            .I(\U712_CHIP_RAM.N_319 ));
    InMux I__493 (
            .O(N__4173),
            .I(N__4168));
    InMux I__492 (
            .O(N__4172),
            .I(N__4163));
    InMux I__491 (
            .O(N__4171),
            .I(N__4163));
    LocalMux I__490 (
            .O(N__4168),
            .I(N__4160));
    LocalMux I__489 (
            .O(N__4163),
            .I(\U712_CHIP_RAM.N_307 ));
    Odrv4 I__488 (
            .O(N__4160),
            .I(\U712_CHIP_RAM.N_307 ));
    InMux I__487 (
            .O(N__4155),
            .I(N__4151));
    InMux I__486 (
            .O(N__4154),
            .I(N__4148));
    LocalMux I__485 (
            .O(N__4151),
            .I(N__4143));
    LocalMux I__484 (
            .O(N__4148),
            .I(N__4140));
    InMux I__483 (
            .O(N__4147),
            .I(N__4137));
    InMux I__482 (
            .O(N__4146),
            .I(N__4134));
    Span4Mux_v I__481 (
            .O(N__4143),
            .I(N__4129));
    Span4Mux_v I__480 (
            .O(N__4140),
            .I(N__4129));
    LocalMux I__479 (
            .O(N__4137),
            .I(\U712_CHIP_RAM.N_177 ));
    LocalMux I__478 (
            .O(N__4134),
            .I(\U712_CHIP_RAM.N_177 ));
    Odrv4 I__477 (
            .O(N__4129),
            .I(\U712_CHIP_RAM.N_177 ));
    CascadeMux I__476 (
            .O(N__4122),
            .I(\U712_CHIP_RAM.N_319_cascade_ ));
    InMux I__475 (
            .O(N__4119),
            .I(N__4115));
    InMux I__474 (
            .O(N__4118),
            .I(N__4112));
    LocalMux I__473 (
            .O(N__4115),
            .I(\U712_CHIP_RAM.N_322 ));
    LocalMux I__472 (
            .O(N__4112),
            .I(\U712_CHIP_RAM.N_322 ));
    InMux I__471 (
            .O(N__4107),
            .I(N__4102));
    InMux I__470 (
            .O(N__4106),
            .I(N__4095));
    InMux I__469 (
            .O(N__4105),
            .I(N__4095));
    LocalMux I__468 (
            .O(N__4102),
            .I(N__4092));
    InMux I__467 (
            .O(N__4101),
            .I(N__4089));
    InMux I__466 (
            .O(N__4100),
            .I(N__4086));
    LocalMux I__465 (
            .O(N__4095),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__464 (
            .O(N__4092),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__463 (
            .O(N__4089),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__462 (
            .O(N__4086),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    InMux I__461 (
            .O(N__4077),
            .I(N__4072));
    InMux I__460 (
            .O(N__4076),
            .I(N__4067));
    InMux I__459 (
            .O(N__4075),
            .I(N__4067));
    LocalMux I__458 (
            .O(N__4072),
            .I(\U712_CHIP_RAM.N_311 ));
    LocalMux I__457 (
            .O(N__4067),
            .I(\U712_CHIP_RAM.N_311 ));
    InMux I__456 (
            .O(N__4062),
            .I(N__4059));
    LocalMux I__455 (
            .O(N__4059),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_i_i_a3_0 ));
    InMux I__454 (
            .O(N__4056),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__453 (
            .O(N__4053),
            .I(N__4050));
    LocalMux I__452 (
            .O(N__4050),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__451 (
            .O(N__4047),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    CascadeMux I__450 (
            .O(N__4044),
            .I(\U712_CHIP_RAM.N_187_cascade_ ));
    CascadeMux I__449 (
            .O(N__4041),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_1_cascade_ ));
    CascadeMux I__448 (
            .O(N__4038),
            .I(\U712_CHIP_RAM.N_264_cascade_ ));
    InMux I__447 (
            .O(N__4035),
            .I(N__4032));
    LocalMux I__446 (
            .O(N__4032),
            .I(\U712_CHIP_RAM.N_262 ));
    CascadeMux I__445 (
            .O(N__4029),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_ ));
    CEMux I__444 (
            .O(N__4026),
            .I(N__4023));
    LocalMux I__443 (
            .O(N__4023),
            .I(N__4020));
    Span4Mux_h I__442 (
            .O(N__4020),
            .I(N__4017));
    Odrv4 I__441 (
            .O(N__4017),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0 ));
    InMux I__440 (
            .O(N__4014),
            .I(N__4011));
    LocalMux I__439 (
            .O(N__4011),
            .I(N__4008));
    Odrv4 I__438 (
            .O(N__4008),
            .I(\U712_CHIP_RAM.N_220 ));
    InMux I__437 (
            .O(N__4005),
            .I(N__4002));
    LocalMux I__436 (
            .O(N__4002),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0_1 ));
    CascadeMux I__435 (
            .O(N__3999),
            .I(N__3996));
    InMux I__434 (
            .O(N__3996),
            .I(N__3993));
    LocalMux I__433 (
            .O(N__3993),
            .I(N__3990));
    Odrv4 I__432 (
            .O(N__3990),
            .I(\U712_CHIP_RAM.N_323 ));
    InMux I__431 (
            .O(N__3987),
            .I(N__3984));
    LocalMux I__430 (
            .O(N__3984),
            .I(\U712_CHIP_RAM.N_176 ));
    InMux I__429 (
            .O(N__3981),
            .I(N__3978));
    LocalMux I__428 (
            .O(N__3978),
            .I(N__3975));
    Span4Mux_v I__427 (
            .O(N__3975),
            .I(N__3972));
    Span4Mux_h I__426 (
            .O(N__3972),
            .I(N__3969));
    Span4Mux_h I__425 (
            .O(N__3969),
            .I(N__3966));
    Odrv4 I__424 (
            .O(N__3966),
            .I(A_c_10));
    InMux I__423 (
            .O(N__3963),
            .I(N__3960));
    LocalMux I__422 (
            .O(N__3960),
            .I(N__3957));
    Span4Mux_v I__421 (
            .O(N__3957),
            .I(N__3954));
    Sp12to4 I__420 (
            .O(N__3954),
            .I(N__3951));
    Span12Mux_h I__419 (
            .O(N__3951),
            .I(N__3948));
    Span12Mux_v I__418 (
            .O(N__3948),
            .I(N__3945));
    Odrv12 I__417 (
            .O(N__3945),
            .I(A_c_3));
    InMux I__416 (
            .O(N__3942),
            .I(N__3939));
    LocalMux I__415 (
            .O(N__3939),
            .I(N__3936));
    Span12Mux_v I__414 (
            .O(N__3936),
            .I(N__3933));
    Odrv12 I__413 (
            .O(N__3933),
            .I(A_c_9));
    InMux I__412 (
            .O(N__3930),
            .I(N__3927));
    LocalMux I__411 (
            .O(N__3927),
            .I(N__3924));
    Span12Mux_v I__410 (
            .O(N__3924),
            .I(N__3921));
    Span12Mux_v I__409 (
            .O(N__3921),
            .I(N__3918));
    Odrv12 I__408 (
            .O(N__3918),
            .I(A_c_2));
    InMux I__407 (
            .O(N__3915),
            .I(N__3912));
    LocalMux I__406 (
            .O(N__3912),
            .I(N__3909));
    Odrv4 I__405 (
            .O(N__3909),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_1 ));
    CascadeMux I__404 (
            .O(N__3906),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_0_cascade_ ));
    InMux I__403 (
            .O(N__3903),
            .I(N__3900));
    LocalMux I__402 (
            .O(N__3900),
            .I(\U712_CHIP_RAM.N_193 ));
    CascadeMux I__401 (
            .O(N__3897),
            .I(\U712_CHIP_RAM.N_177_cascade_ ));
    InMux I__400 (
            .O(N__3894),
            .I(N__3891));
    LocalMux I__399 (
            .O(N__3891),
            .I(\U712_CHIP_RAM.N_223 ));
    InMux I__398 (
            .O(N__3888),
            .I(N__3885));
    LocalMux I__397 (
            .O(N__3885),
            .I(\U712_CHIP_RAM.N_300 ));
    CascadeMux I__396 (
            .O(N__3882),
            .I(\U712_CHIP_RAM.N_223_cascade_ ));
    InMux I__395 (
            .O(N__3879),
            .I(N__3876));
    LocalMux I__394 (
            .O(N__3876),
            .I(N__3872));
    IoInMux I__393 (
            .O(N__3875),
            .I(N__3869));
    Span4Mux_v I__392 (
            .O(N__3872),
            .I(N__3866));
    LocalMux I__391 (
            .O(N__3869),
            .I(N__3863));
    Sp12to4 I__390 (
            .O(N__3866),
            .I(N__3860));
    IoSpan4Mux I__389 (
            .O(N__3863),
            .I(N__3857));
    Span12Mux_h I__388 (
            .O(N__3860),
            .I(N__3854));
    IoSpan4Mux I__387 (
            .O(N__3857),
            .I(N__3851));
    Span12Mux_v I__386 (
            .O(N__3854),
            .I(N__3848));
    IoSpan4Mux I__385 (
            .O(N__3851),
            .I(N__3845));
    Odrv12 I__384 (
            .O(N__3848),
            .I(C3_c));
    Odrv4 I__383 (
            .O(N__3845),
            .I(C3_c));
    InMux I__382 (
            .O(N__3840),
            .I(N__3837));
    LocalMux I__381 (
            .O(N__3837),
            .I(N__3834));
    Odrv4 I__380 (
            .O(N__3834),
            .I(\U712_CHIP_RAM.N_213 ));
    IoInMux I__379 (
            .O(N__3831),
            .I(N__3828));
    LocalMux I__378 (
            .O(N__3828),
            .I(N__3825));
    Span12Mux_s3_v I__377 (
            .O(N__3825),
            .I(N__3822));
    Odrv12 I__376 (
            .O(N__3822),
            .I(VBENn_c));
    InMux I__375 (
            .O(N__3819),
            .I(N__3816));
    LocalMux I__374 (
            .O(N__3816),
            .I(N__3813));
    Span4Mux_v I__373 (
            .O(N__3813),
            .I(N__3810));
    Sp12to4 I__372 (
            .O(N__3810),
            .I(N__3807));
    Span12Mux_h I__371 (
            .O(N__3807),
            .I(N__3804));
    Odrv12 I__370 (
            .O(N__3804),
            .I(A_c_12));
    InMux I__369 (
            .O(N__3801),
            .I(N__3798));
    LocalMux I__368 (
            .O(N__3798),
            .I(N__3795));
    Span12Mux_v I__367 (
            .O(N__3795),
            .I(N__3792));
    Odrv12 I__366 (
            .O(N__3792),
            .I(A_c_5));
    CascadeMux I__365 (
            .O(N__3789),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ));
    InMux I__364 (
            .O(N__3786),
            .I(N__3783));
    LocalMux I__363 (
            .O(N__3783),
            .I(N__3780));
    Span4Mux_h I__362 (
            .O(N__3780),
            .I(N__3777));
    Sp12to4 I__361 (
            .O(N__3777),
            .I(N__3774));
    Span12Mux_v I__360 (
            .O(N__3774),
            .I(N__3771));
    Odrv12 I__359 (
            .O(N__3771),
            .I(A_c_18));
    InMux I__358 (
            .O(N__3768),
            .I(N__3765));
    LocalMux I__357 (
            .O(N__3765),
            .I(N__3762));
    Span4Mux_v I__356 (
            .O(N__3762),
            .I(N__3759));
    Span4Mux_v I__355 (
            .O(N__3759),
            .I(N__3756));
    Span4Mux_h I__354 (
            .O(N__3756),
            .I(N__3753));
    Sp12to4 I__353 (
            .O(N__3753),
            .I(N__3750));
    Odrv12 I__352 (
            .O(N__3750),
            .I(A_c_16));
    CascadeMux I__351 (
            .O(N__3747),
            .I(\U712_CHIP_RAM.N_253_cascade_ ));
    CascadeMux I__350 (
            .O(N__3744),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_cascade_ ));
    CEMux I__349 (
            .O(N__3741),
            .I(N__3738));
    LocalMux I__348 (
            .O(N__3738),
            .I(N__3735));
    Sp12to4 I__347 (
            .O(N__3735),
            .I(N__3732));
    Odrv12 I__346 (
            .O(N__3732),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0 ));
    CascadeMux I__345 (
            .O(N__3729),
            .I(\U712_CHIP_RAM.N_298_cascade_ ));
    CascadeMux I__344 (
            .O(N__3726),
            .I(\U712_CHIP_RAM.N_323_cascade_ ));
    InMux I__343 (
            .O(N__3723),
            .I(N__3716));
    InMux I__342 (
            .O(N__3722),
            .I(N__3716));
    InMux I__341 (
            .O(N__3721),
            .I(N__3713));
    LocalMux I__340 (
            .O(N__3716),
            .I(\U712_CHIP_RAM.N_304 ));
    LocalMux I__339 (
            .O(N__3713),
            .I(\U712_CHIP_RAM.N_304 ));
    InMux I__338 (
            .O(N__3708),
            .I(N__3705));
    LocalMux I__337 (
            .O(N__3705),
            .I(\U712_CHIP_RAM.N_216 ));
    CascadeMux I__336 (
            .O(N__3702),
            .I(\U712_CHIP_RAM.N_216_cascade_ ));
    CascadeMux I__335 (
            .O(N__3699),
            .I(\U712_CHIP_RAM.N_193_cascade_ ));
    CascadeMux I__334 (
            .O(N__3696),
            .I(\U712_CHIP_RAM.N_176_cascade_ ));
    IoInMux I__333 (
            .O(N__3693),
            .I(N__3690));
    LocalMux I__332 (
            .O(N__3690),
            .I(N__3687));
    IoSpan4Mux I__331 (
            .O(N__3687),
            .I(N__3684));
    Span4Mux_s1_h I__330 (
            .O(N__3684),
            .I(N__3681));
    Odrv4 I__329 (
            .O(N__3681),
            .I(CLK40_PLL_i_i));
    IoInMux I__328 (
            .O(N__3678),
            .I(N__3675));
    LocalMux I__327 (
            .O(N__3675),
            .I(N__3672));
    Span4Mux_s3_h I__326 (
            .O(N__3672),
            .I(N__3669));
    Span4Mux_v I__325 (
            .O(N__3669),
            .I(N__3666));
    Odrv4 I__324 (
            .O(N__3666),
            .I(N_897_i));
    IoInMux I__323 (
            .O(N__3663),
            .I(N__3660));
    LocalMux I__322 (
            .O(N__3660),
            .I(N__3657));
    Span4Mux_s2_v I__321 (
            .O(N__3657),
            .I(N__3654));
    Span4Mux_v I__320 (
            .O(N__3654),
            .I(N__3651));
    Span4Mux_h I__319 (
            .O(N__3651),
            .I(N__3648));
    Odrv4 I__318 (
            .O(N__3648),
            .I(CLK80_PLL_i_i));
    IoInMux I__317 (
            .O(N__3645),
            .I(N__3642));
    LocalMux I__316 (
            .O(N__3642),
            .I(N__3639));
    IoSpan4Mux I__315 (
            .O(N__3639),
            .I(N__3636));
    Span4Mux_s2_v I__314 (
            .O(N__3636),
            .I(N__3633));
    Sp12to4 I__313 (
            .O(N__3633),
            .I(N__3630));
    Span12Mux_v I__312 (
            .O(N__3630),
            .I(N__3627));
    Odrv12 I__311 (
            .O(N__3627),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__8866));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__8867));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__8869));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .I(N__8870));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__8868));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_8_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7698),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__4415),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__3875),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLK40_OUT_obuf_RNO_LC_1_9_5.C_ON=1'b0;
    defparam CLK40_OUT_obuf_RNO_LC_1_9_5.SEQ_MODE=4'b0000;
    defparam CLK40_OUT_obuf_RNO_LC_1_9_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLK40_OUT_obuf_RNO_LC_1_9_5 (
            .in0(N__6978),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_obuft_RNO_LC_2_17_0.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_2_17_0.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_2_17_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_obuft_RNO_LC_2_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4206),
            .lcout(N_897_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_7_1_5.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_7_1_5.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_7_1_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_7_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8127),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_5_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_5_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_5_5  (
            .in0(N__4182),
            .in1(N__6614),
            .in2(_gnd_net_),
            .in3(N__4695),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8106),
            .ce(),
            .sr(N__9391));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILL8G1_LC_7_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILL8G1_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILL8G1_LC_7_6_0 .LUT_INIT=16'b1101111100010011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNILL8G1_LC_7_6_0  (
            .in0(N__4107),
            .in1(N__4661),
            .in2(N__4871),
            .in3(N__5603),
            .lcout(\U712_CHIP_RAM.N_217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_7_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_7_6_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__6592),
            .in2(_gnd_net_),
            .in3(N__5485),
            .lcout(\U712_CHIP_RAM.N_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1_1_LC_7_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1_1_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1_1_LC_7_6_4 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1_1_LC_7_6_4  (
            .in0(N__5486),
            .in1(N__7784),
            .in2(_gnd_net_),
            .in3(N__5602),
            .lcout(\U712_CHIP_RAM.N_193 ),
            .ltout(\U712_CHIP_RAM.N_193_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_7_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_7_6_5 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_7_6_5  (
            .in0(N__6555),
            .in1(N__4583),
            .in2(N__3699),
            .in3(N__5615),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_2_1_LC_7_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_2_1_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_2_1_LC_7_6_6 .LUT_INIT=16'b0011001100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_2_1_LC_7_6_6  (
            .in0(N__6593),
            .in1(N__5604),
            .in2(N__5503),
            .in3(N__4147),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_6_7 .LUT_INIT=16'b0010000011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_6_7  (
            .in0(N__6486),
            .in1(N__6439),
            .in2(N__7788),
            .in3(N__6594),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_i_i_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_7_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_7_7_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_7_7_0  (
            .in0(N__5102),
            .in1(N__4077),
            .in2(_gnd_net_),
            .in3(N__6385),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8114),
            .ce(N__3741),
            .sr(N__9376));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIMTA11_LC_7_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIMTA11_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIMTA11_LC_7_7_1 .LUT_INIT=16'b1010101001000100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIMTA11_LC_7_7_1  (
            .in0(N__5478),
            .in1(N__4100),
            .in2(_gnd_net_),
            .in3(N__4856),
            .lcout(\U712_CHIP_RAM.N_176 ),
            .ltout(\U712_CHIP_RAM.N_176_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_7_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_7_7_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_7_7_2  (
            .in0(N__4647),
            .in1(N__4775),
            .in2(N__3696),
            .in3(N__5586),
            .lcout(\U712_CHIP_RAM.N_253 ),
            .ltout(\U712_CHIP_RAM.N_253_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_7_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_7_7_3 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_7_7_3  (
            .in0(N__6384),
            .in1(N__3721),
            .in2(N__3747),
            .in3(N__5101),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_7_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_7_7_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_7_7_4  (
            .in0(N__9416),
            .in1(_gnd_net_),
            .in2(N__3744),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_7_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_7_7_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_7_7_6  (
            .in0(N__4855),
            .in1(N__5477),
            .in2(N__4662),
            .in3(N__5585),
            .lcout(\U712_CHIP_RAM.N_298 ),
            .ltout(\U712_CHIP_RAM.N_298_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_7_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_7_7_7 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_7_7_7  (
            .in0(N__6636),
            .in1(_gnd_net_),
            .in2(N__3729),
            .in3(N__6549),
            .lcout(\U712_CHIP_RAM.N_304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIV2P76_LC_7_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIV2P76_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIV2P76_LC_7_8_0 .LUT_INIT=16'b1010000010100010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIV2P76_LC_7_8_0  (
            .in0(N__3722),
            .in1(N__6484),
            .in2(N__6447),
            .in3(N__5099),
            .lcout(\U712_CHIP_RAM.N_323 ),
            .ltout(\U712_CHIP_RAM.N_323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_7_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_7_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_7_8_1 .LUT_INIT=16'b0101111101010000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_7_8_1  (
            .in0(N__3840),
            .in1(_gnd_net_),
            .in2(N__3726),
            .in3(N__4106),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8118),
            .ce(),
            .sr(N__9369));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILCLN6_LC_7_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILCLN6_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILCLN6_LC_7_8_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILCLN6_LC_7_8_3  (
            .in0(N__7773),
            .in1(N__3723),
            .in2(N__5103),
            .in3(N__6390),
            .lcout(\U712_CHIP_RAM.N_256_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_8_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_8_5  (
            .in0(N__6637),
            .in1(N__3708),
            .in2(_gnd_net_),
            .in3(N__4155),
            .lcout(\U712_CHIP_RAM.N_220 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_7_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_7_8_6 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_7_8_6  (
            .in0(N__5616),
            .in1(N__5480),
            .in2(_gnd_net_),
            .in3(N__4860),
            .lcout(\U712_CHIP_RAM.N_216 ),
            .ltout(\U712_CHIP_RAM.N_216_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_8_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(N__4105),
            .in2(N__3702),
            .in3(N__4658),
            .lcout(\U712_CHIP_RAM.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_0_LC_7_9_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_7_9_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_7_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3879),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8121),
            .ce(),
            .sr(N__9364));
    defparam \U712_REG_SM.C3_SYNC_1_LC_7_9_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_7_9_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_7_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4364),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8121),
            .ce(),
            .sr(N__9364));
    defparam \U712_REG_SM.C3_SYNC_2_LC_7_9_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_2_LC_7_9_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_2_LC_7_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_2_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4912),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8121),
            .ce(),
            .sr(N__9364));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_7_10_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_7_10_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_7_10_5  (
            .in0(N__6123),
            .in1(N__6269),
            .in2(_gnd_net_),
            .in3(N__8496),
            .lcout(\U712_BYTE_ENABLE.N_275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_10_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_10_7  (
            .in0(N__6846),
            .in1(N__6722),
            .in2(_gnd_net_),
            .in3(N__6438),
            .lcout(\U712_CHIP_RAM.N_213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_0_a3_LC_8_3_7 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_0_a3_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_0_a3_LC_8_3_7 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_0_a3_LC_8_3_7  (
            .in0(N__8543),
            .in1(N__6216),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_8_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_8_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_8_4_0  (
            .in0(N__3819),
            .in1(N__3801),
            .in2(_gnd_net_),
            .in3(N__8339),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_8_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_8_4_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_8_4_1  (
            .in0(N__8340),
            .in1(N__8552),
            .in2(N__3789),
            .in3(N__9240),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_8_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_8_4_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_8_4_3  (
            .in0(N__8337),
            .in1(N__3786),
            .in2(_gnd_net_),
            .in3(N__3768),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_8_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_8_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_8_4_4  (
            .in0(N__3981),
            .in1(N__3963),
            .in2(_gnd_net_),
            .in3(N__8338),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_8_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_8_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_8_4_6  (
            .in0(N__3942),
            .in1(N__3930),
            .in2(_gnd_net_),
            .in3(N__8336),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_1_1_LC_8_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_1_1_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_1_1_LC_8_5_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_1_1_LC_8_5_1  (
            .in0(N__4172),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5399),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_8_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_8_5_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_8_5_2  (
            .in0(N__4521),
            .in1(N__3915),
            .in2(N__3906),
            .in3(N__3894),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8104),
            .ce(N__4026),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINN5O1_LC_8_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINN5O1_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINN5O1_LC_8_5_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINN5O1_LC_8_5_4  (
            .in0(N__5623),
            .in1(N__6608),
            .in2(_gnd_net_),
            .in3(N__4146),
            .lcout(\U712_CHIP_RAM.N_300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_8_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_8_5_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(N__4660),
            .in2(_gnd_net_),
            .in3(N__4868),
            .lcout(\U712_CHIP_RAM.N_177 ),
            .ltout(\U712_CHIP_RAM.N_177_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNINB8M4_0_LC_8_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNINB8M4_0_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNINB8M4_0_LC_8_5_6 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNINB8M4_0_LC_8_5_6  (
            .in0(N__5624),
            .in1(N__3903),
            .in2(N__3897),
            .in3(N__6550),
            .lcout(\U712_CHIP_RAM.N_223 ),
            .ltout(\U712_CHIP_RAM.N_223_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI63MN7_2_LC_8_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI63MN7_2_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI63MN7_2_LC_8_5_7 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI63MN7_2_LC_8_5_7  (
            .in0(N__4171),
            .in1(N__3888),
            .in2(N__3882),
            .in3(N__4869),
            .lcout(\U712_CHIP_RAM.N_42_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_8_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_8_6_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_8_6_0  (
            .in0(N__6535),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6650),
            .lcout(\U712_CHIP_RAM.N_311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_6_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__6635),
            .in2(_gnd_net_),
            .in3(N__6534),
            .lcout(\U712_CHIP_RAM.N_187 ),
            .ltout(\U712_CHIP_RAM.N_187_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_8_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_8_6_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_8_6_2  (
            .in0(N__7782),
            .in1(N__4794),
            .in2(N__4044),
            .in3(N__4670),
            .lcout(\U712_CHIP_RAM.N_262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGELS1_2_LC_8_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGELS1_2_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGELS1_2_LC_8_6_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIGELS1_2_LC_8_6_3  (
            .in0(N__5596),
            .in1(N__7781),
            .in2(N__4870),
            .in3(N__5494),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILJN86_2_LC_8_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILJN86_2_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILJN86_2_LC_8_6_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNILJN86_2_LC_8_6_4  (
            .in0(N__6386),
            .in1(N__5100),
            .in2(N__4041),
            .in3(N__4776),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_264_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ3ENG_3_LC_8_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ3ENG_3_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ3ENG_3_LC_8_6_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ3ENG_3_LC_8_6_5  (
            .in0(N__4118),
            .in1(N__7783),
            .in2(N__4038),
            .in3(N__4035),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_8_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_8_6_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4029),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_6_7 .LUT_INIT=16'b1111001111100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_6_7  (
            .in0(N__4014),
            .in1(N__4543),
            .in2(N__7499),
            .in3(N__4005),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8107),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_7_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_7_0  (
            .in0(N__4253),
            .in1(N__7779),
            .in2(N__3999),
            .in3(N__4053),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8111),
            .ce(N__4221),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_8_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_8_7_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_8_7_1  (
            .in0(N__5609),
            .in1(N__3987),
            .in2(N__4788),
            .in3(N__4643),
            .lcout(\U712_CHIP_RAM.N_242 ),
            .ltout(\U712_CHIP_RAM.N_242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9NL8E_3_LC_8_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9NL8E_3_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9NL8E_3_LC_8_7_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9NL8E_3_LC_8_7_2  (
            .in0(N__4119),
            .in1(N__4075),
            .in2(N__4185),
            .in3(N__7780),
            .lcout(\U712_CHIP_RAM.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOO5O1_LC_8_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOO5O1_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOO5O1_LC_8_7_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOO5O1_LC_8_7_3  (
            .in0(N__6615),
            .in1(N__5490),
            .in2(_gnd_net_),
            .in3(N__5385),
            .lcout(\U712_CHIP_RAM.N_319 ),
            .ltout(\U712_CHIP_RAM.N_319_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINL0R5_LC_8_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINL0R5_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINL0R5_LC_8_7_4 .LUT_INIT=16'b1111001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINL0R5_LC_8_7_4  (
            .in0(N__4173),
            .in1(N__4154),
            .in2(N__4122),
            .in3(N__4688),
            .lcout(\U712_CHIP_RAM.N_322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_3_LC_8_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_3_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_3_LC_8_7_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_3_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(N__4642),
            .in2(_gnd_net_),
            .in3(N__4851),
            .lcout(\U712_CHIP_RAM.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_8_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_8_7_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_8_7_6  (
            .in0(N__4852),
            .in1(N__5479),
            .in2(N__5627),
            .in3(N__4101),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_7_7 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_7_7  (
            .in0(N__4076),
            .in1(N__4515),
            .in2(N__4266),
            .in3(N__4062),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8111),
            .ce(N__4221),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_8_8_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_8_8_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__5608),
            .in2(_gnd_net_),
            .in3(N__9093),
            .lcout(\U712_CHIP_RAM.DBENn_7_0 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_1  (
            .in0(N__4257),
            .in1(N__5481),
            .in2(_gnd_net_),
            .in3(N__4056),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__8115),
            .ce(N__4220),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__4864),
            .in2(_gnd_net_),
            .in3(N__4047),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3  (
            .in0(N__4258),
            .in1(N__4659),
            .in2(_gnd_net_),
            .in3(N__4278),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__8115),
            .ce(N__4220),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4  (
            .in0(N__4254),
            .in1(N__4724),
            .in2(_gnd_net_),
            .in3(N__4275),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__8115),
            .ce(N__4220),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5  (
            .in0(N__4259),
            .in1(N__4737),
            .in2(_gnd_net_),
            .in3(N__4272),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__8115),
            .ce(N__4220),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6  (
            .in0(N__4255),
            .in1(N__4749),
            .in2(_gnd_net_),
            .in3(N__4269),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__8115),
            .ce(N__4220),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7  (
            .in0(N__4710),
            .in1(N__4256),
            .in2(_gnd_net_),
            .in3(N__4224),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8115),
            .ce(N__4220),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_9_0 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_9_0  (
            .in0(N__7760),
            .in1(N__6304),
            .in2(N__6900),
            .in3(N__6325),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_207_i_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_9_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_9_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_9_1  (
            .in0(N__9414),
            .in1(_gnd_net_),
            .in2(N__4209),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.N_207_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_9_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_9_2 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_9_2 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_9_2  (
            .in0(N__7759),
            .in1(N__6305),
            .in2(_gnd_net_),
            .in3(N__6326),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8119),
            .ce(N__4194),
            .sr(N__9354));
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_0_2_LC_8_9_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_0_2_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_0_2_LC_8_9_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI9DCD1_0_2_LC_8_9_6  (
            .in0(N__4381),
            .in1(N__4335),
            .in2(N__4313),
            .in3(N__4359),
            .lcout(\U712_REG_SM.N_185 ),
            .ltout(\U712_REG_SM.N_185_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_8_9_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_8_9_7 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__4941),
            .in2(N__4422),
            .in3(N__4903),
            .lcout(\U712_REG_SM.N_188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_0_LC_8_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_8_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_8_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4419),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8122),
            .ce(),
            .sr(N__9346));
    defparam \U712_REG_SM.C1_SYNC_1_LC_8_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_8_10_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_8_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_8_10_1  (
            .in0(N__4312),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8122),
            .ce(),
            .sr(N__9346));
    defparam \U712_REG_SM.C1_SYNC_2_LC_8_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_2_LC_8_10_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_2_LC_8_10_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \U712_REG_SM.C1_SYNC_2_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__4338),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8122),
            .ce(),
            .sr(N__9346));
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_8_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_8_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_8_10_3  (
            .in0(N__4382),
            .in1(N__4336),
            .in2(N__4314),
            .in3(N__4360),
            .lcout(\U712_REG_SM.N_197 ),
            .ltout(\U712_REG_SM.N_197_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_8_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_8_10_4 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_8_10_4  (
            .in0(N__4911),
            .in1(_gnd_net_),
            .in2(N__4386),
            .in3(N__4948),
            .lcout(\U712_REG_SM.N_209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIFFTG1_2_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIFFTG1_2_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIFFTG1_2_LC_8_10_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIFFTG1_2_LC_8_10_5  (
            .in0(N__4383),
            .in1(N__4910),
            .in2(N__4368),
            .in3(N__4942),
            .lcout(),
            .ltout(\U712_REG_SM.DS_EN_0_sqmuxa_0_a2_0_a3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_8_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_8_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_8_10_6  (
            .in0(N__4286),
            .in1(N__4337),
            .in2(N__4317),
            .in3(N__4311),
            .lcout(\U712_REG_SM.DS_EN_0_sqmuxa ),
            .ltout(\U712_REG_SM.DS_EN_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_8_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_8_10_7 .LUT_INIT=16'b0000110000001110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_8_10_7  (
            .in0(N__5817),
            .in1(N__4287),
            .in2(N__4290),
            .in3(N__5201),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8122),
            .ce(),
            .sr(N__9346));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_9_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_9_4_0 .LUT_INIT=16'b0000000001100111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_9_4_0  (
            .in0(N__7674),
            .in1(N__8330),
            .in2(N__7504),
            .in3(N__8702),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_9_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_9_4_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_9_4_1  (
            .in0(N__9417),
            .in1(_gnd_net_),
            .in2(N__4491),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_9_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_9_4_2 .LUT_INIT=16'b1011111110110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_9_4_2  (
            .in0(N__4488),
            .in1(N__7426),
            .in2(N__8576),
            .in3(N__8889),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_9_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_9_4_4 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_9_4_4  (
            .in0(N__4487),
            .in1(N__7425),
            .in2(N__8577),
            .in3(N__8888),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_4_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_4_5  (
            .in0(N__8334),
            .in1(N__4467),
            .in2(N__8578),
            .in3(N__8751),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_9_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_9_4_6 .LUT_INIT=16'b0000010011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_9_4_6  (
            .in0(N__8548),
            .in1(N__8636),
            .in2(N__8225),
            .in3(N__8335),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_9_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_9_4_7 .LUT_INIT=16'b0000111111101111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_9_4_7  (
            .in0(N__8637),
            .in1(N__8544),
            .in2(N__8364),
            .in3(N__8210),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_5_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_5_0  (
            .in0(N__8341),
            .in1(N__4461),
            .in2(_gnd_net_),
            .in3(N__4443),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_5_1 .LUT_INIT=16'b1010101000001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_5_1  (
            .in0(N__6631),
            .in1(N__4872),
            .in2(N__5508),
            .in3(N__5626),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_5_2 .LUT_INIT=16'b1111111000110010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_5_2  (
            .in0(N__4529),
            .in1(N__4544),
            .in2(N__4425),
            .in3(N__7673),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8101),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_5_3 .LUT_INIT=16'b1111010111100100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_5_3  (
            .in0(N__4545),
            .in1(N__4530),
            .in2(N__8719),
            .in3(N__4509),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8101),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_0_LC_9_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_0_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_0_LC_9_5_5 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_0_LC_9_5_5  (
            .in0(N__7672),
            .in1(_gnd_net_),
            .in2(N__7495),
            .in3(N__8342),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_5_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(N__7671),
            .in2(_gnd_net_),
            .in3(N__7476),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_9_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_9_5_7 .LUT_INIT=16'b0000000011010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_9_5_7  (
            .in0(N__6485),
            .in1(N__6443),
            .in2(N__6638),
            .in3(N__5625),
            .lcout(\U712_CHIP_RAM.N_236 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_0  (
            .in0(N__6785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5607),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_6_1 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_6_1  (
            .in0(N__5606),
            .in1(N__5493),
            .in2(N__5398),
            .in3(N__4854),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_6_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_6_2  (
            .in0(N__5492),
            .in1(N__5605),
            .in2(_gnd_net_),
            .in3(N__5386),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_9_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_9_6_3 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_9_6_3  (
            .in0(N__4503),
            .in1(N__4671),
            .in2(N__4497),
            .in3(N__4777),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_LC_9_6_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_LC_9_6_4  (
            .in0(N__9415),
            .in1(_gnd_net_),
            .in2(N__4494),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_9_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_9_6_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(N__5491),
            .in2(_gnd_net_),
            .in3(N__4853),
            .lcout(\U712_CHIP_RAM.N_198_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_7_0 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__5390),
            .in2(N__4787),
            .in3(N__4677),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_7_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_7_1  (
            .in0(N__4748),
            .in1(N__4736),
            .in2(N__4725),
            .in3(N__4709),
            .lcout(\U712_CHIP_RAM.N_355 ),
            .ltout(\U712_CHIP_RAM.N_355_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_9_7_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4698),
            .in3(N__5582),
            .lcout(\U712_CHIP_RAM.N_321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_9_7_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_9_7_3  (
            .in0(N__5583),
            .in1(N__5495),
            .in2(_gnd_net_),
            .in3(N__4654),
            .lcout(\U712_CHIP_RAM.N_235 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_7_4 .LUT_INIT=16'b1111111110101011;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_7_4  (
            .in0(N__5496),
            .in1(N__5584),
            .in2(N__4669),
            .in3(N__6542),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CPU_TACK_8_iv_i_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_7_5 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_7_5  (
            .in0(N__4587),
            .in1(N__8517),
            .in2(N__4569),
            .in3(N__5397),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_117_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_9_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_9_7_6 .LUT_INIT=16'b1010101010001011;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_9_7_6  (
            .in0(N__5112),
            .in1(N__4566),
            .in2(N__4554),
            .in3(N__4551),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8108),
            .ce(),
            .sr(N__9365));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_7_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_7_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_9_7_7  (
            .in0(N__5972),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5111),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861_1_LC_9_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861_1_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861_1_LC_9_8_1 .LUT_INIT=16'b0000111101111111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861_1_LC_9_8_1  (
            .in0(N__5876),
            .in1(N__5961),
            .in2(N__5043),
            .in3(N__5027),
            .lcout(\U712_CHIP_RAM.REFRESH_SYNC_RNI5J861Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_8_4 .LUT_INIT=16'b0000001110101011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_8_4  (
            .in0(N__5042),
            .in1(N__5265),
            .in2(N__5067),
            .in3(N__8562),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8112),
            .ce(),
            .sr(N__9355));
    defparam DBR_SYNC_1_LC_9_8_5.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_9_8_5.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_9_8_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 DBR_SYNC_1_LC_9_8_5 (
            .in0(N__5142),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8112),
            .ce(),
            .sr(N__9355));
    defparam \U712_REG_SM.C3_SYNC_RNIBM0G2_2_LC_9_8_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIBM0G2_2_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIBM0G2_2_LC_9_8_6 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIBM0G2_2_LC_9_8_6  (
            .in0(N__5028),
            .in1(N__5141),
            .in2(_gnd_net_),
            .in3(N__5940),
            .lcout(\U712_REG_SM.N_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_9_1 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_9_9_1  (
            .in0(N__5187),
            .in1(N__5157),
            .in2(N__5019),
            .in3(N__5312),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8116),
            .ce(),
            .sr(N__9347));
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_9_9_2 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_9_9_2  (
            .in0(N__4950),
            .in1(N__5015),
            .in2(N__4920),
            .in3(N__5007),
            .lcout(\U712_REG_SM.N_215 ),
            .ltout(\U712_REG_SM.N_215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_1_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_1_LC_9_9_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_1_LC_9_9_3 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \U712_REG_SM.REGENn_1_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__4963),
            .in2(N__5001),
            .in3(N__5172),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8116),
            .ce(),
            .sr(N__9347));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_9_9_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_9_9_4  (
            .in0(N__4949),
            .in1(N__4913),
            .in2(_gnd_net_),
            .in3(N__4878),
            .lcout(\U712_REG_SM.N_204 ),
            .ltout(\U712_REG_SM.N_204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_9_9_5 .LUT_INIT=16'b0000000010101110;
    LogicCell40 \U712_REG_SM.DS_EN_LC_9_9_5  (
            .in0(N__6032),
            .in1(N__5279),
            .in2(N__5319),
            .in3(N__5171),
            .lcout(DS_ENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8116),
            .ce(),
            .sr(N__9347));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_9_7 .LUT_INIT=16'b0010111000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_9_9_7  (
            .in0(N__5865),
            .in1(N__5278),
            .in2(N__5295),
            .in3(N__5846),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8116),
            .ce(),
            .sr(N__9347));
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_9_10_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_GO_LC_9_10_0  (
            .in0(N__5155),
            .in1(N__5210),
            .in2(N__5316),
            .in3(N__5189),
            .lcout(\U712_REG_SM.REG_CYCLE_GOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8120),
            .ce(),
            .sr(N__9340));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_10_1 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_9_10_1  (
            .in0(N__5311),
            .in1(N__5280),
            .in2(_gnd_net_),
            .in3(N__5294),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8120),
            .ce(),
            .sr(N__9340));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_10_2 .LUT_INIT=16'b0000010111001101;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_9_10_2  (
            .in0(N__5261),
            .in1(N__5190),
            .in2(N__5235),
            .in3(N__5211),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8120),
            .ce(),
            .sr(N__9340));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_9_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_9_10_3 .LUT_INIT=16'b1010000010101000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_9_10_3  (
            .in0(N__5202),
            .in1(N__5918),
            .in2(N__5823),
            .in3(N__5941),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8120),
            .ce(),
            .sr(N__9340));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_10_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_10_6 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_9_10_6  (
            .in0(N__5156),
            .in1(N__5188),
            .in2(_gnd_net_),
            .in3(N__5170),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8120),
            .ce(),
            .sr(N__9340));
    defparam DBR_SYNC_0_LC_9_11_2.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_9_11_2.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_9_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_9_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8840),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8123),
            .ce(),
            .sr(N__9338));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_10_2_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_10_2_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_10_2_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_10_2_5  (
            .in0(N__7682),
            .in1(N__8394),
            .in2(N__7512),
            .in3(N__8718),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8092),
            .ce(N__7985),
            .sr(N__9392));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_4_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_10_4_4  (
            .in0(N__5793),
            .in1(N__5784),
            .in2(_gnd_net_),
            .in3(N__5778),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8099),
            .ce(N__7984),
            .sr(N__9377));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_10_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_10_4_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_10_4_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_10_4_7  (
            .in0(N__5754),
            .in1(N__5748),
            .in2(_gnd_net_),
            .in3(N__5634),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8099),
            .ce(N__7984),
            .sr(N__9377));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_5_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_5_1  (
            .in0(N__5721),
            .in1(N__8358),
            .in2(_gnd_net_),
            .in3(N__5706),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_10_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_10_5_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_10_5_2  (
            .in0(N__8359),
            .in1(N__8530),
            .in2(N__5694),
            .in3(N__8973),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_5_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_5_5  (
            .in0(N__5691),
            .in1(N__8357),
            .in2(_gnd_net_),
            .in3(N__5676),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_5_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_5_6  (
            .in0(N__5658),
            .in1(N__8531),
            .in2(_gnd_net_),
            .in3(N__9231),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_324_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_7 .LUT_INIT=16'b0011001111110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_7  (
            .in0(_gnd_net_),
            .in1(N__8360),
            .in2(N__5637),
            .in3(N__8224),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_10_6_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_10_6_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_LC_10_6_0  (
            .in0(N__5628),
            .in1(N__5507),
            .in2(_gnd_net_),
            .in3(N__5403),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8102),
            .ce(N__5328),
            .sr(N__9366));
    defparam \U712_CHIP_RAM.DBENn_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_10_7_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_10_7_1 .LUT_INIT=16'b0000001011111110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_10_7_1  (
            .in0(N__7243),
            .in1(N__6006),
            .in2(N__6504),
            .in3(N__5997),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8105),
            .ce(),
            .sr(N__9356));
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_10_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_10_7_4 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_LC_10_7_4  (
            .in0(N__7207),
            .in1(N__6502),
            .in2(_gnd_net_),
            .in3(N__5985),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8105),
            .ce(),
            .sr(N__9356));
    defparam \U712_REG_SM.REG_TACK_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_10_7_7 .LUT_INIT=16'b1101100011011100;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_10_7_7  (
            .in0(N__5821),
            .in1(N__5917),
            .in2(N__5976),
            .in3(N__5955),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8105),
            .ce(),
            .sr(N__9356));
    defparam \U712_CHIP_RAM.REFRESH_SYNC_1_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_1_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_1_LC_10_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_SYNC_1_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5877),
            .lcout(\U712_CHIP_RAM.REFRESH_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8109),
            .ce(),
            .sr(N__9348));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_10_8_1 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_10_8_1  (
            .in0(N__5864),
            .in1(N__5842),
            .in2(N__5919),
            .in3(N__5954),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8109),
            .ce(),
            .sr(N__9348));
    defparam \U712_CHIP_RAM.REFRESH_SYNC_0_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_0_LC_10_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_0_LC_10_8_3 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \U712_CHIP_RAM.REFRESH_SYNC_0_LC_10_8_3  (
            .in0(N__5895),
            .in1(N__8948),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.REFRESH_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8109),
            .ce(),
            .sr(N__9348));
    defparam \U712_REG_SM.REG_CYCLE_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_10_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_10_8_5 .LUT_INIT=16'b1010101011001110;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_10_8_5  (
            .in0(N__5863),
            .in1(N__6199),
            .in2(N__5850),
            .in3(N__5822),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8109),
            .ce(),
            .sr(N__9348));
    defparam \U712_CHIP_RAM.REFRESH_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_8_7 .LUT_INIT=16'b1111001111111011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_10_8_7  (
            .in0(N__7887),
            .in1(N__6999),
            .in2(N__7818),
            .in3(N__6987),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8109),
            .ce(),
            .sr(N__9348));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_10_9_3 .LUT_INIT=16'b1100100011111000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_10_9_3  (
            .in0(N__6980),
            .in1(N__6941),
            .in2(N__6306),
            .in3(N__6333),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8113),
            .ce(),
            .sr(N__9341));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_9_4 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_9_4 .LUT_INIT=16'b1111110011110100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_10_9_4  (
            .in0(N__6940),
            .in1(N__6344),
            .in2(N__7338),
            .in3(N__6981),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8113),
            .ce(),
            .sr(N__9341));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_9_5 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_9_5 .LUT_INIT=16'b0011001000110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_10_9_5  (
            .in0(N__7305),
            .in1(N__6939),
            .in2(N__6899),
            .in3(N__6332),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8113),
            .ce(),
            .sr(N__9341));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_10_10_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_10_10_2  (
            .in0(N__6138),
            .in1(N__6285),
            .in2(_gnd_net_),
            .in3(N__8569),
            .lcout(\U712_BYTE_ENABLE.N_271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_10_10_3 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_10_10_3  (
            .in0(N__6283),
            .in1(N__6136),
            .in2(N__8583),
            .in3(N__6241),
            .lcout(\U712_BYTE_ENABLE.N_277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_10_10_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_10_10_5 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_10_10_5  (
            .in0(N__6284),
            .in1(N__6137),
            .in2(N__8584),
            .in3(N__6242),
            .lcout(\U712_BYTE_ENABLE.N_273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_LC_10_10_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_LC_10_10_7 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_LC_10_10_7  (
            .in0(N__8570),
            .in1(N__6243),
            .in2(_gnd_net_),
            .in3(N__6084),
            .lcout(\U712_BYTE_ENABLE.N_270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_10_15_7 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_10_15_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_10_15_7  (
            .in0(N__7226),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6212),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_10_17_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_10_17_0 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_10_17_0  (
            .in0(N__6044),
            .in1(N__6124),
            .in2(_gnd_net_),
            .in3(N__6073),
            .lcout(un1_LDSn_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_10_17_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_10_17_7 .LUT_INIT=16'b1010000011111111;
    LogicCell40 \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_10_17_7  (
            .in0(N__6125),
            .in1(_gnd_net_),
            .in2(N__6080),
            .in3(N__6045),
            .lcout(un1_UDSn_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_10_18_3 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_10_18_3 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_10_18_3  (
            .in0(N__6721),
            .in1(N__6842),
            .in2(_gnd_net_),
            .in3(N__7227),
            .lcout(N_212),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_11_2_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_2_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_2_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_2_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_3_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_3_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_3_6 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_11_3_6  (
            .in0(N__8182),
            .in1(N__8787),
            .in2(N__8257),
            .in3(N__6744),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8093),
            .ce(N__8015),
            .sr(N__9378));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_4 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_4  (
            .in0(N__6750),
            .in1(N__8572),
            .in2(N__8398),
            .in3(N__8964),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_5_0 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_5_0  (
            .in0(N__8571),
            .in1(N__9222),
            .in2(N__8393),
            .in3(N__6738),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBDIR_LC_11_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_11_6_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_11_6_1 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_11_6_1  (
            .in0(N__6729),
            .in1(N__6503),
            .in2(_gnd_net_),
            .in3(N__6668),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8100),
            .ce(),
            .sr(N__9357));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_11_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_11_7_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_11_7_0  (
            .in0(N__6413),
            .in1(N__6657),
            .in2(N__6639),
            .in3(N__6551),
            .lcout(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_7_4 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_7_4  (
            .in0(N__6414),
            .in1(N__7206),
            .in2(N__6912),
            .in3(N__6993),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8103),
            .ce(),
            .sr(N__9349));
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_11_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_11_7_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIRILU_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__6468),
            .in2(_gnd_net_),
            .in3(N__6412),
            .lcout(\U712_CHIP_RAM.N_305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__7835),
            .in2(_gnd_net_),
            .in3(N__7850),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_8_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_8_3  (
            .in0(N__7028),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6923),
            .lcout(\U712_CHIP_RAM.un5_DMA_CYCLE_START_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_4 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_4  (
            .in0(N__7901),
            .in1(N__7352),
            .in2(N__7869),
            .in3(N__7367),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_9_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7317),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8110),
            .ce(),
            .sr(N__9339));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_9_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_9_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__6979),
            .in2(_gnd_net_),
            .in3(N__6942),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8110),
            .ce(),
            .sr(N__9339));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_9_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7029),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8110),
            .ce(),
            .sr(N__9339));
    defparam \U712_CHIP_RAM.CAS_SYNC_2_LC_11_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_2_LC_11_9_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_2_LC_11_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_2_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6924),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8110),
            .ce(),
            .sr(N__9339));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__7334),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8110),
            .ce(),
            .sr(N__9339));
    defparam \U712_BYTE_ENABLE.N_148_i_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_148_i_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_148_i_LC_11_10_0 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \U712_BYTE_ENABLE.N_148_i_LC_11_10_0  (
            .in0(N__7185),
            .in1(N__6879),
            .in2(N__7062),
            .in3(N__7146),
            .lcout(N_148_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_10_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_10_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__7333),
            .in2(_gnd_net_),
            .in3(N__7316),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0_0_LC_11_10_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0_0_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0_0_LC_11_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0_0_LC_11_10_2  (
            .in0(N__7259),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7219),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0 ),
            .ltout(\U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_171_i_LC_11_10_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_171_i_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_171_i_LC_11_10_3 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_171_i_LC_11_10_3  (
            .in0(N__7299),
            .in1(N__7149),
            .in2(N__7290),
            .in3(N__7061),
            .lcout(N_171_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0_LC_11_10_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0_LC_11_10_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0_LC_11_10_4  (
            .in0(N__7258),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7218),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0 ),
            .ltout(\U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_150_i_LC_11_10_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_150_i_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_150_i_LC_11_10_5 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_150_i_LC_11_10_5  (
            .in0(N__7147),
            .in1(N__7179),
            .in2(N__7173),
            .in3(N__7091),
            .lcout(N_150_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_172_i_LC_11_10_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_172_i_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_172_i_LC_11_10_7 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_172_i_LC_11_10_7  (
            .in0(N__7148),
            .in1(N__7131),
            .in2(N__7125),
            .in3(N__7092),
            .lcout(N_172_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_11_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_11_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_11_11_4  (
            .in0(N__7085),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7049),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8117),
            .ce(),
            .sr(N__9337));
    defparam \U712_CHIP_RAM.WEn_LC_12_2_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_12_2_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_12_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_12_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7508),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8088),
            .ce(),
            .sr(N__9375));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_3_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_3_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_3_1  (
            .in0(N__8386),
            .in1(N__8539),
            .in2(N__7629),
            .in3(N__7911),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496_1_LC_12_3_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496_1_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496_1_LC_12_3_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496_1_LC_12_3_6  (
            .in0(_gnd_net_),
            .in1(N__8538),
            .in2(_gnd_net_),
            .in3(N__8385),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_4_0 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_12_4_0  (
            .in0(N__8184),
            .in1(N__8245),
            .in2(N__9522),
            .in3(N__7614),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8091),
            .ce(N__8000),
            .sr(N__9363));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_4_1 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_12_4_1  (
            .in0(N__8183),
            .in1(N__9174),
            .in2(N__8256),
            .in3(N__7584),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8091),
            .ce(N__8000),
            .sr(N__9363));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_4_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_4_6 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_12_4_6  (
            .in0(N__7551),
            .in1(N__7439),
            .in2(N__8588),
            .in3(N__9162),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8091),
            .ce(N__8000),
            .sr(N__9363));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_12_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_12_5_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_12_5_2  (
            .in0(N__7681),
            .in1(N__8356),
            .in2(N__8720),
            .in3(N__7500),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_6_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_12_6_0  (
            .in0(N__7440),
            .in1(N__7407),
            .in2(N__8589),
            .in3(N__8922),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8095),
            .ce(N__8016),
            .sr(N__9345));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_8_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_8_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(N__7368),
            .in2(_gnd_net_),
            .in3(N__7356),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_12_8_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__8865),
            .ce(),
            .sr(N__7800));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_8_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_8_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__7353),
            .in2(_gnd_net_),
            .in3(N__7341),
            .lcout(\U712_CHIP_RAM.REFRESH5lto1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__8865),
            .ce(),
            .sr(N__7800));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_8_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_8_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(N__7902),
            .in2(_gnd_net_),
            .in3(N__7890),
            .lcout(\U712_CHIP_RAM.REFRESH5lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__8865),
            .ce(),
            .sr(N__7800));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_8_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_8_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(N__7886),
            .in2(_gnd_net_),
            .in3(N__7872),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__8865),
            .ce(),
            .sr(N__7800));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_8_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_8_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(N__7868),
            .in2(_gnd_net_),
            .in3(N__7854),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__8865),
            .ce(),
            .sr(N__7800));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_8_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_8_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(N__7851),
            .in2(_gnd_net_),
            .in3(N__7839),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__8865),
            .ce(),
            .sr(N__7800));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_8_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_8_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_8_6  (
            .in0(_gnd_net_),
            .in1(N__7836),
            .in2(_gnd_net_),
            .in3(N__7824),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__8865),
            .ce(),
            .sr(N__7800));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_8_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_8_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__7814),
            .in2(_gnd_net_),
            .in3(N__7821),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8865),
            .ce(),
            .sr(N__7800));
    defparam RESETn_ibuf_RNIM9SF_LC_12_11_0.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_11_0.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_11_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7728),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RASn_LC_13_1_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_13_1_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_13_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_13_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7686),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8089),
            .ce(),
            .sr(N__9393));
    defparam \U712_CHIP_RAM.CASn_LC_13_1_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_13_1_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_13_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_13_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8399),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8089),
            .ce(),
            .sr(N__9393));
    defparam \U712_CHIP_RAM.CRCSn_LC_13_1_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_1_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_13_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8721),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8089),
            .ce(),
            .sr(N__9393));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_2_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_2_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_2_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_13_2_2  (
            .in0(N__8185),
            .in1(N__8793),
            .in2(N__8262),
            .in3(N__8658),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8090),
            .ce(N__8008),
            .sr(N__9385));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_3_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_3_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7947),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9500),
            .ce(N__9469),
            .sr(N__9379));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_4_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_4_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_13_4_2  (
            .in0(N__8186),
            .in1(N__9009),
            .in2(N__8258),
            .in3(N__8622),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8094),
            .ce(N__8007),
            .sr(N__9370));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_4_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_4_5  (
            .in0(N__8579),
            .in1(N__8412),
            .in2(N__8400),
            .in3(N__9126),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_4_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_4_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_13_4_6  (
            .in0(N__8252),
            .in1(N__8187),
            .in2(N__8151),
            .in3(N__9567),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8094),
            .ce(N__8007),
            .sr(N__9370));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7940),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__9083),
            .sr(N__9367));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_5_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8916),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__9083),
            .sr(N__9367));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9213),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__9083),
            .sr(N__9367));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_13_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_13_6_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_13_6_3  (
            .in0(N__8952),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9498),
            .ce(N__9451),
            .sr(N__9358));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8912),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9498),
            .ce(N__9451),
            .sr(N__9358));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_13_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_13_7_4 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_13_7_4  (
            .in0(N__9413),
            .in1(N__8841),
            .in2(_gnd_net_),
            .in3(N__8874),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_13_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_13_8_1 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_13_8_1  (
            .in0(N__9412),
            .in1(N__8836),
            .in2(_gnd_net_),
            .in3(N__9507),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_3_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_3_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9117),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9502),
            .ce(N__9474),
            .sr(N__9386));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_3_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_3_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_3_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_3_5  (
            .in0(N__8778),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9502),
            .ce(N__9474),
            .sr(N__9386));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_4_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8777),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__9082),
            .sr(N__9380));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_4_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9033),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__9082),
            .sr(N__9380));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9555),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__9081),
            .sr(N__9371));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9000),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__9081),
            .sr(N__9371));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_6_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_6_5  (
            .in0(N__9212),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9499),
            .ce(N__9467),
            .sr(N__9368));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_6_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_6_7  (
            .in0(N__9150),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9499),
            .ce(N__9467),
            .sr(N__9368));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9149),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__9084),
            .sr(N__9359));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_14_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_14_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_14_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9116),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__9065),
            .sr(N__9350));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_4_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_4_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_4_4  (
            .in0(N__9032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9503),
            .ce(N__9468),
            .sr(N__9387));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8996),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9501),
            .ce(N__9470),
            .sr(N__9381));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9551),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9501),
            .ce(N__9470),
            .sr(N__9381));
endmodule // U712_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 25 2025 11:06:30

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    TT : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(31 downto 1);
    TICK50 : out std_logic;
    nROMEN : out std_logic;
    nCIACS1 : out std_logic;
    TICK60 : out std_logic;
    CLKCIA : out std_logic;
    CLK6 : in std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    TSn : in std_logic;
    nBUFEN : out std_logic;
    nREGSPACE : out std_logic;
    nRAMSPACE : out std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    TACKn : inout std_logic;
    nCIACS0 : out std_logic;
    PORTSIZE : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__6284\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2586\ : std_logic;
signal \N__2583\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2566\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2526\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2446\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_17\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U409_CIA.g0Z0Z_8_cascade_\ : std_logic;
signal \U409_CIA.g0Z0Z_11\ : std_logic;
signal \A_c_25\ : std_logic;
signal \A_c_24\ : std_logic;
signal \A_c_26\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \A_c_31\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7_cascade_\ : std_logic;
signal \U409_CIA.g0Z0Z_10\ : std_logic;
signal \U409_CIA.g0Z0Z_2_cascade_\ : std_logic;
signal \A_c_29\ : std_logic;
signal \A_c_28\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_30\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_10\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEm_6\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEm_3\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_CIA.N_9_cascade_\ : std_logic;
signal \U409_CIA.N_20_cascade_\ : std_logic;
signal \U409_CIA.CLKCIA8_0_a2_0\ : std_logic;
signal \U409_CIA.CLKCIA6_0_a2_1\ : std_logic;
signal \U409_CIA.CLKCIAZ0_cascade_\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a2_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nREGSPACE_i\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nCIACS1_i\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nCIACS0_i\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \CIA_ENABLEm\ : std_logic;
signal \A_c_22\ : std_logic;
signal \A_c_23\ : std_logic;
signal \A_c_21\ : std_logic;
signal \AUTOVECTORm\ : std_logic;
signal \ROMENm_i\ : std_logic;
signal \U409_ADDRESS_DECODE.LOWROMZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.HIROMZ0\ : std_logic;
signal \ROMENm\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\ : std_logic;
signal \U409_TRANSFER_ACK.m9_am_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.i6_mux_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0\ : std_logic;
signal \OVL_c\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \U409_CIA.g0Z0Z_14\ : std_logic;
signal \U409_CIA.g0Z0Z_13\ : std_logic;
signal \U409_CIA.CIA_HOLDZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\ : std_logic;
signal \U409_TICK.TICK603_8_cascade_\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.TICK603_11\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \U409_TICK.TICK603_10_cascade_\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \U409_TRANSFER_ACK.N_107\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_107_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.m9_bm\ : std_logic;
signal \U409_TRANSFER_ACK.N_4\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \CLKCIA_c\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \bfn_12_7_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_EN_e_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_OUTnC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_EN_iC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\ : std_logic;
signal \TACK_EN_i\ : std_logic;
signal \N_373_i\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \nBUFEN_c\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \CLKCIA_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \nCIACS0_wire\ : std_logic;
signal \nCIACS1_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \nRAMSPACE_wire\ : std_logic;
signal \nROMEN_wire\ : std_logic;
signal \nBUFEN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \nREGSPACE_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    \TT_wire\ <= TT;
    CLKCIA <= \CLKCIA_wire\;
    \A_wire\ <= A;
    nCIACS0 <= \nCIACS0_wire\;
    nCIACS1 <= \nCIACS1_wire\;
    \TSn_wire\ <= TSn;
    PORTSIZE <= \PORTSIZE_wire\;
    nRAMSPACE <= \nRAMSPACE_wire\;
    nROMEN <= \nROMEN_wire\;
    nBUFEN <= \nBUFEN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    nREGSPACE <= \nREGSPACE_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TICK60 <= \TICK60_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__5110\,
            RESETB => \N__4891\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6282\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6284\,
            DIN => \N__6283\,
            DOUT => \N__6282\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6284\,
            PADOUT => \N__6283\,
            PADIN => \N__6282\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6272\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6274\,
            DIN => \N__6273\,
            DOUT => \N__6272\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6274\,
            PADOUT => \N__6273\,
            PADIN => \N__6272\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6263\,
            DIN => \N__6262\,
            DOUT => \N__6261\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6263\,
            PADOUT => \N__6262\,
            PADIN => \N__6261\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKCIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6254\,
            DIN => \N__6253\,
            DOUT => \N__6252\,
            PACKAGEPIN => \CLKCIA_wire\
        );

    \CLKCIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6254\,
            PADOUT => \N__6253\,
            PADIN => \N__6252\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4948\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6245\,
            DIN => \N__6244\,
            DOUT => \N__6243\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6245\,
            PADOUT => \N__6244\,
            PADIN => \N__6243\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6236\,
            DIN => \N__6235\,
            DOUT => \N__6234\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6236\,
            PADOUT => \N__6235\,
            PADIN => \N__6234\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCIACS0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6227\,
            DIN => \N__6226\,
            DOUT => \N__6225\,
            PACKAGEPIN => \nCIACS0_wire\
        );

    \nCIACS0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6227\,
            PADOUT => \N__6226\,
            PADIN => \N__6225\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3076\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCIACS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6218\,
            DIN => \N__6217\,
            DOUT => \N__6216\,
            PACKAGEPIN => \nCIACS1_wire\
        );

    \nCIACS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6218\,
            PADOUT => \N__6217\,
            PADIN => \N__6216\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3109\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6209\,
            DIN => \N__6208\,
            DOUT => \N__6207\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6209\,
            PADOUT => \N__6208\,
            PADIN => \N__6207\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6200\,
            DIN => \N__6199\,
            DOUT => \N__6198\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6200\,
            PADOUT => \N__6199\,
            PADIN => \N__6198\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6191\,
            DIN => \N__6190\,
            DOUT => \N__6189\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6191\,
            PADOUT => \N__6190\,
            PADIN => \N__6189\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6182\,
            DIN => \N__6181\,
            DOUT => \N__6180\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6182\,
            PADOUT => \N__6181\,
            PADIN => \N__6180\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5878\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__5515\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6173\,
            DIN => \N__6172\,
            DOUT => \N__6171\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6173\,
            PADOUT => \N__6172\,
            PADIN => \N__6171\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6164\,
            DIN => \N__6163\,
            DOUT => \N__6162\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6164\,
            PADOUT => \N__6163\,
            PADIN => \N__6162\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6155\,
            DIN => \N__6154\,
            DOUT => \N__6153\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6155\,
            PADOUT => \N__6154\,
            PADIN => \N__6153\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6146\,
            DIN => \N__6145\,
            DOUT => \N__6144\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6146\,
            PADOUT => \N__6145\,
            PADIN => \N__6144\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2989\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nRAMSPACE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6137\,
            DIN => \N__6136\,
            DOUT => \N__6135\,
            PACKAGEPIN => \nRAMSPACE_wire\
        );

    \nRAMSPACE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6137\,
            PADOUT => \N__6136\,
            PADIN => \N__6135\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3574\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nROMEN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6128\,
            DIN => \N__6127\,
            DOUT => \N__6126\,
            PACKAGEPIN => \nROMEN_wire\
        );

    \nROMEN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6128\,
            PADOUT => \N__6127\,
            PADIN => \N__6126\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3883\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6119\,
            DIN => \N__6118\,
            DOUT => \N__6117\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6119\,
            PADOUT => \N__6118\,
            PADIN => \N__6117\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6110\,
            DIN => \N__6109\,
            DOUT => \N__6108\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6110\,
            PADOUT => \N__6109\,
            PADIN => \N__6108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nBUFEN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6101\,
            DIN => \N__6100\,
            DOUT => \N__6099\,
            PACKAGEPIN => \nBUFEN_wire\
        );

    \nBUFEN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6101\,
            PADOUT => \N__6100\,
            PADIN => \N__6099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5713\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6092\,
            DIN => \N__6091\,
            DOUT => \N__6090\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6092\,
            PADOUT => \N__6091\,
            PADIN => \N__6090\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6083\,
            DIN => \N__6082\,
            DOUT => \N__6081\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6083\,
            PADOUT => \N__6082\,
            PADIN => \N__6081\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6074\,
            DIN => \N__6073\,
            DOUT => \N__6072\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6074\,
            PADOUT => \N__6073\,
            PADIN => \N__6072\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6065\,
            DIN => \N__6064\,
            DOUT => \N__6063\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6065\,
            PADOUT => \N__6064\,
            PADIN => \N__6063\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6056\,
            DIN => \N__6055\,
            DOUT => \N__6054\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6056\,
            PADOUT => \N__6055\,
            PADIN => \N__6054\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6047\,
            DIN => \N__6046\,
            DOUT => \N__6045\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6047\,
            PADOUT => \N__6046\,
            PADIN => \N__6045\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6038\,
            DIN => \N__6037\,
            DOUT => \N__6036\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6038\,
            PADOUT => \N__6037\,
            PADIN => \N__6036\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nREGSPACE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6029\,
            DIN => \N__6028\,
            DOUT => \N__6027\,
            PACKAGEPIN => \nREGSPACE_wire\
        );

    \nREGSPACE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6029\,
            PADOUT => \N__6028\,
            PADIN => \N__6027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3148\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6020\,
            DIN => \N__6019\,
            DOUT => \N__6018\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6020\,
            PADOUT => \N__6019\,
            PADIN => \N__6018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3448\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6011\,
            DIN => \N__6010\,
            DOUT => \N__6009\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6011\,
            PADOUT => \N__6010\,
            PADIN => \N__6009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6002\,
            DIN => \N__6001\,
            DOUT => \N__6000\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6002\,
            PADOUT => \N__6001\,
            PADIN => \N__6000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5993\,
            DIN => \N__5992\,
            DOUT => \N__5991\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5993\,
            PADOUT => \N__5992\,
            PADIN => \N__5991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5984\,
            DIN => \N__5983\,
            DOUT => \N__5982\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5984\,
            PADOUT => \N__5983\,
            PADIN => \N__5982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5975\,
            DIN => \N__5974\,
            DOUT => \N__5973\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5975\,
            PADOUT => \N__5974\,
            PADIN => \N__5973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5966\,
            DIN => \N__5965\,
            DOUT => \N__5964\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5966\,
            PADOUT => \N__5965\,
            PADIN => \N__5964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4576\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5957\,
            DIN => \N__5956\,
            DOUT => \N__5955\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5957\,
            PADOUT => \N__5956\,
            PADIN => \N__5955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1376\ : InMux
    port map (
            O => \N__5938\,
            I => \N__5929\
        );

    \I__1375\ : InMux
    port map (
            O => \N__5937\,
            I => \N__5929\
        );

    \I__1374\ : InMux
    port map (
            O => \N__5936\,
            I => \N__5929\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__5929\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1372\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5917\
        );

    \I__1371\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5917\
        );

    \I__1370\ : InMux
    port map (
            O => \N__5924\,
            I => \N__5917\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__5917\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1368\ : InMux
    port map (
            O => \N__5914\,
            I => \N__5910\
        );

    \I__1367\ : InMux
    port map (
            O => \N__5913\,
            I => \N__5907\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__5910\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__5907\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\
        );

    \I__1364\ : CEMux
    port map (
            O => \N__5902\,
            I => \N__5899\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__5899\,
            I => \N__5896\
        );

    \I__1362\ : Span4Mux_h
    port map (
            O => \N__5896\,
            I => \N__5893\
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__5893\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\
        );

    \I__1360\ : InMux
    port map (
            O => \N__5890\,
            I => \N__5887\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__5887\,
            I => \N__5884\
        );

    \I__1358\ : Span4Mux_v
    port map (
            O => \N__5884\,
            I => \N__5881\
        );

    \I__1357\ : Odrv4
    port map (
            O => \N__5881\,
            I => \TACK_EN_i\
        );

    \I__1356\ : IoInMux
    port map (
            O => \N__5878\,
            I => \N__5875\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__5875\,
            I => \N__5872\
        );

    \I__1354\ : Span4Mux_s0_v
    port map (
            O => \N__5872\,
            I => \N__5869\
        );

    \I__1353\ : Sp12to4
    port map (
            O => \N__5869\,
            I => \N__5866\
        );

    \I__1352\ : Span12Mux_h
    port map (
            O => \N__5866\,
            I => \N__5863\
        );

    \I__1351\ : Odrv12
    port map (
            O => \N__5863\,
            I => \N_373_i\
        );

    \I__1350\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5853\
        );

    \I__1349\ : InMux
    port map (
            O => \N__5859\,
            I => \N__5848\
        );

    \I__1348\ : InMux
    port map (
            O => \N__5858\,
            I => \N__5848\
        );

    \I__1347\ : InMux
    port map (
            O => \N__5857\,
            I => \N__5845\
        );

    \I__1346\ : InMux
    port map (
            O => \N__5856\,
            I => \N__5842\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__5853\,
            I => \N__5835\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__5848\,
            I => \N__5832\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__5845\,
            I => \N__5829\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__5842\,
            I => \N__5826\
        );

    \I__1341\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5821\
        );

    \I__1340\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5821\
        );

    \I__1339\ : CascadeMux
    port map (
            O => \N__5839\,
            I => \N__5818\
        );

    \I__1338\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5814\
        );

    \I__1337\ : Span4Mux_v
    port map (
            O => \N__5835\,
            I => \N__5811\
        );

    \I__1336\ : Span4Mux_v
    port map (
            O => \N__5832\,
            I => \N__5808\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__5829\,
            I => \N__5805\
        );

    \I__1334\ : Span4Mux_v
    port map (
            O => \N__5826\,
            I => \N__5799\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__5821\,
            I => \N__5799\
        );

    \I__1332\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5794\
        );

    \I__1331\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5794\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__5814\,
            I => \N__5789\
        );

    \I__1329\ : Sp12to4
    port map (
            O => \N__5811\,
            I => \N__5785\
        );

    \I__1328\ : Span4Mux_h
    port map (
            O => \N__5808\,
            I => \N__5782\
        );

    \I__1327\ : Sp12to4
    port map (
            O => \N__5805\,
            I => \N__5779\
        );

    \I__1326\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5776\
        );

    \I__1325\ : Span4Mux_h
    port map (
            O => \N__5799\,
            I => \N__5771\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__5794\,
            I => \N__5771\
        );

    \I__1323\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5766\
        );

    \I__1322\ : InMux
    port map (
            O => \N__5792\,
            I => \N__5766\
        );

    \I__1321\ : Span4Mux_v
    port map (
            O => \N__5789\,
            I => \N__5763\
        );

    \I__1320\ : InMux
    port map (
            O => \N__5788\,
            I => \N__5760\
        );

    \I__1319\ : Span12Mux_h
    port map (
            O => \N__5785\,
            I => \N__5757\
        );

    \I__1318\ : Sp12to4
    port map (
            O => \N__5782\,
            I => \N__5754\
        );

    \I__1317\ : Span12Mux_h
    port map (
            O => \N__5779\,
            I => \N__5745\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__5776\,
            I => \N__5745\
        );

    \I__1315\ : Sp12to4
    port map (
            O => \N__5771\,
            I => \N__5745\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__5766\,
            I => \N__5745\
        );

    \I__1313\ : Sp12to4
    port map (
            O => \N__5763\,
            I => \N__5740\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__5760\,
            I => \N__5740\
        );

    \I__1311\ : Span12Mux_v
    port map (
            O => \N__5757\,
            I => \N__5737\
        );

    \I__1310\ : Span12Mux_h
    port map (
            O => \N__5754\,
            I => \N__5734\
        );

    \I__1309\ : Span12Mux_v
    port map (
            O => \N__5745\,
            I => \N__5731\
        );

    \I__1308\ : Span12Mux_h
    port map (
            O => \N__5740\,
            I => \N__5728\
        );

    \I__1307\ : Span12Mux_h
    port map (
            O => \N__5737\,
            I => \N__5723\
        );

    \I__1306\ : Span12Mux_v
    port map (
            O => \N__5734\,
            I => \N__5723\
        );

    \I__1305\ : Span12Mux_h
    port map (
            O => \N__5731\,
            I => \N__5718\
        );

    \I__1304\ : Span12Mux_v
    port map (
            O => \N__5728\,
            I => \N__5718\
        );

    \I__1303\ : Odrv12
    port map (
            O => \N__5723\,
            I => \RESETn_c\
        );

    \I__1302\ : Odrv12
    port map (
            O => \N__5718\,
            I => \RESETn_c\
        );

    \I__1301\ : IoInMux
    port map (
            O => \N__5713\,
            I => \N__5710\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__5710\,
            I => \N__5707\
        );

    \I__1299\ : Span12Mux_s10_v
    port map (
            O => \N__5707\,
            I => \N__5703\
        );

    \I__1298\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5700\
        );

    \I__1297\ : Span12Mux_h
    port map (
            O => \N__5703\,
            I => \N__5697\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__5700\,
            I => \N__5694\
        );

    \I__1295\ : Odrv12
    port map (
            O => \N__5697\,
            I => \nBUFEN_c\
        );

    \I__1294\ : Odrv12
    port map (
            O => \N__5694\,
            I => \nBUFEN_c\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5686\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__5686\,
            I => \N__5683\
        );

    \I__1291\ : Span4Mux_h
    port map (
            O => \N__5683\,
            I => \N__5680\
        );

    \I__1290\ : Span4Mux_h
    port map (
            O => \N__5680\,
            I => \N__5677\
        );

    \I__1289\ : Sp12to4
    port map (
            O => \N__5677\,
            I => \N__5674\
        );

    \I__1288\ : Span12Mux_v
    port map (
            O => \N__5674\,
            I => \N__5671\
        );

    \I__1287\ : Odrv12
    port map (
            O => \N__5671\,
            I => \TACKn_in\
        );

    \I__1286\ : SRMux
    port map (
            O => \N__5668\,
            I => \N__5665\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__5665\,
            I => \N__5661\
        );

    \I__1284\ : SRMux
    port map (
            O => \N__5664\,
            I => \N__5658\
        );

    \I__1283\ : Span4Mux_v
    port map (
            O => \N__5661\,
            I => \N__5655\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__5658\,
            I => \N__5652\
        );

    \I__1281\ : Sp12to4
    port map (
            O => \N__5655\,
            I => \N__5647\
        );

    \I__1280\ : Span12Mux_v
    port map (
            O => \N__5652\,
            I => \N__5647\
        );

    \I__1279\ : Odrv12
    port map (
            O => \N__5647\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1278\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5641\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5641\,
            I => \U409_TRANSFER_ACK.ROM_TACK_EN_e_1\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__5638\,
            I => \N__5634\
        );

    \I__1275\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5626\
        );

    \I__1274\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5626\
        );

    \I__1273\ : InMux
    port map (
            O => \N__5633\,
            I => \N__5626\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__5626\,
            I => \N__5623\
        );

    \I__1271\ : Span4Mux_v
    port map (
            O => \N__5623\,
            I => \N__5620\
        );

    \I__1270\ : Span4Mux_v
    port map (
            O => \N__5620\,
            I => \N__5617\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__5617\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5607\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5613\,
            I => \N__5607\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5612\,
            I => \N__5604\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__5607\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5604\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1263\ : InMux
    port map (
            O => \N__5599\,
            I => \N__5589\
        );

    \I__1262\ : InMux
    port map (
            O => \N__5598\,
            I => \N__5589\
        );

    \I__1261\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5589\
        );

    \I__1260\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5586\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__5589\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__5586\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__5581\,
            I => \N__5576\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5570\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5579\,
            I => \N__5570\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5576\,
            I => \N__5565\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5575\,
            I => \N__5565\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__5570\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__5565\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1250\ : SRMux
    port map (
            O => \N__5560\,
            I => \N__5555\
        );

    \I__1249\ : SRMux
    port map (
            O => \N__5559\,
            I => \N__5552\
        );

    \I__1248\ : SRMux
    port map (
            O => \N__5558\,
            I => \N__5549\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__5555\,
            I => \N__5545\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__5552\,
            I => \N__5542\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__5549\,
            I => \N__5539\
        );

    \I__1244\ : SRMux
    port map (
            O => \N__5548\,
            I => \N__5536\
        );

    \I__1243\ : Span4Mux_v
    port map (
            O => \N__5545\,
            I => \N__5533\
        );

    \I__1242\ : Span4Mux_v
    port map (
            O => \N__5542\,
            I => \N__5530\
        );

    \I__1241\ : Span4Mux_h
    port map (
            O => \N__5539\,
            I => \N__5527\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__5536\,
            I => \N__5524\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__5533\,
            I => \RESETn_c_i\
        );

    \I__1238\ : Odrv4
    port map (
            O => \N__5530\,
            I => \RESETn_c_i\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__5527\,
            I => \RESETn_c_i\
        );

    \I__1236\ : Odrv12
    port map (
            O => \N__5524\,
            I => \RESETn_c_i\
        );

    \I__1235\ : IoInMux
    port map (
            O => \N__5515\,
            I => \N__5512\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5512\,
            I => \N__5509\
        );

    \I__1233\ : Span12Mux_s7_v
    port map (
            O => \N__5509\,
            I => \N__5506\
        );

    \I__1232\ : Span12Mux_h
    port map (
            O => \N__5506\,
            I => \N__5502\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5505\,
            I => \N__5499\
        );

    \I__1230\ : Odrv12
    port map (
            O => \N__5502\,
            I => \TACK_OUTn\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__5499\,
            I => \TACK_OUTn\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__5494\,
            I => \N__5491\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5486\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5483\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5480\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5486\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5483\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__5480\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5473\,
            I => \N__5469\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5472\,
            I => \N__5466\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5469\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5466\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__5461\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_\
        );

    \I__1216\ : InMux
    port map (
            O => \N__5458\,
            I => \N__5454\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5457\,
            I => \N__5451\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__5454\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5451\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__5446\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5439\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5436\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__5439\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__5436\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5431\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5428\,
            I => \N__5424\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5427\,
            I => \N__5421\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__5424\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__5421\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5416\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5413\,
            I => \N__5409\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5412\,
            I => \N__5406\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5409\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5406\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__1197\ : InMux
    port map (
            O => \N__5401\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__5398\,
            I => \N__5395\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5391\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5388\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5391\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5388\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5383\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5376\
        );

    \I__1189\ : InMux
    port map (
            O => \N__5379\,
            I => \N__5373\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__5376\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5373\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5368\,
            I => \N__5365\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__5365\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5362\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5355\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5358\,
            I => \N__5352\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5355\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__5352\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5344\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5344\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5341\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5338\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5331\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5334\,
            I => \N__5328\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5331\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__5328\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__1171\ : ClkMux
    port map (
            O => \N__5323\,
            I => \N__5299\
        );

    \I__1170\ : ClkMux
    port map (
            O => \N__5322\,
            I => \N__5299\
        );

    \I__1169\ : ClkMux
    port map (
            O => \N__5321\,
            I => \N__5299\
        );

    \I__1168\ : ClkMux
    port map (
            O => \N__5320\,
            I => \N__5299\
        );

    \I__1167\ : ClkMux
    port map (
            O => \N__5319\,
            I => \N__5299\
        );

    \I__1166\ : ClkMux
    port map (
            O => \N__5318\,
            I => \N__5299\
        );

    \I__1165\ : ClkMux
    port map (
            O => \N__5317\,
            I => \N__5299\
        );

    \I__1164\ : ClkMux
    port map (
            O => \N__5316\,
            I => \N__5299\
        );

    \I__1163\ : GlobalMux
    port map (
            O => \N__5299\,
            I => \N__5296\
        );

    \I__1162\ : gio2CtrlBuf
    port map (
            O => \N__5296\,
            I => \CLK6_c_g\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__5293\,
            I => \N__5290\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5290\,
            I => \N__5286\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5289\,
            I => \N__5283\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5286\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5283\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5278\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5272\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5272\,
            I => \N__5268\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5271\,
            I => \N__5265\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__5268\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5265\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5260\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5253\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5256\,
            I => \N__5250\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__5253\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5250\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5245\,
            I => \N__5242\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__5242\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5239\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5232\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5235\,
            I => \N__5229\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5232\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5229\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__1138\ : InMux
    port map (
            O => \N__5224\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5221\,
            I => \N__5217\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5214\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5217\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__5214\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5206\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__5206\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5203\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5200\,
            I => \N__5196\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5199\,
            I => \N__5193\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5196\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5193\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1126\ : InMux
    port map (
            O => \N__5188\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5185\,
            I => \N__5181\
        );

    \I__1124\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5178\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__5181\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__5178\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__5173\,
            I => \N__5170\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5167\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__5167\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5164\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__5161\,
            I => \N__5158\
        );

    \I__1116\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5154\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5151\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__5154\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__5151\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__5146\,
            I => \N__5143\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5143\,
            I => \N__5140\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__5140\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5137\,
            I => \bfn_12_7_0_\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5127\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5120\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5120\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5131\,
            I => \N__5120\
        );

    \I__1104\ : InMux
    port map (
            O => \N__5130\,
            I => \N__5117\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5127\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5120\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5117\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1100\ : IoInMux
    port map (
            O => \N__5110\,
            I => \N__5107\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5107\,
            I => \N__5104\
        );

    \I__1098\ : IoSpan4Mux
    port map (
            O => \N__5104\,
            I => \N__5097\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5094\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5091\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__5101\,
            I => \N__5088\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5085\
        );

    \I__1093\ : Span4Mux_s0_v
    port map (
            O => \N__5097\,
            I => \N__5082\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__5094\,
            I => \N__5077\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5091\,
            I => \N__5077\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5074\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5085\,
            I => \N__5071\
        );

    \I__1088\ : Sp12to4
    port map (
            O => \N__5082\,
            I => \N__5068\
        );

    \I__1087\ : Span4Mux_h
    port map (
            O => \N__5077\,
            I => \N__5063\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5074\,
            I => \N__5063\
        );

    \I__1085\ : Span4Mux_h
    port map (
            O => \N__5071\,
            I => \N__5060\
        );

    \I__1084\ : Span12Mux_v
    port map (
            O => \N__5068\,
            I => \N__5055\
        );

    \I__1083\ : Sp12to4
    port map (
            O => \N__5063\,
            I => \N__5055\
        );

    \I__1082\ : Sp12to4
    port map (
            O => \N__5060\,
            I => \N__5052\
        );

    \I__1081\ : Span12Mux_v
    port map (
            O => \N__5055\,
            I => \N__5049\
        );

    \I__1080\ : Odrv12
    port map (
            O => \N__5052\,
            I => \CLK40_IN_c\
        );

    \I__1079\ : Odrv12
    port map (
            O => \N__5049\,
            I => \CLK40_IN_c\
        );

    \I__1078\ : CascadeMux
    port map (
            O => \N__5044\,
            I => \N__5041\
        );

    \I__1077\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5038\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5038\,
            I => \U409_TRANSFER_ACK.N_107\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__5035\,
            I => \N__5029\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5034\,
            I => \N__5026\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5033\,
            I => \N__5023\
        );

    \I__1072\ : InMux
    port map (
            O => \N__5032\,
            I => \N__5018\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5029\,
            I => \N__5018\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__5026\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5023\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__5018\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__5011\,
            I => \U409_TRANSFER_ACK.N_107_cascade_\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5008\,
            I => \N__5005\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5005\,
            I => \U409_TRANSFER_ACK.m9_bm\
        );

    \I__1064\ : InMux
    port map (
            O => \N__5002\,
            I => \N__4996\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4996\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__4996\,
            I => \U409_TRANSFER_ACK.N_4\
        );

    \I__1061\ : InMux
    port map (
            O => \N__4993\,
            I => \N__4987\
        );

    \I__1060\ : InMux
    port map (
            O => \N__4992\,
            I => \N__4984\
        );

    \I__1059\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4981\
        );

    \I__1058\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4978\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__4987\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__4984\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__4981\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__4978\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__4969\,
            I => \N__4966\
        );

    \I__1052\ : InMux
    port map (
            O => \N__4966\,
            I => \N__4960\
        );

    \I__1051\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4960\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__4960\,
            I => \N__4956\
        );

    \I__1049\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4953\
        );

    \I__1048\ : Odrv4
    port map (
            O => \N__4956\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__4953\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__1046\ : IoInMux
    port map (
            O => \N__4948\,
            I => \N__4945\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__4945\,
            I => \N__4942\
        );

    \I__1044\ : IoSpan4Mux
    port map (
            O => \N__4942\,
            I => \N__4939\
        );

    \I__1043\ : Span4Mux_s1_v
    port map (
            O => \N__4939\,
            I => \N__4936\
        );

    \I__1042\ : Sp12to4
    port map (
            O => \N__4936\,
            I => \N__4932\
        );

    \I__1041\ : InMux
    port map (
            O => \N__4935\,
            I => \N__4929\
        );

    \I__1040\ : Span12Mux_v
    port map (
            O => \N__4932\,
            I => \N__4923\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__4929\,
            I => \N__4923\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4920\
        );

    \I__1037\ : Odrv12
    port map (
            O => \N__4923\,
            I => \CLKCIA_c\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4920\,
            I => \CLKCIA_c\
        );

    \I__1035\ : InMux
    port map (
            O => \N__4915\,
            I => \N__4910\
        );

    \I__1034\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4905\
        );

    \I__1033\ : InMux
    port map (
            O => \N__4913\,
            I => \N__4905\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__4910\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__4905\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1030\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4894\
        );

    \I__1029\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4894\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__4894\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__1027\ : IoInMux
    port map (
            O => \N__4891\,
            I => \N__4888\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__4888\,
            I => \N__4885\
        );

    \I__1025\ : Span4Mux_s2_v
    port map (
            O => \N__4885\,
            I => \N__4882\
        );

    \I__1024\ : Span4Mux_v
    port map (
            O => \N__4882\,
            I => \N__4879\
        );

    \I__1023\ : Odrv4
    port map (
            O => \N__4879\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4876\,
            I => \N__4869\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4875\,
            I => \N__4869\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4874\,
            I => \N__4866\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__4869\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4866\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__4861\,
            I => \N__4855\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4848\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4848\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4848\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4845\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__4848\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4845\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4835\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4832\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4829\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4835\,
            I => \N__4826\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4832\,
            I => \N__4821\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__4829\,
            I => \N__4821\
        );

    \I__1004\ : Span4Mux_v
    port map (
            O => \N__4826\,
            I => \N__4818\
        );

    \I__1003\ : Span12Mux_h
    port map (
            O => \N__4821\,
            I => \N__4815\
        );

    \I__1002\ : Sp12to4
    port map (
            O => \N__4818\,
            I => \N__4812\
        );

    \I__1001\ : Span12Mux_v
    port map (
            O => \N__4815\,
            I => \N__4809\
        );

    \I__1000\ : Span12Mux_h
    port map (
            O => \N__4812\,
            I => \N__4806\
        );

    \I__999\ : Odrv12
    port map (
            O => \N__4809\,
            I => \TSn_c\
        );

    \I__998\ : Odrv12
    port map (
            O => \N__4806\,
            I => \TSn_c\
        );

    \I__997\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4795\
        );

    \I__996\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4790\
        );

    \I__995\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4790\
        );

    \I__994\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4787\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4795\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__4790\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__4787\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__4780\,
            I => \N__4775\
        );

    \I__989\ : CascadeMux
    port map (
            O => \N__4779\,
            I => \N__4769\
        );

    \I__988\ : CascadeMux
    port map (
            O => \N__4778\,
            I => \N__4766\
        );

    \I__987\ : InMux
    port map (
            O => \N__4775\,
            I => \N__4758\
        );

    \I__986\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4758\
        );

    \I__985\ : InMux
    port map (
            O => \N__4773\,
            I => \N__4758\
        );

    \I__984\ : InMux
    port map (
            O => \N__4772\,
            I => \N__4753\
        );

    \I__983\ : InMux
    port map (
            O => \N__4769\,
            I => \N__4753\
        );

    \I__982\ : InMux
    port map (
            O => \N__4766\,
            I => \N__4750\
        );

    \I__981\ : InMux
    port map (
            O => \N__4765\,
            I => \N__4747\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4758\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4753\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__4750\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4747\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__976\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4729\
        );

    \I__975\ : InMux
    port map (
            O => \N__4737\,
            I => \N__4729\
        );

    \I__974\ : InMux
    port map (
            O => \N__4736\,
            I => \N__4724\
        );

    \I__973\ : InMux
    port map (
            O => \N__4735\,
            I => \N__4724\
        );

    \I__972\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4721\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4729\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4724\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4721\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__968\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4711\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4711\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__966\ : InMux
    port map (
            O => \N__4708\,
            I => \N__4701\
        );

    \I__965\ : InMux
    port map (
            O => \N__4707\,
            I => \N__4701\
        );

    \I__964\ : InMux
    port map (
            O => \N__4706\,
            I => \N__4698\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__4701\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__4698\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__961\ : InMux
    port map (
            O => \N__4693\,
            I => \N__4690\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4690\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\
        );

    \I__959\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4681\
        );

    \I__958\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4678\
        );

    \I__957\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4673\
        );

    \I__956\ : InMux
    port map (
            O => \N__4684\,
            I => \N__4673\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4681\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4678\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4673\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__952\ : InMux
    port map (
            O => \N__4666\,
            I => \N__4657\
        );

    \I__951\ : InMux
    port map (
            O => \N__4665\,
            I => \N__4657\
        );

    \I__950\ : InMux
    port map (
            O => \N__4664\,
            I => \N__4654\
        );

    \I__949\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4651\
        );

    \I__948\ : InMux
    port map (
            O => \N__4662\,
            I => \N__4648\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4657\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4654\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4651\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4648\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__4639\,
            I => \N__4636\
        );

    \I__942\ : InMux
    port map (
            O => \N__4636\,
            I => \N__4630\
        );

    \I__941\ : InMux
    port map (
            O => \N__4635\,
            I => \N__4630\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4630\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\
        );

    \I__939\ : InMux
    port map (
            O => \N__4627\,
            I => \N__4620\
        );

    \I__938\ : InMux
    port map (
            O => \N__4626\,
            I => \N__4611\
        );

    \I__937\ : InMux
    port map (
            O => \N__4625\,
            I => \N__4611\
        );

    \I__936\ : InMux
    port map (
            O => \N__4624\,
            I => \N__4611\
        );

    \I__935\ : InMux
    port map (
            O => \N__4623\,
            I => \N__4611\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4620\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4611\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__932\ : CascadeMux
    port map (
            O => \N__4606\,
            I => \N__4600\
        );

    \I__931\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4597\
        );

    \I__930\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4594\
        );

    \I__929\ : InMux
    port map (
            O => \N__4603\,
            I => \N__4589\
        );

    \I__928\ : InMux
    port map (
            O => \N__4600\,
            I => \N__4589\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4597\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4594\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4589\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__4582\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__923\ : CascadeMux
    port map (
            O => \N__4579\,
            I => \U409_TICK.TICK603_10_cascade_\
        );

    \I__922\ : IoInMux
    port map (
            O => \N__4576\,
            I => \N__4573\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4573\,
            I => \N__4570\
        );

    \I__920\ : Span4Mux_s0_v
    port map (
            O => \N__4570\,
            I => \N__4567\
        );

    \I__919\ : Sp12to4
    port map (
            O => \N__4567\,
            I => \N__4564\
        );

    \I__918\ : Span12Mux_h
    port map (
            O => \N__4564\,
            I => \N__4561\
        );

    \I__917\ : Span12Mux_v
    port map (
            O => \N__4561\,
            I => \N__4557\
        );

    \I__916\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4554\
        );

    \I__915\ : Odrv12
    port map (
            O => \N__4557\,
            I => \TICK60_c\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4554\,
            I => \TICK60_c\
        );

    \I__913\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4536\
        );

    \I__912\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4536\
        );

    \I__911\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4536\
        );

    \I__910\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4527\
        );

    \I__909\ : InMux
    port map (
            O => \N__4545\,
            I => \N__4527\
        );

    \I__908\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4527\
        );

    \I__907\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4527\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4536\,
            I => \U409_TICK.TICK603_10\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4527\,
            I => \U409_TICK.TICK603_10\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__4522\,
            I => \N__4518\
        );

    \I__903\ : InMux
    port map (
            O => \N__4521\,
            I => \N__4510\
        );

    \I__902\ : InMux
    port map (
            O => \N__4518\,
            I => \N__4507\
        );

    \I__901\ : InMux
    port map (
            O => \N__4517\,
            I => \N__4496\
        );

    \I__900\ : InMux
    port map (
            O => \N__4516\,
            I => \N__4496\
        );

    \I__899\ : InMux
    port map (
            O => \N__4515\,
            I => \N__4496\
        );

    \I__898\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4496\
        );

    \I__897\ : InMux
    port map (
            O => \N__4513\,
            I => \N__4496\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4510\,
            I => \U409_TICK.TICK603_14\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4507\,
            I => \U409_TICK.TICK603_14\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4496\,
            I => \U409_TICK.TICK603_14\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__4489\,
            I => \N__4480\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__4488\,
            I => \N__4477\
        );

    \I__891\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4472\
        );

    \I__890\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4472\
        );

    \I__889\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4461\
        );

    \I__888\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4461\
        );

    \I__887\ : InMux
    port map (
            O => \N__4483\,
            I => \N__4461\
        );

    \I__886\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4461\
        );

    \I__885\ : InMux
    port map (
            O => \N__4477\,
            I => \N__4461\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4472\,
            I => \U409_TICK.TICK603_9\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__4461\,
            I => \U409_TICK.TICK603_9\
        );

    \I__882\ : CascadeMux
    port map (
            O => \N__4456\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__4453\,
            I => \N__4450\
        );

    \I__880\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4444\
        );

    \I__879\ : InMux
    port map (
            O => \N__4449\,
            I => \N__4444\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4444\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__877\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4438\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4438\,
            I => \N__4434\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__4437\,
            I => \N__4431\
        );

    \I__874\ : Span4Mux_v
    port map (
            O => \N__4434\,
            I => \N__4428\
        );

    \I__873\ : InMux
    port map (
            O => \N__4431\,
            I => \N__4425\
        );

    \I__872\ : Odrv4
    port map (
            O => \N__4428\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4425\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\
        );

    \I__870\ : InMux
    port map (
            O => \N__4420\,
            I => \N__4416\
        );

    \I__869\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4413\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4416\,
            I => \N__4410\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4413\,
            I => \N__4407\
        );

    \I__866\ : Odrv4
    port map (
            O => \N__4410\,
            I => \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__4407\,
            I => \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0\
        );

    \I__864\ : CascadeMux
    port map (
            O => \N__4402\,
            I => \N__4399\
        );

    \I__863\ : InMux
    port map (
            O => \N__4399\,
            I => \N__4396\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4396\,
            I => \N__4391\
        );

    \I__861\ : InMux
    port map (
            O => \N__4395\,
            I => \N__4387\
        );

    \I__860\ : InMux
    port map (
            O => \N__4394\,
            I => \N__4382\
        );

    \I__859\ : Span4Mux_v
    port map (
            O => \N__4391\,
            I => \N__4379\
        );

    \I__858\ : InMux
    port map (
            O => \N__4390\,
            I => \N__4376\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4387\,
            I => \N__4373\
        );

    \I__856\ : InMux
    port map (
            O => \N__4386\,
            I => \N__4368\
        );

    \I__855\ : InMux
    port map (
            O => \N__4385\,
            I => \N__4368\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4382\,
            I => \N__4364\
        );

    \I__853\ : Sp12to4
    port map (
            O => \N__4379\,
            I => \N__4359\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__4376\,
            I => \N__4359\
        );

    \I__851\ : Span4Mux_v
    port map (
            O => \N__4373\,
            I => \N__4356\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4368\,
            I => \N__4353\
        );

    \I__849\ : InMux
    port map (
            O => \N__4367\,
            I => \N__4350\
        );

    \I__848\ : Span12Mux_v
    port map (
            O => \N__4364\,
            I => \N__4347\
        );

    \I__847\ : Span12Mux_h
    port map (
            O => \N__4359\,
            I => \N__4344\
        );

    \I__846\ : Span4Mux_h
    port map (
            O => \N__4356\,
            I => \N__4341\
        );

    \I__845\ : Span4Mux_h
    port map (
            O => \N__4353\,
            I => \N__4338\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4350\,
            I => \N__4335\
        );

    \I__843\ : Odrv12
    port map (
            O => \N__4347\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0\
        );

    \I__842\ : Odrv12
    port map (
            O => \N__4344\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0\
        );

    \I__841\ : Odrv4
    port map (
            O => \N__4341\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__4338\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0\
        );

    \I__839\ : Odrv4
    port map (
            O => \N__4335\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0\
        );

    \I__838\ : InMux
    port map (
            O => \N__4324\,
            I => \N__4321\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4321\,
            I => \N__4318\
        );

    \I__836\ : Span4Mux_v
    port map (
            O => \N__4318\,
            I => \N__4313\
        );

    \I__835\ : InMux
    port map (
            O => \N__4317\,
            I => \N__4310\
        );

    \I__834\ : InMux
    port map (
            O => \N__4316\,
            I => \N__4307\
        );

    \I__833\ : Sp12to4
    port map (
            O => \N__4313\,
            I => \N__4300\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4310\,
            I => \N__4300\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4307\,
            I => \N__4300\
        );

    \I__830\ : Span12Mux_h
    port map (
            O => \N__4300\,
            I => \N__4297\
        );

    \I__829\ : Span12Mux_v
    port map (
            O => \N__4297\,
            I => \N__4294\
        );

    \I__828\ : Odrv12
    port map (
            O => \N__4294\,
            I => \OVL_c\
        );

    \I__827\ : InMux
    port map (
            O => \N__4291\,
            I => \N__4286\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__4290\,
            I => \N__4282\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__4289\,
            I => \N__4279\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4286\,
            I => \N__4276\
        );

    \I__823\ : InMux
    port map (
            O => \N__4285\,
            I => \N__4273\
        );

    \I__822\ : InMux
    port map (
            O => \N__4282\,
            I => \N__4268\
        );

    \I__821\ : InMux
    port map (
            O => \N__4279\,
            I => \N__4268\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__4276\,
            I => \U409_CIA.VMAZ0\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4273\,
            I => \U409_CIA.VMAZ0\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4268\,
            I => \U409_CIA.VMAZ0\
        );

    \I__817\ : InMux
    port map (
            O => \N__4261\,
            I => \N__4258\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4258\,
            I => \N__4253\
        );

    \I__815\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4248\
        );

    \I__814\ : InMux
    port map (
            O => \N__4256\,
            I => \N__4248\
        );

    \I__813\ : Sp12to4
    port map (
            O => \N__4253\,
            I => \N__4243\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__4248\,
            I => \N__4243\
        );

    \I__811\ : Odrv12
    port map (
            O => \N__4243\,
            I => \U409_CIA.g0Z0Z_14\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__4240\,
            I => \N__4237\
        );

    \I__809\ : InMux
    port map (
            O => \N__4237\,
            I => \N__4232\
        );

    \I__808\ : InMux
    port map (
            O => \N__4236\,
            I => \N__4227\
        );

    \I__807\ : InMux
    port map (
            O => \N__4235\,
            I => \N__4227\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4232\,
            I => \N__4222\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__4227\,
            I => \N__4222\
        );

    \I__804\ : Span4Mux_h
    port map (
            O => \N__4222\,
            I => \N__4219\
        );

    \I__803\ : Span4Mux_v
    port map (
            O => \N__4219\,
            I => \N__4216\
        );

    \I__802\ : Span4Mux_h
    port map (
            O => \N__4216\,
            I => \N__4213\
        );

    \I__801\ : Odrv4
    port map (
            O => \N__4213\,
            I => \U409_CIA.g0Z0Z_13\
        );

    \I__800\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4205\
        );

    \I__799\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4200\
        );

    \I__798\ : InMux
    port map (
            O => \N__4208\,
            I => \N__4200\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4205\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4200\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__4195\,
            I => \U409_TICK.TICK603_8_cascade_\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__4192\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__793\ : InMux
    port map (
            O => \N__4189\,
            I => \N__4186\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4186\,
            I => \U409_TICK.TICK603_11\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__4183\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\
        );

    \I__790\ : InMux
    port map (
            O => \N__4180\,
            I => \N__4173\
        );

    \I__789\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4173\
        );

    \I__788\ : InMux
    port map (
            O => \N__4178\,
            I => \N__4170\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4173\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4170\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__4165\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\
        );

    \I__784\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4156\
        );

    \I__783\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4156\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__4156\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__781\ : CascadeMux
    port map (
            O => \N__4153\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__4150\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__779\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4139\
        );

    \I__778\ : InMux
    port map (
            O => \N__4146\,
            I => \N__4139\
        );

    \I__777\ : InMux
    port map (
            O => \N__4145\,
            I => \N__4134\
        );

    \I__776\ : InMux
    port map (
            O => \N__4144\,
            I => \N__4134\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4139\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4134\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__773\ : CascadeMux
    port map (
            O => \N__4129\,
            I => \U409_TRANSFER_ACK.m9_am_cascade_\
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__4126\,
            I => \U409_TRANSFER_ACK.i6_mux_0_cascade_\
        );

    \I__771\ : InMux
    port map (
            O => \N__4123\,
            I => \N__4120\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4120\,
            I => \N__4116\
        );

    \I__769\ : InMux
    port map (
            O => \N__4119\,
            I => \N__4113\
        );

    \I__768\ : Span12Mux_h
    port map (
            O => \N__4116\,
            I => \N__4108\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4113\,
            I => \N__4108\
        );

    \I__766\ : Odrv12
    port map (
            O => \N__4108\,
            I => \CIA_ENABLEm\
        );

    \I__765\ : InMux
    port map (
            O => \N__4105\,
            I => \N__4099\
        );

    \I__764\ : InMux
    port map (
            O => \N__4104\,
            I => \N__4096\
        );

    \I__763\ : InMux
    port map (
            O => \N__4103\,
            I => \N__4089\
        );

    \I__762\ : InMux
    port map (
            O => \N__4102\,
            I => \N__4089\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4099\,
            I => \N__4086\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4096\,
            I => \N__4083\
        );

    \I__759\ : InMux
    port map (
            O => \N__4095\,
            I => \N__4078\
        );

    \I__758\ : InMux
    port map (
            O => \N__4094\,
            I => \N__4078\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__4089\,
            I => \N__4075\
        );

    \I__756\ : Span4Mux_v
    port map (
            O => \N__4086\,
            I => \N__4068\
        );

    \I__755\ : Span4Mux_h
    port map (
            O => \N__4083\,
            I => \N__4068\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__4078\,
            I => \N__4068\
        );

    \I__753\ : Sp12to4
    port map (
            O => \N__4075\,
            I => \N__4064\
        );

    \I__752\ : Span4Mux_v
    port map (
            O => \N__4068\,
            I => \N__4061\
        );

    \I__751\ : InMux
    port map (
            O => \N__4067\,
            I => \N__4058\
        );

    \I__750\ : Span12Mux_v
    port map (
            O => \N__4064\,
            I => \N__4055\
        );

    \I__749\ : Span4Mux_v
    port map (
            O => \N__4061\,
            I => \N__4052\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4058\,
            I => \N__4049\
        );

    \I__747\ : Span12Mux_h
    port map (
            O => \N__4055\,
            I => \N__4046\
        );

    \I__746\ : Sp12to4
    port map (
            O => \N__4052\,
            I => \N__4041\
        );

    \I__745\ : Span12Mux_v
    port map (
            O => \N__4049\,
            I => \N__4041\
        );

    \I__744\ : Odrv12
    port map (
            O => \N__4046\,
            I => \A_c_22\
        );

    \I__743\ : Odrv12
    port map (
            O => \N__4041\,
            I => \A_c_22\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__4036\,
            I => \N__4033\
        );

    \I__741\ : InMux
    port map (
            O => \N__4033\,
            I => \N__4023\
        );

    \I__740\ : InMux
    port map (
            O => \N__4032\,
            I => \N__4023\
        );

    \I__739\ : InMux
    port map (
            O => \N__4031\,
            I => \N__4019\
        );

    \I__738\ : InMux
    port map (
            O => \N__4030\,
            I => \N__4014\
        );

    \I__737\ : InMux
    port map (
            O => \N__4029\,
            I => \N__4014\
        );

    \I__736\ : InMux
    port map (
            O => \N__4028\,
            I => \N__4011\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__4023\,
            I => \N__4008\
        );

    \I__734\ : InMux
    port map (
            O => \N__4022\,
            I => \N__4005\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4019\,
            I => \N__4002\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4014\,
            I => \N__3998\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4011\,
            I => \N__3995\
        );

    \I__730\ : Span4Mux_v
    port map (
            O => \N__4008\,
            I => \N__3992\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__4005\,
            I => \N__3989\
        );

    \I__728\ : Span4Mux_v
    port map (
            O => \N__4002\,
            I => \N__3986\
        );

    \I__727\ : InMux
    port map (
            O => \N__4001\,
            I => \N__3983\
        );

    \I__726\ : Sp12to4
    port map (
            O => \N__3998\,
            I => \N__3980\
        );

    \I__725\ : Span4Mux_v
    port map (
            O => \N__3995\,
            I => \N__3977\
        );

    \I__724\ : Sp12to4
    port map (
            O => \N__3992\,
            I => \N__3968\
        );

    \I__723\ : Span12Mux_v
    port map (
            O => \N__3989\,
            I => \N__3968\
        );

    \I__722\ : Sp12to4
    port map (
            O => \N__3986\,
            I => \N__3968\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__3983\,
            I => \N__3968\
        );

    \I__720\ : Span12Mux_v
    port map (
            O => \N__3980\,
            I => \N__3965\
        );

    \I__719\ : Span4Mux_h
    port map (
            O => \N__3977\,
            I => \N__3962\
        );

    \I__718\ : Odrv12
    port map (
            O => \N__3968\,
            I => \A_c_23\
        );

    \I__717\ : Odrv12
    port map (
            O => \N__3965\,
            I => \A_c_23\
        );

    \I__716\ : Odrv4
    port map (
            O => \N__3962\,
            I => \A_c_23\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__3955\,
            I => \N__3951\
        );

    \I__714\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3946\
        );

    \I__713\ : InMux
    port map (
            O => \N__3951\,
            I => \N__3946\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__3946\,
            I => \N__3940\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__3945\,
            I => \N__3937\
        );

    \I__710\ : InMux
    port map (
            O => \N__3944\,
            I => \N__3932\
        );

    \I__709\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3932\
        );

    \I__708\ : Span4Mux_v
    port map (
            O => \N__3940\,
            I => \N__3929\
        );

    \I__707\ : InMux
    port map (
            O => \N__3937\,
            I => \N__3926\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3932\,
            I => \N__3923\
        );

    \I__705\ : Span4Mux_h
    port map (
            O => \N__3929\,
            I => \N__3920\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__3926\,
            I => \N__3917\
        );

    \I__703\ : Span4Mux_v
    port map (
            O => \N__3923\,
            I => \N__3914\
        );

    \I__702\ : Span4Mux_h
    port map (
            O => \N__3920\,
            I => \N__3909\
        );

    \I__701\ : Span4Mux_v
    port map (
            O => \N__3917\,
            I => \N__3909\
        );

    \I__700\ : Span4Mux_h
    port map (
            O => \N__3914\,
            I => \N__3906\
        );

    \I__699\ : Span4Mux_h
    port map (
            O => \N__3909\,
            I => \N__3903\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__3906\,
            I => \A_c_21\
        );

    \I__697\ : Odrv4
    port map (
            O => \N__3903\,
            I => \A_c_21\
        );

    \I__696\ : InMux
    port map (
            O => \N__3898\,
            I => \N__3895\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__3895\,
            I => \N__3892\
        );

    \I__694\ : Span4Mux_h
    port map (
            O => \N__3892\,
            I => \N__3889\
        );

    \I__693\ : Span4Mux_h
    port map (
            O => \N__3889\,
            I => \N__3886\
        );

    \I__692\ : Odrv4
    port map (
            O => \N__3886\,
            I => \AUTOVECTORm\
        );

    \I__691\ : IoInMux
    port map (
            O => \N__3883\,
            I => \N__3880\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3880\,
            I => \N__3877\
        );

    \I__689\ : IoSpan4Mux
    port map (
            O => \N__3877\,
            I => \N__3874\
        );

    \I__688\ : Span4Mux_s2_v
    port map (
            O => \N__3874\,
            I => \N__3871\
        );

    \I__687\ : Span4Mux_v
    port map (
            O => \N__3871\,
            I => \N__3868\
        );

    \I__686\ : Span4Mux_v
    port map (
            O => \N__3868\,
            I => \N__3865\
        );

    \I__685\ : Odrv4
    port map (
            O => \N__3865\,
            I => \ROMENm_i\
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__3862\,
            I => \N__3858\
        );

    \I__683\ : InMux
    port map (
            O => \N__3861\,
            I => \N__3853\
        );

    \I__682\ : InMux
    port map (
            O => \N__3858\,
            I => \N__3853\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3853\,
            I => \N__3850\
        );

    \I__680\ : Odrv4
    port map (
            O => \N__3850\,
            I => \U409_ADDRESS_DECODE.LOWROMZ0\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__3847\,
            I => \N__3844\
        );

    \I__678\ : InMux
    port map (
            O => \N__3844\,
            I => \N__3838\
        );

    \I__677\ : InMux
    port map (
            O => \N__3843\,
            I => \N__3838\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3838\,
            I => \N__3835\
        );

    \I__675\ : Span4Mux_h
    port map (
            O => \N__3835\,
            I => \N__3832\
        );

    \I__674\ : Odrv4
    port map (
            O => \N__3832\,
            I => \U409_ADDRESS_DECODE.HIROMZ0\
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__3829\,
            I => \N__3826\
        );

    \I__672\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3823\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3823\,
            I => \ROMENm\
        );

    \I__670\ : InMux
    port map (
            O => \N__3820\,
            I => \N__3816\
        );

    \I__669\ : InMux
    port map (
            O => \N__3819\,
            I => \N__3813\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3816\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3813\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__666\ : InMux
    port map (
            O => \N__3808\,
            I => \N__3804\
        );

    \I__665\ : InMux
    port map (
            O => \N__3807\,
            I => \N__3801\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__3804\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__3801\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__3796\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__661\ : InMux
    port map (
            O => \N__3793\,
            I => \N__3790\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3790\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__659\ : InMux
    port map (
            O => \N__3787\,
            I => \N__3783\
        );

    \I__658\ : InMux
    port map (
            O => \N__3786\,
            I => \N__3780\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3783\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3780\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__655\ : InMux
    port map (
            O => \N__3775\,
            I => \N__3772\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3772\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__653\ : InMux
    port map (
            O => \N__3769\,
            I => \N__3765\
        );

    \I__652\ : InMux
    port map (
            O => \N__3768\,
            I => \N__3762\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3765\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__3762\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__649\ : CascadeMux
    port map (
            O => \N__3757\,
            I => \N__3754\
        );

    \I__648\ : InMux
    port map (
            O => \N__3754\,
            I => \N__3750\
        );

    \I__647\ : InMux
    port map (
            O => \N__3753\,
            I => \N__3747\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3750\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3747\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__644\ : InMux
    port map (
            O => \N__3742\,
            I => \N__3738\
        );

    \I__643\ : InMux
    port map (
            O => \N__3741\,
            I => \N__3735\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3738\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3735\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__640\ : InMux
    port map (
            O => \N__3730\,
            I => \N__3727\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__3727\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__638\ : CascadeMux
    port map (
            O => \N__3724\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__637\ : CascadeMux
    port map (
            O => \N__3721\,
            I => \N__3718\
        );

    \I__636\ : InMux
    port map (
            O => \N__3718\,
            I => \N__3714\
        );

    \I__635\ : InMux
    port map (
            O => \N__3717\,
            I => \N__3711\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3714\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3711\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__632\ : InMux
    port map (
            O => \N__3706\,
            I => \N__3690\
        );

    \I__631\ : InMux
    port map (
            O => \N__3705\,
            I => \N__3690\
        );

    \I__630\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3690\
        );

    \I__629\ : InMux
    port map (
            O => \N__3703\,
            I => \N__3690\
        );

    \I__628\ : InMux
    port map (
            O => \N__3702\,
            I => \N__3681\
        );

    \I__627\ : InMux
    port map (
            O => \N__3701\,
            I => \N__3681\
        );

    \I__626\ : InMux
    port map (
            O => \N__3700\,
            I => \N__3681\
        );

    \I__625\ : InMux
    port map (
            O => \N__3699\,
            I => \N__3681\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3690\,
            I => \U409_TICK.TICK503_10\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3681\,
            I => \U409_TICK.TICK503_10\
        );

    \I__622\ : CascadeMux
    port map (
            O => \N__3676\,
            I => \N__3668\
        );

    \I__621\ : InMux
    port map (
            O => \N__3675\,
            I => \N__3655\
        );

    \I__620\ : InMux
    port map (
            O => \N__3674\,
            I => \N__3655\
        );

    \I__619\ : InMux
    port map (
            O => \N__3673\,
            I => \N__3655\
        );

    \I__618\ : InMux
    port map (
            O => \N__3672\,
            I => \N__3655\
        );

    \I__617\ : InMux
    port map (
            O => \N__3671\,
            I => \N__3655\
        );

    \I__616\ : InMux
    port map (
            O => \N__3668\,
            I => \N__3652\
        );

    \I__615\ : InMux
    port map (
            O => \N__3667\,
            I => \N__3647\
        );

    \I__614\ : InMux
    port map (
            O => \N__3666\,
            I => \N__3647\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3655\,
            I => \N__3644\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3652\,
            I => \U409_TICK.TICK503_14\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3647\,
            I => \U409_TICK.TICK503_14\
        );

    \I__610\ : Odrv4
    port map (
            O => \N__3644\,
            I => \U409_TICK.TICK503_14\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__3637\,
            I => \N__3628\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__3636\,
            I => \N__3625\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__3635\,
            I => \N__3621\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__3634\,
            I => \N__3618\
        );

    \I__605\ : InMux
    port map (
            O => \N__3633\,
            I => \N__3609\
        );

    \I__604\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3609\
        );

    \I__603\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3609\
        );

    \I__602\ : InMux
    port map (
            O => \N__3628\,
            I => \N__3609\
        );

    \I__601\ : InMux
    port map (
            O => \N__3625\,
            I => \N__3606\
        );

    \I__600\ : InMux
    port map (
            O => \N__3624\,
            I => \N__3599\
        );

    \I__599\ : InMux
    port map (
            O => \N__3621\,
            I => \N__3599\
        );

    \I__598\ : InMux
    port map (
            O => \N__3618\,
            I => \N__3599\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3609\,
            I => \U409_TICK.TICK503_9\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3606\,
            I => \U409_TICK.TICK503_9\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3599\,
            I => \U409_TICK.TICK503_9\
        );

    \I__594\ : InMux
    port map (
            O => \N__3592\,
            I => \N__3589\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3589\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__592\ : InMux
    port map (
            O => \N__3586\,
            I => \N__3582\
        );

    \I__591\ : InMux
    port map (
            O => \N__3585\,
            I => \N__3579\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3582\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3579\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__588\ : IoInMux
    port map (
            O => \N__3574\,
            I => \N__3571\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3571\,
            I => \N__3568\
        );

    \I__586\ : IoSpan4Mux
    port map (
            O => \N__3568\,
            I => \N__3565\
        );

    \I__585\ : Span4Mux_s2_v
    port map (
            O => \N__3565\,
            I => \N__3562\
        );

    \I__584\ : Sp12to4
    port map (
            O => \N__3562\,
            I => \N__3559\
        );

    \I__583\ : Span12Mux_s11_v
    port map (
            O => \N__3559\,
            I => \N__3556\
        );

    \I__582\ : Odrv12
    port map (
            O => \N__3556\,
            I => \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\
        );

    \I__581\ : ClkMux
    port map (
            O => \N__3553\,
            I => \N__3541\
        );

    \I__580\ : ClkMux
    port map (
            O => \N__3552\,
            I => \N__3541\
        );

    \I__579\ : ClkMux
    port map (
            O => \N__3551\,
            I => \N__3541\
        );

    \I__578\ : ClkMux
    port map (
            O => \N__3550\,
            I => \N__3541\
        );

    \I__577\ : GlobalMux
    port map (
            O => \N__3541\,
            I => \N__3538\
        );

    \I__576\ : gio2CtrlBuf
    port map (
            O => \N__3538\,
            I => \CLK28_IN_c_g\
        );

    \I__575\ : InMux
    port map (
            O => \N__3535\,
            I => \N__3531\
        );

    \I__574\ : InMux
    port map (
            O => \N__3534\,
            I => \N__3528\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3531\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3528\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__571\ : InMux
    port map (
            O => \N__3523\,
            I => \N__3519\
        );

    \I__570\ : InMux
    port map (
            O => \N__3522\,
            I => \N__3516\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3519\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3516\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__3511\,
            I => \N__3507\
        );

    \I__566\ : InMux
    port map (
            O => \N__3510\,
            I => \N__3504\
        );

    \I__565\ : InMux
    port map (
            O => \N__3507\,
            I => \N__3501\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__3504\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3501\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__562\ : InMux
    port map (
            O => \N__3496\,
            I => \N__3492\
        );

    \I__561\ : InMux
    port map (
            O => \N__3495\,
            I => \N__3489\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3492\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3489\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__558\ : InMux
    port map (
            O => \N__3484\,
            I => \N__3481\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3481\,
            I => \U409_TICK.TICK503_11\
        );

    \I__556\ : InMux
    port map (
            O => \N__3478\,
            I => \N__3474\
        );

    \I__555\ : InMux
    port map (
            O => \N__3477\,
            I => \N__3471\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3474\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3471\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__552\ : CascadeMux
    port map (
            O => \N__3466\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__551\ : InMux
    port map (
            O => \N__3463\,
            I => \N__3459\
        );

    \I__550\ : InMux
    port map (
            O => \N__3462\,
            I => \N__3456\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3459\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3456\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__547\ : CascadeMux
    port map (
            O => \N__3451\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__546\ : IoInMux
    port map (
            O => \N__3448\,
            I => \N__3445\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3445\,
            I => \N__3442\
        );

    \I__544\ : Span4Mux_s1_v
    port map (
            O => \N__3442\,
            I => \N__3439\
        );

    \I__543\ : Sp12to4
    port map (
            O => \N__3439\,
            I => \N__3436\
        );

    \I__542\ : Span12Mux_h
    port map (
            O => \N__3436\,
            I => \N__3433\
        );

    \I__541\ : Span12Mux_v
    port map (
            O => \N__3433\,
            I => \N__3429\
        );

    \I__540\ : InMux
    port map (
            O => \N__3432\,
            I => \N__3426\
        );

    \I__539\ : Odrv12
    port map (
            O => \N__3429\,
            I => \TICK50_c\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3426\,
            I => \TICK50_c\
        );

    \I__537\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3418\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3418\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__3415\,
            I => \N__3411\
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__3414\,
            I => \N__3406\
        );

    \I__533\ : InMux
    port map (
            O => \N__3411\,
            I => \N__3403\
        );

    \I__532\ : InMux
    port map (
            O => \N__3410\,
            I => \N__3398\
        );

    \I__531\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3398\
        );

    \I__530\ : InMux
    port map (
            O => \N__3406\,
            I => \N__3395\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3403\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3398\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3395\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__526\ : InMux
    port map (
            O => \N__3388\,
            I => \N__3381\
        );

    \I__525\ : InMux
    port map (
            O => \N__3387\,
            I => \N__3381\
        );

    \I__524\ : InMux
    port map (
            O => \N__3386\,
            I => \N__3378\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3381\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3378\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__521\ : InMux
    port map (
            O => \N__3373\,
            I => \N__3370\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3370\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__519\ : InMux
    port map (
            O => \N__3367\,
            I => \N__3363\
        );

    \I__518\ : InMux
    port map (
            O => \N__3366\,
            I => \N__3360\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3363\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3360\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__515\ : InMux
    port map (
            O => \N__3355\,
            I => \N__3352\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__3352\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__513\ : InMux
    port map (
            O => \N__3349\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__512\ : InMux
    port map (
            O => \N__3346\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__3343\,
            I => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\
        );

    \I__510\ : InMux
    port map (
            O => \N__3340\,
            I => \N__3332\
        );

    \I__509\ : InMux
    port map (
            O => \N__3339\,
            I => \N__3332\
        );

    \I__508\ : InMux
    port map (
            O => \N__3338\,
            I => \N__3327\
        );

    \I__507\ : InMux
    port map (
            O => \N__3337\,
            I => \N__3327\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3332\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3327\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__504\ : CascadeMux
    port map (
            O => \N__3322\,
            I => \N__3317\
        );

    \I__503\ : InMux
    port map (
            O => \N__3321\,
            I => \N__3311\
        );

    \I__502\ : InMux
    port map (
            O => \N__3320\,
            I => \N__3311\
        );

    \I__501\ : InMux
    port map (
            O => \N__3317\,
            I => \N__3306\
        );

    \I__500\ : InMux
    port map (
            O => \N__3316\,
            I => \N__3306\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3311\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3306\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__3301\,
            I => \N__3297\
        );

    \I__496\ : InMux
    port map (
            O => \N__3300\,
            I => \N__3292\
        );

    \I__495\ : InMux
    port map (
            O => \N__3297\,
            I => \N__3287\
        );

    \I__494\ : InMux
    port map (
            O => \N__3296\,
            I => \N__3287\
        );

    \I__493\ : InMux
    port map (
            O => \N__3295\,
            I => \N__3284\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3292\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3287\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3284\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__489\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3269\
        );

    \I__488\ : InMux
    port map (
            O => \N__3276\,
            I => \N__3262\
        );

    \I__487\ : InMux
    port map (
            O => \N__3275\,
            I => \N__3262\
        );

    \I__486\ : InMux
    port map (
            O => \N__3274\,
            I => \N__3262\
        );

    \I__485\ : InMux
    port map (
            O => \N__3273\,
            I => \N__3257\
        );

    \I__484\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3257\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__3269\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3262\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3257\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__480\ : InMux
    port map (
            O => \N__3250\,
            I => \N__3247\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3247\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\
        );

    \I__478\ : InMux
    port map (
            O => \N__3244\,
            I => \N__3241\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3241\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__3238\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_\
        );

    \I__475\ : CascadeMux
    port map (
            O => \N__3235\,
            I => \N__3225\
        );

    \I__474\ : InMux
    port map (
            O => \N__3234\,
            I => \N__3220\
        );

    \I__473\ : InMux
    port map (
            O => \N__3233\,
            I => \N__3220\
        );

    \I__472\ : InMux
    port map (
            O => \N__3232\,
            I => \N__3217\
        );

    \I__471\ : InMux
    port map (
            O => \N__3231\,
            I => \N__3212\
        );

    \I__470\ : InMux
    port map (
            O => \N__3230\,
            I => \N__3212\
        );

    \I__469\ : InMux
    port map (
            O => \N__3229\,
            I => \N__3205\
        );

    \I__468\ : InMux
    port map (
            O => \N__3228\,
            I => \N__3205\
        );

    \I__467\ : InMux
    port map (
            O => \N__3225\,
            I => \N__3205\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3220\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3217\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3212\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__3205\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__462\ : InMux
    port map (
            O => \N__3196\,
            I => \N__3187\
        );

    \I__461\ : InMux
    port map (
            O => \N__3195\,
            I => \N__3180\
        );

    \I__460\ : InMux
    port map (
            O => \N__3194\,
            I => \N__3180\
        );

    \I__459\ : InMux
    port map (
            O => \N__3193\,
            I => \N__3180\
        );

    \I__458\ : InMux
    port map (
            O => \N__3192\,
            I => \N__3173\
        );

    \I__457\ : InMux
    port map (
            O => \N__3191\,
            I => \N__3173\
        );

    \I__456\ : InMux
    port map (
            O => \N__3190\,
            I => \N__3173\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__3187\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__3180\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3173\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__452\ : InMux
    port map (
            O => \N__3166\,
            I => \N__3163\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__3163\,
            I => \N__3159\
        );

    \I__450\ : InMux
    port map (
            O => \N__3162\,
            I => \N__3156\
        );

    \I__449\ : Span12Mux_v
    port map (
            O => \N__3159\,
            I => \N__3151\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3156\,
            I => \N__3151\
        );

    \I__447\ : Odrv12
    port map (
            O => \N__3151\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\
        );

    \I__446\ : IoInMux
    port map (
            O => \N__3148\,
            I => \N__3145\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3145\,
            I => \N__3142\
        );

    \I__444\ : IoSpan4Mux
    port map (
            O => \N__3142\,
            I => \N__3139\
        );

    \I__443\ : Span4Mux_s3_v
    port map (
            O => \N__3139\,
            I => \N__3136\
        );

    \I__442\ : Sp12to4
    port map (
            O => \N__3136\,
            I => \N__3133\
        );

    \I__441\ : Span12Mux_s11_v
    port map (
            O => \N__3133\,
            I => \N__3130\
        );

    \I__440\ : Odrv12
    port map (
            O => \N__3130\,
            I => \U409_ADDRESS_DECODE_un1_nREGSPACE_i\
        );

    \I__439\ : InMux
    port map (
            O => \N__3127\,
            I => \N__3124\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__3124\,
            I => \N__3121\
        );

    \I__437\ : Span4Mux_v
    port map (
            O => \N__3121\,
            I => \N__3118\
        );

    \I__436\ : Sp12to4
    port map (
            O => \N__3118\,
            I => \N__3115\
        );

    \I__435\ : Span12Mux_h
    port map (
            O => \N__3115\,
            I => \N__3112\
        );

    \I__434\ : Odrv12
    port map (
            O => \N__3112\,
            I => \A_c_13\
        );

    \I__433\ : IoInMux
    port map (
            O => \N__3109\,
            I => \N__3106\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__3106\,
            I => \N__3103\
        );

    \I__431\ : Span4Mux_s1_h
    port map (
            O => \N__3103\,
            I => \N__3100\
        );

    \I__430\ : Sp12to4
    port map (
            O => \N__3100\,
            I => \N__3097\
        );

    \I__429\ : Span12Mux_s9_v
    port map (
            O => \N__3097\,
            I => \N__3094\
        );

    \I__428\ : Span12Mux_h
    port map (
            O => \N__3094\,
            I => \N__3091\
        );

    \I__427\ : Odrv12
    port map (
            O => \N__3091\,
            I => \U409_ADDRESS_DECODE_un1_nCIACS1_i\
        );

    \I__426\ : InMux
    port map (
            O => \N__3088\,
            I => \N__3085\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3085\,
            I => \N__3082\
        );

    \I__424\ : Span12Mux_h
    port map (
            O => \N__3082\,
            I => \N__3079\
        );

    \I__423\ : Odrv12
    port map (
            O => \N__3079\,
            I => \A_c_12\
        );

    \I__422\ : IoInMux
    port map (
            O => \N__3076\,
            I => \N__3073\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3073\,
            I => \N__3070\
        );

    \I__420\ : Span4Mux_s1_h
    port map (
            O => \N__3070\,
            I => \N__3067\
        );

    \I__419\ : Sp12to4
    port map (
            O => \N__3067\,
            I => \N__3064\
        );

    \I__418\ : Span12Mux_s10_v
    port map (
            O => \N__3064\,
            I => \N__3061\
        );

    \I__417\ : Span12Mux_h
    port map (
            O => \N__3061\,
            I => \N__3058\
        );

    \I__416\ : Odrv12
    port map (
            O => \N__3058\,
            I => \U409_ADDRESS_DECODE_un1_nCIACS0_i\
        );

    \I__415\ : CascadeMux
    port map (
            O => \N__3055\,
            I => \U409_CIA.N_9_cascade_\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__3052\,
            I => \U409_CIA.N_20_cascade_\
        );

    \I__413\ : InMux
    port map (
            O => \N__3049\,
            I => \N__3043\
        );

    \I__412\ : InMux
    port map (
            O => \N__3048\,
            I => \N__3043\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__3043\,
            I => \U409_CIA.CLKCIA8_0_a2_0\
        );

    \I__410\ : InMux
    port map (
            O => \N__3040\,
            I => \N__3037\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3037\,
            I => \U409_CIA.CLKCIA6_0_a2_1\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__3034\,
            I => \U409_CIA.CLKCIAZ0_cascade_\
        );

    \I__407\ : InMux
    port map (
            O => \N__3031\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__406\ : InMux
    port map (
            O => \N__3028\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__405\ : InMux
    port map (
            O => \N__3025\,
            I => \bfn_8_9_0_\
        );

    \I__404\ : InMux
    port map (
            O => \N__3022\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__403\ : InMux
    port map (
            O => \N__3019\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__402\ : InMux
    port map (
            O => \N__3016\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__401\ : InMux
    port map (
            O => \N__3013\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__400\ : InMux
    port map (
            O => \N__3010\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__399\ : InMux
    port map (
            O => \N__3007\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__398\ : InMux
    port map (
            O => \N__3004\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__397\ : InMux
    port map (
            O => \N__3001\,
            I => \N__2998\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2998\,
            I => \N__2995\
        );

    \I__395\ : Span4Mux_h
    port map (
            O => \N__2995\,
            I => \N__2992\
        );

    \I__394\ : Odrv4
    port map (
            O => \N__2992\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\
        );

    \I__393\ : IoInMux
    port map (
            O => \N__2989\,
            I => \N__2986\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2986\,
            I => \N__2983\
        );

    \I__391\ : IoSpan4Mux
    port map (
            O => \N__2983\,
            I => \N__2980\
        );

    \I__390\ : Sp12to4
    port map (
            O => \N__2980\,
            I => \N__2977\
        );

    \I__389\ : Span12Mux_v
    port map (
            O => \N__2977\,
            I => \N__2974\
        );

    \I__388\ : Odrv12
    port map (
            O => \N__2974\,
            I => \PORTSIZE_0_i\
        );

    \I__387\ : InMux
    port map (
            O => \N__2971\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__386\ : InMux
    port map (
            O => \N__2968\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__385\ : InMux
    port map (
            O => \N__2965\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__384\ : InMux
    port map (
            O => \N__2962\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__383\ : InMux
    port map (
            O => \N__2959\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__382\ : InMux
    port map (
            O => \N__2956\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__381\ : InMux
    port map (
            O => \N__2953\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__380\ : InMux
    port map (
            O => \N__2950\,
            I => \N__2941\
        );

    \I__379\ : InMux
    port map (
            O => \N__2949\,
            I => \N__2941\
        );

    \I__378\ : InMux
    port map (
            O => \N__2948\,
            I => \N__2941\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2941\,
            I => \N__2938\
        );

    \I__376\ : Span12Mux_v
    port map (
            O => \N__2938\,
            I => \N__2935\
        );

    \I__375\ : Odrv12
    port map (
            O => \N__2935\,
            I => \A_c_29\
        );

    \I__374\ : InMux
    port map (
            O => \N__2932\,
            I => \N__2927\
        );

    \I__373\ : InMux
    port map (
            O => \N__2931\,
            I => \N__2922\
        );

    \I__372\ : InMux
    port map (
            O => \N__2930\,
            I => \N__2922\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2927\,
            I => \N__2917\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2922\,
            I => \N__2917\
        );

    \I__369\ : Span4Mux_h
    port map (
            O => \N__2917\,
            I => \N__2914\
        );

    \I__368\ : Span4Mux_v
    port map (
            O => \N__2914\,
            I => \N__2911\
        );

    \I__367\ : Span4Mux_v
    port map (
            O => \N__2911\,
            I => \N__2908\
        );

    \I__366\ : Odrv4
    port map (
            O => \N__2908\,
            I => \A_c_28\
        );

    \I__365\ : CascadeMux
    port map (
            O => \N__2905\,
            I => \N__2902\
        );

    \I__364\ : InMux
    port map (
            O => \N__2902\,
            I => \N__2897\
        );

    \I__363\ : InMux
    port map (
            O => \N__2901\,
            I => \N__2894\
        );

    \I__362\ : InMux
    port map (
            O => \N__2900\,
            I => \N__2891\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2897\,
            I => \N__2884\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2894\,
            I => \N__2884\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2891\,
            I => \N__2884\
        );

    \I__358\ : Odrv12
    port map (
            O => \N__2884\,
            I => \A_c_27\
        );

    \I__357\ : CascadeMux
    port map (
            O => \N__2881\,
            I => \N__2877\
        );

    \I__356\ : InMux
    port map (
            O => \N__2880\,
            I => \N__2869\
        );

    \I__355\ : InMux
    port map (
            O => \N__2877\,
            I => \N__2869\
        );

    \I__354\ : InMux
    port map (
            O => \N__2876\,
            I => \N__2869\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2869\,
            I => \N__2866\
        );

    \I__352\ : Span12Mux_v
    port map (
            O => \N__2866\,
            I => \N__2863\
        );

    \I__351\ : Odrv12
    port map (
            O => \N__2863\,
            I => \A_c_30\
        );

    \I__350\ : InMux
    port map (
            O => \N__2860\,
            I => \N__2857\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2857\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_10\
        );

    \I__348\ : InMux
    port map (
            O => \N__2854\,
            I => \N__2848\
        );

    \I__347\ : InMux
    port map (
            O => \N__2853\,
            I => \N__2848\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2848\,
            I => \N__2845\
        );

    \I__345\ : Span4Mux_v
    port map (
            O => \N__2845\,
            I => \N__2841\
        );

    \I__344\ : InMux
    port map (
            O => \N__2844\,
            I => \N__2838\
        );

    \I__343\ : Sp12to4
    port map (
            O => \N__2841\,
            I => \N__2833\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2838\,
            I => \N__2833\
        );

    \I__341\ : Odrv12
    port map (
            O => \N__2833\,
            I => \A_c_20\
        );

    \I__340\ : CascadeMux
    port map (
            O => \N__2830\,
            I => \N__2826\
        );

    \I__339\ : InMux
    port map (
            O => \N__2829\,
            I => \N__2822\
        );

    \I__338\ : InMux
    port map (
            O => \N__2826\,
            I => \N__2819\
        );

    \I__337\ : InMux
    port map (
            O => \N__2825\,
            I => \N__2816\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2822\,
            I => \N__2811\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__2819\,
            I => \N__2811\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2816\,
            I => \N__2808\
        );

    \I__333\ : Span4Mux_v
    port map (
            O => \N__2811\,
            I => \N__2805\
        );

    \I__332\ : Odrv12
    port map (
            O => \N__2808\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEm_6\
        );

    \I__331\ : Odrv4
    port map (
            O => \N__2805\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEm_6\
        );

    \I__330\ : InMux
    port map (
            O => \N__2800\,
            I => \N__2795\
        );

    \I__329\ : InMux
    port map (
            O => \N__2799\,
            I => \N__2790\
        );

    \I__328\ : InMux
    port map (
            O => \N__2798\,
            I => \N__2790\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2795\,
            I => \N__2787\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2790\,
            I => \N__2784\
        );

    \I__325\ : Span4Mux_v
    port map (
            O => \N__2787\,
            I => \N__2781\
        );

    \I__324\ : Span4Mux_v
    port map (
            O => \N__2784\,
            I => \N__2778\
        );

    \I__323\ : Span4Mux_h
    port map (
            O => \N__2781\,
            I => \N__2775\
        );

    \I__322\ : Sp12to4
    port map (
            O => \N__2778\,
            I => \N__2772\
        );

    \I__321\ : Sp12to4
    port map (
            O => \N__2775\,
            I => \N__2767\
        );

    \I__320\ : Span12Mux_s3_h
    port map (
            O => \N__2772\,
            I => \N__2767\
        );

    \I__319\ : Span12Mux_v
    port map (
            O => \N__2767\,
            I => \N__2764\
        );

    \I__318\ : Odrv12
    port map (
            O => \N__2764\,
            I => \A_c_19\
        );

    \I__317\ : CascadeMux
    port map (
            O => \N__2761\,
            I => \N__2757\
        );

    \I__316\ : CascadeMux
    port map (
            O => \N__2760\,
            I => \N__2754\
        );

    \I__315\ : InMux
    port map (
            O => \N__2757\,
            I => \N__2748\
        );

    \I__314\ : InMux
    port map (
            O => \N__2754\,
            I => \N__2748\
        );

    \I__313\ : CascadeMux
    port map (
            O => \N__2753\,
            I => \N__2745\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2748\,
            I => \N__2742\
        );

    \I__311\ : InMux
    port map (
            O => \N__2745\,
            I => \N__2739\
        );

    \I__310\ : Odrv4
    port map (
            O => \N__2742\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEm_3\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2739\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEm_3\
        );

    \I__308\ : InMux
    port map (
            O => \N__2734\,
            I => \N__2731\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2731\,
            I => \N__2728\
        );

    \I__306\ : Span4Mux_v
    port map (
            O => \N__2728\,
            I => \N__2725\
        );

    \I__305\ : Span4Mux_v
    port map (
            O => \N__2725\,
            I => \N__2722\
        );

    \I__304\ : IoSpan4Mux
    port map (
            O => \N__2722\,
            I => \N__2719\
        );

    \I__303\ : Odrv4
    port map (
            O => \N__2719\,
            I => \TT_c_1\
        );

    \I__302\ : InMux
    port map (
            O => \N__2716\,
            I => \N__2713\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2713\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8\
        );

    \I__300\ : InMux
    port map (
            O => \N__2710\,
            I => \N__2707\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2707\,
            I => \N__2704\
        );

    \I__298\ : Span4Mux_h
    port map (
            O => \N__2704\,
            I => \N__2701\
        );

    \I__297\ : Span4Mux_v
    port map (
            O => \N__2701\,
            I => \N__2696\
        );

    \I__296\ : InMux
    port map (
            O => \N__2700\,
            I => \N__2691\
        );

    \I__295\ : InMux
    port map (
            O => \N__2699\,
            I => \N__2691\
        );

    \I__294\ : Sp12to4
    port map (
            O => \N__2696\,
            I => \N__2686\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2691\,
            I => \N__2686\
        );

    \I__292\ : Odrv12
    port map (
            O => \N__2686\,
            I => \A_c_25\
        );

    \I__291\ : CascadeMux
    port map (
            O => \N__2683\,
            I => \N__2679\
        );

    \I__290\ : CascadeMux
    port map (
            O => \N__2682\,
            I => \N__2675\
        );

    \I__289\ : InMux
    port map (
            O => \N__2679\,
            I => \N__2672\
        );

    \I__288\ : InMux
    port map (
            O => \N__2678\,
            I => \N__2667\
        );

    \I__287\ : InMux
    port map (
            O => \N__2675\,
            I => \N__2667\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2672\,
            I => \N__2662\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2667\,
            I => \N__2662\
        );

    \I__284\ : Span4Mux_v
    port map (
            O => \N__2662\,
            I => \N__2659\
        );

    \I__283\ : Span4Mux_v
    port map (
            O => \N__2659\,
            I => \N__2656\
        );

    \I__282\ : Sp12to4
    port map (
            O => \N__2656\,
            I => \N__2653\
        );

    \I__281\ : Odrv12
    port map (
            O => \N__2653\,
            I => \A_c_24\
        );

    \I__280\ : InMux
    port map (
            O => \N__2650\,
            I => \N__2641\
        );

    \I__279\ : InMux
    port map (
            O => \N__2649\,
            I => \N__2641\
        );

    \I__278\ : InMux
    port map (
            O => \N__2648\,
            I => \N__2641\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2641\,
            I => \N__2638\
        );

    \I__276\ : Span4Mux_v
    port map (
            O => \N__2638\,
            I => \N__2635\
        );

    \I__275\ : Span4Mux_v
    port map (
            O => \N__2635\,
            I => \N__2632\
        );

    \I__274\ : Span4Mux_h
    port map (
            O => \N__2632\,
            I => \N__2629\
        );

    \I__273\ : Odrv4
    port map (
            O => \N__2629\,
            I => \A_c_26\
        );

    \I__272\ : CascadeMux
    port map (
            O => \N__2626\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_\
        );

    \I__271\ : InMux
    port map (
            O => \N__2623\,
            I => \N__2620\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2620\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\
        );

    \I__269\ : InMux
    port map (
            O => \N__2617\,
            I => \N__2614\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2614\,
            I => \N__2611\
        );

    \I__267\ : Span12Mux_v
    port map (
            O => \N__2611\,
            I => \N__2608\
        );

    \I__266\ : Odrv12
    port map (
            O => \N__2608\,
            I => \TT_c_0\
        );

    \I__265\ : CascadeMux
    port map (
            O => \N__2605\,
            I => \N__2600\
        );

    \I__264\ : InMux
    port map (
            O => \N__2604\,
            I => \N__2595\
        );

    \I__263\ : InMux
    port map (
            O => \N__2603\,
            I => \N__2595\
        );

    \I__262\ : InMux
    port map (
            O => \N__2600\,
            I => \N__2592\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2595\,
            I => \N__2589\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2592\,
            I => \N__2586\
        );

    \I__259\ : Span4Mux_v
    port map (
            O => \N__2589\,
            I => \N__2583\
        );

    \I__258\ : Span4Mux_v
    port map (
            O => \N__2586\,
            I => \N__2580\
        );

    \I__257\ : Sp12to4
    port map (
            O => \N__2583\,
            I => \N__2575\
        );

    \I__256\ : Sp12to4
    port map (
            O => \N__2580\,
            I => \N__2575\
        );

    \I__255\ : Odrv12
    port map (
            O => \N__2575\,
            I => \A_c_31\
        );

    \I__254\ : InMux
    port map (
            O => \N__2572\,
            I => \N__2569\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__2569\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9\
        );

    \I__252\ : CascadeMux
    port map (
            O => \N__2566\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7_cascade_\
        );

    \I__251\ : InMux
    port map (
            O => \N__2563\,
            I => \N__2560\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2560\,
            I => \U409_CIA.g0Z0Z_10\
        );

    \I__249\ : CascadeMux
    port map (
            O => \N__2557\,
            I => \U409_CIA.g0Z0Z_2_cascade_\
        );

    \I__248\ : InMux
    port map (
            O => \N__2554\,
            I => \N__2548\
        );

    \I__247\ : InMux
    port map (
            O => \N__2553\,
            I => \N__2548\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__2548\,
            I => \N__2545\
        );

    \I__245\ : Span4Mux_v
    port map (
            O => \N__2545\,
            I => \N__2542\
        );

    \I__244\ : Sp12to4
    port map (
            O => \N__2542\,
            I => \N__2539\
        );

    \I__243\ : Span12Mux_s7_h
    port map (
            O => \N__2539\,
            I => \N__2536\
        );

    \I__242\ : Span12Mux_v
    port map (
            O => \N__2536\,
            I => \N__2533\
        );

    \I__241\ : Odrv12
    port map (
            O => \N__2533\,
            I => \A_c_18\
        );

    \I__240\ : CascadeMux
    port map (
            O => \N__2530\,
            I => \N__2526\
        );

    \I__239\ : InMux
    port map (
            O => \N__2529\,
            I => \N__2521\
        );

    \I__238\ : InMux
    port map (
            O => \N__2526\,
            I => \N__2521\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__2521\,
            I => \N__2518\
        );

    \I__236\ : Span4Mux_v
    port map (
            O => \N__2518\,
            I => \N__2515\
        );

    \I__235\ : Sp12to4
    port map (
            O => \N__2515\,
            I => \N__2512\
        );

    \I__234\ : Span12Mux_v
    port map (
            O => \N__2512\,
            I => \N__2509\
        );

    \I__233\ : Odrv12
    port map (
            O => \N__2509\,
            I => \A_c_17\
        );

    \I__232\ : InMux
    port map (
            O => \N__2506\,
            I => \N__2500\
        );

    \I__231\ : InMux
    port map (
            O => \N__2505\,
            I => \N__2500\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__2500\,
            I => \N__2497\
        );

    \I__229\ : Span4Mux_v
    port map (
            O => \N__2497\,
            I => \N__2494\
        );

    \I__228\ : Sp12to4
    port map (
            O => \N__2494\,
            I => \N__2491\
        );

    \I__227\ : Span12Mux_s3_h
    port map (
            O => \N__2491\,
            I => \N__2488\
        );

    \I__226\ : Span12Mux_v
    port map (
            O => \N__2488\,
            I => \N__2485\
        );

    \I__225\ : Odrv12
    port map (
            O => \N__2485\,
            I => \A_c_16\
        );

    \I__224\ : CascadeMux
    port map (
            O => \N__2482\,
            I => \U409_CIA.g0Z0Z_8_cascade_\
        );

    \I__223\ : InMux
    port map (
            O => \N__2479\,
            I => \N__2476\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__2476\,
            I => \U409_CIA.g0Z0Z_11\
        );

    \I__221\ : ClkMux
    port map (
            O => \N__2473\,
            I => \N__2446\
        );

    \I__220\ : ClkMux
    port map (
            O => \N__2472\,
            I => \N__2446\
        );

    \I__219\ : ClkMux
    port map (
            O => \N__2471\,
            I => \N__2446\
        );

    \I__218\ : ClkMux
    port map (
            O => \N__2470\,
            I => \N__2446\
        );

    \I__217\ : ClkMux
    port map (
            O => \N__2469\,
            I => \N__2446\
        );

    \I__216\ : ClkMux
    port map (
            O => \N__2468\,
            I => \N__2446\
        );

    \I__215\ : ClkMux
    port map (
            O => \N__2467\,
            I => \N__2446\
        );

    \I__214\ : ClkMux
    port map (
            O => \N__2466\,
            I => \N__2446\
        );

    \I__213\ : ClkMux
    port map (
            O => \N__2465\,
            I => \N__2446\
        );

    \I__212\ : GlobalMux
    port map (
            O => \N__2446\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.TACK_EN_iC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            I => \N__2468\
        );

    \INVU409_TRANSFER_ACK.TACK_OUTnC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            I => \N__2466\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            I => \N__2465\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            I => \N__2472\
        );

    \INVU409_TRANSFER_ACK.CIA_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            I => \N__2470\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            I => \N__2467\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            I => \N__2473\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__2471\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            I => \N__2469\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_12_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_12_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2798\,
            in1 => \N__2553\,
            in2 => \N__2530\,
            in3 => \N__2505\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_11_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2710\,
            in1 => \N__2844\,
            in2 => \N__3945\,
            in3 => \N__2554\,
            lcout => \U409_CIA.g0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_8_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2529\,
            in1 => \N__4028\,
            in2 => \_gnd_net_\,
            in3 => \N__5857\,
            lcout => OPEN,
            ltout => \U409_CIA.g0Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_14_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2506\,
            in1 => \N__2799\,
            in2 => \N__2482\,
            in3 => \N__2479\,
            lcout => \U409_CIA.g0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2648\,
            in1 => \N__2699\,
            in2 => \N__2682\,
            in3 => \N__2825\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_10_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2901\,
            in1 => \N__2678\,
            in2 => \N__2605\,
            in3 => \N__2650\,
            lcout => \U409_CIA.g0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2700\,
            in1 => \N__2900\,
            in2 => \N__2683\,
            in3 => \N__2649\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__2604\,
            in1 => \_gnd_net_\,
            in2 => \N__2881\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__2949\,
            in1 => \N__2931\,
            in2 => \N__2626\,
            in3 => \N__2623\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5860\,
            in1 => \N__2617\,
            in2 => \_gnd_net_\,
            in3 => \N__2603\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2860\,
            in1 => \N__2572\,
            in2 => \N__2566\,
            in3 => \N__2716\,
            lcout => \AUTOVECTORm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_2_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__2950\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2880\,
            lcout => OPEN,
            ltout => \U409_CIA.g0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_13_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__2563\,
            in1 => \N__2932\,
            in2 => \N__2557\,
            in3 => \N__4067\,
            lcout => \U409_CIA.g0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_10_0_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2948\,
            in1 => \N__2930\,
            in2 => \N__2905\,
            in3 => \N__2876\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.HIROM_0_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3943\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2853\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEm_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__2854\,
            in1 => \N__4105\,
            in2 => \N__2830\,
            in3 => \N__3944\,
            lcout => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__4104\,
            in1 => \N__4367\,
            in2 => \N__2753\,
            in3 => \N__2829\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.HIROM_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4095\,
            in1 => \N__4030\,
            in2 => \N__2761\,
            in3 => \N__2800\,
            lcout => \U409_ADDRESS_DECODE.HIROMZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4094\,
            in1 => \N__4029\,
            in2 => \N__2760\,
            in3 => \N__2734\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4390\,
            in1 => \N__4031\,
            in2 => \_gnd_net_\,
            in3 => \N__3162\,
            lcout => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3233\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3234\,
            in2 => \_gnd_net_\,
            in3 => \N__3277\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5856\,
            in1 => \N__4001\,
            in2 => \N__4437\,
            in3 => \N__3001\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3386\,
            in2 => \N__3414\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3522\,
            in2 => \_gnd_net_\,
            in3 => \N__2971\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__5321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3495\,
            in2 => \_gnd_net_\,
            in3 => \N__2968\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__5321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3753\,
            in2 => \_gnd_net_\,
            in3 => \N__2965\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__5321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3366\,
            in2 => \_gnd_net_\,
            in3 => \N__2962\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3807\,
            in2 => \_gnd_net_\,
            in3 => \N__2959\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3768\,
            in2 => \_gnd_net_\,
            in3 => \N__2956\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__5321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3534\,
            in2 => \_gnd_net_\,
            in3 => \N__2953\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__5321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3717\,
            in2 => \_gnd_net_\,
            in3 => \N__3025\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3462\,
            in2 => \_gnd_net_\,
            in3 => \N__3022\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__5323\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3819\,
            in2 => \_gnd_net_\,
            in3 => \N__3019\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3477\,
            in2 => \_gnd_net_\,
            in3 => \N__3016\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__5323\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3786\,
            in2 => \_gnd_net_\,
            in3 => \N__3013\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3585\,
            in2 => \_gnd_net_\,
            in3 => \N__3010\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3741\,
            in2 => \_gnd_net_\,
            in3 => \N__3007\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3510\,
            in2 => \_gnd_net_\,
            in3 => \N__3004\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5323\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_1_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3300\,
            in1 => \N__3340\,
            in2 => \N__3322\,
            in3 => \N__3195\,
            lcout => \U409_CIA.CLKCIA6_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001000100"
        )
    port map (
            in0 => \N__3275\,
            in1 => \N__3194\,
            in2 => \_gnd_net_\,
            in3 => \N__3232\,
            lcout => OPEN,
            ltout => \U409_CIA.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011101100"
        )
    port map (
            in0 => \N__3049\,
            in1 => \N__4285\,
            in2 => \N__3055\,
            in3 => \N__3196\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__3316\,
            in1 => \N__3339\,
            in2 => \_gnd_net_\,
            in3 => \N__3295\,
            lcout => \U409_CIA.CLKCIA8_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_2_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3193\,
            in1 => \N__3230\,
            in2 => \_gnd_net_\,
            in3 => \N__3274\,
            lcout => OPEN,
            ltout => \U409_CIA.N_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_0_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4928\,
            in2 => \N__3052\,
            in3 => \N__3048\,
            lcout => OPEN,
            ltout => \U409_CIA.CLKCIAZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__3040\,
            in1 => \N__3231\,
            in2 => \N__3034\,
            in3 => \N__3276\,
            lcout => \CLKCIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3272\,
            in2 => \N__3235\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3337\,
            in2 => \_gnd_net_\,
            in3 => \N__3031\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__3552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3190\,
            in2 => \_gnd_net_\,
            in3 => \N__3028\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3296\,
            in2 => \_gnd_net_\,
            in3 => \N__3349\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__3552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3320\,
            in2 => \_gnd_net_\,
            in3 => \N__3346\,
            lcout => OPEN,
            ltout => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__3192\,
            in1 => \N__3250\,
            in2 => \N__3343\,
            in3 => \N__3228\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__3338\,
            in1 => \N__3321\,
            in2 => \N__3301\,
            in3 => \N__3273\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\,
            ltout => \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011001100110"
        )
    port map (
            in0 => \N__3191\,
            in1 => \N__3244\,
            in2 => \N__3238\,
            in3 => \N__3229\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__3166\,
            in1 => \N__4022\,
            in2 => \_gnd_net_\,
            in3 => \N__4395\,
            lcout => \U409_ADDRESS_DECODE_un1_nREGSPACE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__3127\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4123\,
            lcout => \U409_ADDRESS_DECODE_un1_nCIACS1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3088\,
            in2 => \_gnd_net_\,
            in3 => \N__4119\,
            lcout => \U409_ADDRESS_DECODE_un1_nCIACS0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3535\,
            in1 => \N__3523\,
            in2 => \N__3511\,
            in3 => \N__3387\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3367\,
            in1 => \N__3496\,
            in2 => \_gnd_net_\,
            in3 => \N__3409\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3484\,
            in1 => \N__3478\,
            in2 => \N__3466\,
            in3 => \N__3463\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__3706\,
            in1 => \N__3432\,
            in2 => \N__3451\,
            in3 => \N__3633\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3666\,
            in1 => \N__3705\,
            in2 => \N__3637\,
            in3 => \N__3421\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__3703\,
            in1 => \N__3667\,
            in2 => \N__3415\,
            in3 => \N__3631\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3410\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3388\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__3704\,
            in1 => \N__3373\,
            in2 => \N__3676\,
            in3 => \N__3632\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3671\,
            in1 => \N__3699\,
            in2 => \N__3636\,
            in3 => \N__3355\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3820\,
            in1 => \N__3808\,
            in2 => \N__3721\,
            in3 => \N__3787\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3672\,
            in1 => \N__3700\,
            in2 => \N__3796\,
            in3 => \N__3793\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3702\,
            in1 => \N__3674\,
            in2 => \N__3635\,
            in3 => \N__3775\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__3586\,
            in1 => \N__3769\,
            in2 => \N__3757\,
            in3 => \N__3742\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__3624\,
            in1 => \N__3730\,
            in2 => \N__3724\,
            in3 => \N__3675\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3701\,
            in1 => \N__3673\,
            in2 => \N__3634\,
            in3 => \N__3592\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__4394\,
            in1 => \N__4419\,
            in2 => \_gnd_net_\,
            in3 => \N__4317\,
            lcout => \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_HOLD_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__4235\,
            in1 => \N__4256\,
            in2 => \N__4289\,
            in3 => \N__4208\,
            lcout => \U409_CIA.CIA_HOLDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__4236\,
            in1 => \N__4257\,
            in2 => \N__4290\,
            in3 => \N__4209\,
            lcout => \CIA_ENABLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.LOWROM_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4324\,
            in1 => \N__4032\,
            in2 => \N__3955\,
            in3 => \N__4102\,
            lcout => \U409_ADDRESS_DECODE.LOWROMZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__4103\,
            in1 => \_gnd_net_\,
            in2 => \N__4036\,
            in3 => \N__3954\,
            lcout => \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__4840\,
            in1 => \N__3898\,
            in2 => \N__3829\,
            in3 => \N__5100\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMENm_i_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011111111111"
        )
    port map (
            in0 => \N__4386\,
            in1 => \N__3861\,
            in2 => \N__3847\,
            in3 => \N__5859\,
            lcout => \ROMENm_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__5858\,
            in1 => \N__4385\,
            in2 => \N__3862\,
            in3 => \N__3843\,
            lcout => \ROMENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__4180\,
            in1 => \N__4145\,
            in2 => \N__4453\,
            in3 => \N__4627\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__5668\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4734\,
            in2 => \_gnd_net_\,
            in3 => \N__4798\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4662\,
            in1 => \N__4684\,
            in2 => \N__4606\,
            in3 => \N__4178\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4765\,
            in1 => \N__4146\,
            in2 => \N__4183\,
            in3 => \N__4161\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4179\,
            in1 => \N__4685\,
            in2 => \N__4778\,
            in3 => \N__4144\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4663\,
            in1 => \N__4603\,
            in2 => \N__4165\,
            in3 => \N__4162\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__4838\,
            in1 => \N__5103\,
            in2 => \N__4153\,
            in3 => \N__4706\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4449\,
            in2 => \N__4150\,
            in3 => \N__4147\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__5668\
        );

    \RESETn_ibuf_RNIM9SF_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5838\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100000111"
        )
    port map (
            in0 => \N__4965\,
            in1 => \N__4991\,
            in2 => \N__5035\,
            in3 => \N__5001\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.m9_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010010001100"
        )
    port map (
            in0 => \N__5133\,
            in1 => \N__5840\,
            in2 => \N__4129\,
            in3 => \N__5008\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000110111"
        )
    port map (
            in0 => \N__4992\,
            in1 => \N__5131\,
            in2 => \N__4969\,
            in3 => \N__5002\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.i6_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010001000"
        )
    port map (
            in0 => \N__5132\,
            in1 => \N__5841\,
            in2 => \N__4126\,
            in3 => \N__5032\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__4441\,
            in1 => \N__4420\,
            in2 => \N__4402\,
            in3 => \N__4316\,
            lcout => \nBUFEN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__4291\,
            in1 => \N__4261\,
            in2 => \N__4240\,
            in3 => \N__4210\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__5558\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5236\,
            in1 => \N__5257\,
            in2 => \_gnd_net_\,
            in3 => \N__4858\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4189\,
            in1 => \N__5428\,
            in2 => \N__4195\,
            in3 => \N__5275\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__4547\,
            in1 => \N__4486\,
            in2 => \N__4192\,
            in3 => \N__4859\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5334\,
            in1 => \N__4875\,
            in2 => \N__5293\,
            in3 => \N__5413\,
            lcout => \U409_TICK.TICK603_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__4548\,
            in1 => \N__5245\,
            in2 => \N__4522\,
            in3 => \N__4487\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5380\,
            in1 => \N__5185\,
            in2 => \N__5161\,
            in3 => \N__5221\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4549\,
            in1 => \N__4521\,
            in2 => \N__4582\,
            in3 => \N__5209\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__4860\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4876\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4514\,
            in1 => \N__4546\,
            in2 => \N__5146\,
            in3 => \N__4484\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4544\,
            in1 => \N__4517\,
            in2 => \N__4489\,
            in3 => \N__5347\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4513\,
            in1 => \N__4545\,
            in2 => \N__5173\,
            in3 => \N__4483\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__5359\,
            in1 => \N__5443\,
            in2 => \N__5398\,
            in3 => \N__5200\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => \U409_TICK.TICK603_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__4515\,
            in1 => \N__4560\,
            in2 => \N__4579\,
            in3 => \N__4485\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4543\,
            in1 => \N__4516\,
            in2 => \N__4488\,
            in3 => \N__5368\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4686\,
            in1 => \N__4799\,
            in2 => \N__4779\,
            in3 => \N__4735\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4604\,
            in2 => \N__4456\,
            in3 => \N__4664\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4772\,
            in1 => \N__4800\,
            in2 => \_gnd_net_\,
            in3 => \N__4736\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100000101"
        )
    port map (
            in0 => \N__4708\,
            in1 => \N__4839\,
            in2 => \N__4780\,
            in3 => \N__5102\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5664\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__4737\,
            in1 => \N__4774\,
            in2 => \_gnd_net_\,
            in3 => \N__4801\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5664\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4773\,
            in1 => \N__4738\,
            in2 => \_gnd_net_\,
            in3 => \N__4625\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5664\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__4714\,
            in1 => \N__5458\,
            in2 => \_gnd_net_\,
            in3 => \N__4707\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5664\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4693\,
            in1 => \N__4687\,
            in2 => \_gnd_net_\,
            in3 => \N__4624\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5664\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4623\,
            in1 => \N__4635\,
            in2 => \_gnd_net_\,
            in3 => \N__4666\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5664\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__4665\,
            in1 => \N__4605\,
            in2 => \N__4639\,
            in3 => \N__4626\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5664\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011101000000"
        )
    port map (
            in0 => \N__5034\,
            in1 => \N__5134\,
            in2 => \N__5044\,
            in3 => \N__5473\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5548\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__5130\,
            in1 => \N__4900\,
            in2 => \N__5101\,
            in3 => \N__4914\,
            lcout => \U409_TRANSFER_ACK.N_107\,
            ltout => \U409_TRANSFER_ACK.N_107_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100100111"
        )
    port map (
            in0 => \N__5033\,
            in1 => \N__4959\,
            in2 => \N__5011\,
            in3 => \N__4990\,
            lcout => \U409_TRANSFER_ACK.m9_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4899\,
            in2 => \_gnd_net_\,
            in3 => \N__4913\,
            lcout => \U409_TRANSFER_ACK.N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4993\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            ce => 'H',
            sr => \N__5559\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4935\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            ce => 'H',
            sr => \N__5559\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4915\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            ce => 'H',
            sr => \N__5559\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4874\,
            in2 => \N__4861\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5289\,
            in2 => \_gnd_net_\,
            in3 => \N__5278\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__5316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5271\,
            in2 => \_gnd_net_\,
            in3 => \N__5260\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__5316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5256\,
            in2 => \_gnd_net_\,
            in3 => \N__5239\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5235\,
            in2 => \_gnd_net_\,
            in3 => \N__5224\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__5316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5220\,
            in2 => \_gnd_net_\,
            in3 => \N__5203\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5199\,
            in2 => \_gnd_net_\,
            in3 => \N__5188\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__5316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5184\,
            in2 => \_gnd_net_\,
            in3 => \N__5164\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5157\,
            in2 => \_gnd_net_\,
            in3 => \N__5137\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_7_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5442\,
            in2 => \_gnd_net_\,
            in3 => \N__5431\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__5318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5427\,
            in2 => \_gnd_net_\,
            in3 => \N__5416\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__5318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5412\,
            in2 => \_gnd_net_\,
            in3 => \N__5401\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__5318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5394\,
            in2 => \_gnd_net_\,
            in3 => \N__5383\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__5318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5379\,
            in2 => \_gnd_net_\,
            in3 => \N__5362\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5358\,
            in2 => \_gnd_net_\,
            in3 => \N__5341\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5335\,
            in2 => \_gnd_net_\,
            in3 => \N__5338\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001100"
        )
    port map (
            in0 => \N__5612\,
            in1 => \N__5490\,
            in2 => \_gnd_net_\,
            in3 => \N__5596\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_EN_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110100"
        )
    port map (
            in0 => \N__5575\,
            in1 => \N__5644\,
            in2 => \N__5494\,
            in3 => \N__5637\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5560\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001100"
        )
    port map (
            in0 => \N__5580\,
            in1 => \N__5614\,
            in2 => \N__5638\,
            in3 => \N__5599\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5560\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010000"
        )
    port map (
            in0 => \N__5598\,
            in1 => \_gnd_net_\,
            in2 => \N__5581\,
            in3 => \N__5633\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5560\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__5579\,
            in1 => \N__5613\,
            in2 => \_gnd_net_\,
            in3 => \N__5597\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5560\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__5925\,
            in1 => \N__5817\,
            in2 => \_gnd_net_\,
            in3 => \N__5937\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011101010"
        )
    port map (
            in0 => \N__5505\,
            in1 => \N__5926\,
            in2 => \N__5839\,
            in3 => \N__5914\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNI7KT7_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5489\,
            in2 => \_gnd_net_\,
            in3 => \N__5472\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIURL11_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__5924\,
            in1 => \N__5936\,
            in2 => \N__5461\,
            in3 => \N__5457\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5446\,
            in3 => \N__5792\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5938\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5793\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5804\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5913\,
            lcout => \TACK_EN_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            ce => \N__5902\,
            sr => \_gnd_net_\
        );

    \TACKn_iobuf_RNO_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5890\,
            lcout => \N_373_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__5788\,
            in1 => \N__5706\,
            in2 => \_gnd_net_\,
            in3 => \N__5689\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     May 31 2025 14:22:48

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U111_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U111_TOP
entity U111_TOP is
port (
    D_UU_AMIGA : inout std_logic_vector(7 downto 0);
    D_LL_AMIGA : inout std_logic_vector(7 downto 0);
    D_UM_AMIGA : inout std_logic_vector(7 downto 0);
    D_LM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_040 : inout std_logic_vector(7 downto 0);
    D_LM_040 : inout std_logic_vector(7 downto 0);
    D_UM_040 : inout std_logic_vector(7 downto 0);
    D_LL_040 : inout std_logic_vector(7 downto 0);
    A_AMIGA : out std_logic_vector(1 downto 0);
    A_040 : in std_logic_vector(1 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    TEAn : in std_logic;
    TSn : out std_logic;
    RESETn : in std_logic;
    CLKRAMA : out std_logic;
    PORTSIZE : in std_logic;
    TEA_CPUn : out std_logic;
    LBENn : in std_logic;
    CLK40B : out std_logic;
    TBI_CPUn : out std_logic;
    TAn : inout std_logic;
    CPUBGn : out std_logic;
    BUFENn : out std_logic;
    RnW : in std_logic;
    CLK80_CPU : out std_logic;
    BUFDIR : out std_logic;
    TCI_CPUn : out std_logic;
    TS_CPUn : in std_logic;
    CLKRAMB : out std_logic;
    CLK40A : out std_logic;
    TCIn : in std_logic;
    TBIn : in std_logic;
    DMAn : out std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    TACKn : inout std_logic;
    BGn : in std_logic);
end U111_TOP;

-- Architecture of U111_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U111_TOP is

signal \N__13729\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \TCIn_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \TAn_in\ : std_logic;
signal \N_240_i\ : std_logic;
signal \N_237_i\ : std_logic;
signal \N_239_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep26_i_ess\ : std_logic;
signal \N_238_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep24_i_ess\ : std_logic;
signal \N_242_i\ : std_logic;
signal \N_243_i\ : std_logic;
signal \N_229_i\ : std_logic;
signal \N_244_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep29_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep17_i_ess\ : std_logic;
signal \N_230_i\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_0\ : std_logic;
signal \N_221_i\ : std_logic;
signal \N_223_i\ : std_logic;
signal \N_233_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep10_i_ess\ : std_logic;
signal \N_234_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep9_i_ess\ : std_logic;
signal \N_222_i\ : std_logic;
signal \N_236_i\ : std_logic;
signal \N_235_i\ : std_logic;
signal \N_224_i\ : std_logic;
signal \N_227_i\ : std_logic;
signal \N_214_i\ : std_logic;
signal \N_228_i\ : std_logic;
signal \N_225_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep15_i_ess\ : std_logic;
signal \N_241_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep25_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep30_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep16_i_ess\ : std_logic;
signal \N_232_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep8_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep20_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep11_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep22_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep14_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep1_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep12_i_ess\ : std_logic;
signal \N_216_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep5_i_ess\ : std_logic;
signal \N_218_i\ : std_logic;
signal \A_040_c_0\ : std_logic;
signal \A_AMIGA_c_0\ : std_logic;
signal \U111_CYCLE_SM_A_AMIGA_0_i_1\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep28_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep27_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep19_i_ess\ : std_logic;
signal \N_231_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep18_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep21_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep23_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep7_i_ess\ : std_logic;
signal \N_220_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep3_i_ess\ : std_logic;
signal \N_219_i\ : std_logic;
signal \D_LL_AMIGA_in_0\ : std_logic;
signal \un2_D_LL_AMIGA_0\ : std_logic;
signal \D_LM_AMIGA_in_1\ : std_logic;
signal \un2_D_LM_AMIGA_1\ : std_logic;
signal \D_UM_040_in_2\ : std_logic;
signal \D_LL_040_in_2\ : std_logic;
signal \un1_D_UM_040_2\ : std_logic;
signal \D_UM_040_in_6\ : std_logic;
signal \D_LL_040_in_6\ : std_logic;
signal \un1_D_UM_040_6\ : std_logic;
signal \D_LM_AMIGA_in_2\ : std_logic;
signal \un2_D_LM_AMIGA_2\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep0_i_ess\ : std_logic;
signal \N_213_i\ : std_logic;
signal \N_226_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep6_i_ess\ : std_logic;
signal \D_LL_AMIGA_in_1\ : std_logic;
signal \un2_D_LL_AMIGA_1\ : std_logic;
signal \A_040_c_1\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep13_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep4_i_ess\ : std_logic;
signal \N_217_i\ : std_logic;
signal \D_LL_AMIGA_in_4\ : std_logic;
signal \un2_D_LL_AMIGA_4\ : std_logic;
signal \D_LL_040_in_0\ : std_logic;
signal \D_UM_040_in_0\ : std_logic;
signal \un1_D_UM_040_0\ : std_logic;
signal \D_LM_AMIGA_in_3\ : std_logic;
signal \un2_D_LM_AMIGA_3\ : std_logic;
signal \LBENn_c_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep2_i_ess\ : std_logic;
signal \N_215_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \D_LL_AMIGA_in_2\ : std_logic;
signal \un2_D_LL_AMIGA_2\ : std_logic;
signal \D_LM_AMIGA_in_0\ : std_logic;
signal \un2_D_LM_AMIGA_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \INVU111_CYCLE_SM.TSnC_net\ : std_logic;
signal \U111_CYCLE_SM.TS_ENZ0\ : std_logic;
signal \D_UM_040_in_1\ : std_logic;
signal \D_LL_040_in_1\ : std_logic;
signal \un1_D_UM_040_1\ : std_logic;
signal \D_LM_AMIGA_in_6\ : std_logic;
signal \un2_D_LM_AMIGA_6\ : std_logic;
signal \D_LM_040_in_1\ : std_logic;
signal \D_UU_040_in_1\ : std_logic;
signal \un1_D_UU_040_1\ : std_logic;
signal \D_LL_040_in_5\ : std_logic;
signal \D_UM_040_in_5\ : std_logic;
signal \un1_D_UM_040_5\ : std_logic;
signal \D_UU_040_in_6\ : std_logic;
signal \D_LM_040_in_6\ : std_logic;
signal \un1_D_UU_040_6\ : std_logic;
signal \D_LL_AMIGA_in_3\ : std_logic;
signal \un2_D_LL_AMIGA_3\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa_cascade_\ : std_logic;
signal \U111_CYCLE_SM.un1_CYCLE_STATE_0\ : std_logic;
signal \U111_CYCLE_SM.TS_EN_6\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U111_CYCLE_SM.FLIP_WORD_2\ : std_logic;
signal \PORTSIZE_c\ : std_logic;
signal \U111_CYCLE_SM.LW_TRANSZ0\ : std_logic;
signal \U111_CYCLE_SM.PORT_MISMATCH_2\ : std_logic;
signal \U111_CYCLE_SM.A2_ENZ0\ : std_logic;
signal \D_LM_AMIGA_in_5\ : std_logic;
signal \un2_D_LM_AMIGA_5\ : std_logic;
signal \D_LM_040_in_0\ : std_logic;
signal \D_UU_040_in_0\ : std_logic;
signal \un1_D_UU_040_0\ : std_logic;
signal \D_LL_AMIGA_in_6\ : std_logic;
signal \un2_D_LL_AMIGA_6\ : std_logic;
signal \U111_CYCLE_SM.N_124_0\ : std_logic;
signal \U111_CYCLE_SM.N_132_cascade_\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNTZ0Z_1\ : std_logic;
signal \TBIn_c\ : std_logic;
signal \U111_CYCLE_SM.un7_CYCLE_STATE_0\ : std_logic;
signal \U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\ : std_logic;
signal \U111_CYCLE_SM.PORT_MISMATCHZ0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNTZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.BURSTZ0\ : std_logic;
signal \U111_CYCLE_SM.N_131_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0\ : std_logic;
signal \U111_CYCLE_SM.TS_EN6\ : std_logic;
signal \U111_CYCLE_SM.N_144\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\ : std_logic;
signal \D_UU_AMIGA_in_1\ : std_logic;
signal \un1_D_UU_AMIGA_1\ : std_logic;
signal \D_UM_040_in_3\ : std_logic;
signal \D_LL_040_in_3\ : std_logic;
signal \un1_D_UM_040_3\ : std_logic;
signal \D_LM_040_in_3\ : std_logic;
signal \D_UU_040_in_3\ : std_logic;
signal \un1_D_UU_040_3\ : std_logic;
signal \LBENn_c_i_0\ : std_logic;
signal \D_LL_AMIGA_in_7\ : std_logic;
signal \un2_D_LL_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.N_119_0\ : std_logic;
signal \U111_CYCLE_SM.N_117_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_cascade_\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1_cascade_\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \TEAn_c\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\ : std_logic;
signal \U111_CYCLE_SM.TA_DISZ0\ : std_logic;
signal \TAn_1_i\ : std_logic;
signal \D_LM_AMIGA_in_4\ : std_logic;
signal \un2_D_LM_AMIGA_4\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\ : std_logic;
signal \D_UU_AMIGA_in_5\ : std_logic;
signal \un1_D_UU_AMIGA_5\ : std_logic;
signal \D_UM_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\ : std_logic;
signal \un1_D_UM_AMIGA_1\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\ : std_logic;
signal \D_UU_AMIGA_in_0\ : std_logic;
signal \un1_D_UU_AMIGA_0\ : std_logic;
signal \D_LL_AMIGA_in_5\ : std_logic;
signal \un2_D_LL_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1\ : std_logic;
signal \CLK80\ : std_logic;
signal \GB_BUFFER_CLK80_THRU_CO\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\ : std_logic;
signal \D_UU_AMIGA_in_2\ : std_logic;
signal \un1_D_UU_AMIGA_2\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\ : std_logic;
signal \un1_D_UU_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\ : std_logic;
signal \D_UU_AMIGA_in_4\ : std_logic;
signal \un1_D_UU_AMIGA_4\ : std_logic;
signal \D_UM_AMIGA_in_3\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\ : std_logic;
signal \un1_D_UM_AMIGA_3\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\ : std_logic;
signal \D_UM_AMIGA_in_4\ : std_logic;
signal \un1_D_UM_AMIGA_4\ : std_logic;
signal \D_LM_AMIGA_in_7\ : std_logic;
signal \D_UU_AMIGA_in_7\ : std_logic;
signal \un2_D_LM_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\ : std_logic;
signal \D_UM_AMIGA_in_7\ : std_logic;
signal \un1_D_UM_AMIGA_7\ : std_logic;
signal \D_UM_AMIGA_in_5\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\ : std_logic;
signal \un1_D_UM_AMIGA_5\ : std_logic;
signal \D_UU_040_in_2\ : std_logic;
signal \D_LM_040_in_2\ : std_logic;
signal \un1_D_UU_040_2\ : std_logic;
signal \D_UU_040_in_5\ : std_logic;
signal \D_LM_040_in_5\ : std_logic;
signal \un1_D_UU_040_5\ : std_logic;
signal \D_UU_AMIGA_in_3\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\ : std_logic;
signal \un1_D_UU_AMIGA_3\ : std_logic;
signal \D_UU_AMIGA_in_6\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\ : std_logic;
signal \un1_D_UU_AMIGA_6\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\ : std_logic;
signal \D_UM_AMIGA_in_2\ : std_logic;
signal \un1_D_UM_AMIGA_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\ : std_logic;
signal \D_UM_AMIGA_in_6\ : std_logic;
signal \un1_D_UM_AMIGA_6\ : std_logic;
signal \D_LL_040_in_4\ : std_logic;
signal \D_UM_040_in_4\ : std_logic;
signal \un1_D_UM_040_4\ : std_logic;
signal \D_UU_040_in_4\ : std_logic;
signal \D_LM_040_in_4\ : std_logic;
signal \un1_D_UU_040_4\ : std_logic;
signal \U111_CYCLE_SM.LATCH_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\ : std_logic;
signal \D_UM_AMIGA_in_0\ : std_logic;
signal \un1_D_UM_AMIGA_0\ : std_logic;
signal \D_UM_040_in_7\ : std_logic;
signal \D_LL_040_in_7\ : std_logic;
signal \un1_D_UM_040_7\ : std_logic;
signal \U111_CYCLE_SM.FLIP_WORDZ0\ : std_logic;
signal \D_UU_040_in_7\ : std_logic;
signal \D_LM_040_in_7\ : std_logic;
signal \un1_D_UU_040_7\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep4_i_ess\ : std_logic;
signal \N_185_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep2_i_ess\ : std_logic;
signal \N_183_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep0_i_ess\ : std_logic;
signal \N_181_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep7_i_ess\ : std_logic;
signal \N_188_i\ : std_logic;
signal \N_209_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep28_i_ess\ : std_logic;
signal \GB_BUFFER_CLK40_THRU_CO\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep5_i_ess\ : std_logic;
signal \N_186_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep6_i_ess\ : std_logic;
signal \N_187_i\ : std_logic;
signal \N_193_i\ : std_logic;
signal \N_194_i\ : std_logic;
signal \N_205_i\ : std_logic;
signal \N_206_i\ : std_logic;
signal \N_208_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep25_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep24_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep27_i_ess\ : std_logic;
signal \N_211_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep26_i_ess\ : std_logic;
signal \N_207_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep30_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep17_i_ess\ : std_logic;
signal \N_198_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep18_i_ess\ : std_logic;
signal \N_199_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep31_i_ess\ : std_logic;
signal \N_212_i\ : std_logic;
signal \N_197_i\ : std_logic;
signal \N_200_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep19_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep16_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep20_i_ess\ : std_logic;
signal \N_201_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep8_i_ess\ : std_logic;
signal \N_189_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep21_i_ess\ : std_logic;
signal \N_202_i\ : std_logic;
signal \N_210_i\ : std_logic;
signal \N_191_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep10_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep29_i_ess\ : std_logic;
signal \N_195_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep14_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep22_i_ess\ : std_logic;
signal \N_203_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep23_i_ess\ : std_logic;
signal \N_204_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep9_i_ess\ : std_logic;
signal \N_190_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep11_i_ess\ : std_logic;
signal \N_192_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep3_i_ess\ : std_logic;
signal \N_184_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep15_i_ess\ : std_logic;
signal \N_196_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep1_i_ess\ : std_logic;
signal \N_182_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep13_i_ess\ : std_logic;
signal \BGn_c\ : std_logic;
signal \TS_CPUn_c\ : std_logic;
signal \LBENn_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep12_i_ess\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK40\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_g_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \LBENn_wire\ : std_logic;
signal \CPUBGn_wire\ : std_logic;
signal \A_040_wire\ : std_logic_vector(1 downto 0);
signal \CLK40B_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \BUFDIR_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \TS_CPUn_wire\ : std_logic;
signal \CLKRAMB_wire\ : std_logic;
signal \TEAn_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \DMAn_wire\ : std_logic;
signal \CLK80_CPU_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \A_AMIGA_wire\ : std_logic_vector(1 downto 0);
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \BGn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \TBI_CPUn_wire\ : std_logic;
signal \CLK40A_wire\ : std_logic;
signal \CLKRAMA_wire\ : std_logic;
signal \TCI_CPUn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \TEA_CPUn_wire\ : std_logic;
signal \pll_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \LBENn_wire\ <= LBENn;
    CPUBGn <= \CPUBGn_wire\;
    \A_040_wire\ <= A_040;
    CLK40B <= \CLK40B_wire\;
    \TBIn_wire\ <= TBIn;
    BUFDIR <= \BUFDIR_wire\;
    \SIZ_wire\ <= SIZ;
    \TS_CPUn_wire\ <= TS_CPUn;
    CLKRAMB <= \CLKRAMB_wire\;
    \TEAn_wire\ <= TEAn;
    BUFENn <= \BUFENn_wire\;
    DMAn <= \DMAn_wire\;
    CLK80_CPU <= \CLK80_CPU_wire\;
    TSn <= \TSn_wire\;
    \PORTSIZE_wire\ <= PORTSIZE;
    A_AMIGA <= \A_AMIGA_wire\;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    \BGn_wire\ <= BGn;
    \TCIn_wire\ <= TCIn;
    TBI_CPUn <= \TBI_CPUn_wire\;
    CLK40A <= \CLK40A_wire\;
    CLKRAMA <= \CLKRAMA_wire\;
    TCI_CPUn <= \TCI_CPUn_wire\;
    \RnW_wire\ <= RnW;
    TEA_CPUn <= \TEA_CPUn_wire\;
    \pll_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_pll\ : PLL40_2F
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            SCLK => '0',
            PLLOUTGLOBALA => \CLK80\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALB => \CLK40\,
            SDI => '0',
            PLLOUTCOREA => OPEN,
            BYPASS => '0',
            RESETB => \N__5708\,
            PLLOUTCOREB => OPEN,
            LOCK => OPEN,
            SDO => OPEN,
            EXTFEEDBACK => '0',
            DYNAMICDELAY => \pll_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__13729\
        );

    \pll_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__13729\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \LBENn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13713\,
            DIN => \N__13712\,
            DOUT => \N__13711\,
            PACKAGEPIN => \LBENn_wire\
        );

    \LBENn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13713\,
            PADOUT => \N__13712\,
            PADIN => \N__13711\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \LBENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13704\,
            DIN => \N__13703\,
            DOUT => \N__13702\,
            PACKAGEPIN => TAn
        );

    \TAn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13704\,
            PADOUT => \N__13703\,
            PADIN => \N__13702\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7106\,
            DIN0 => \TAn_in\,
            DOUT0 => \N__7418\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13695\,
            DIN => \N__13694\,
            DOUT => \N__13693\,
            PACKAGEPIN => D_LL_AMIGA(1)
        );

    \D_LL_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13695\,
            PADOUT => \N__13694\,
            PADIN => \N__13693\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4103\,
            DIN0 => \D_LL_AMIGA_in_1\,
            DOUT0 => \N__5561\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13686\,
            DIN => \N__13685\,
            DOUT => \N__13684\,
            PACKAGEPIN => D_UU_040(6)
        );

    \D_UU_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13686\,
            PADOUT => \N__13685\,
            PADIN => \N__13684\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9524\,
            DIN0 => \D_UU_040_in_6\,
            DOUT0 => \N__7886\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUBGn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13677\,
            DIN => \N__13676\,
            DOUT => \N__13675\,
            PACKAGEPIN => \CPUBGn_wire\
        );

    \CPUBGn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13677\,
            PADOUT => \N__13676\,
            PADIN => \N__13675\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13668\,
            DIN => \N__13667\,
            DOUT => \N__13666\,
            PACKAGEPIN => D_UM_AMIGA(3)
        );

    \D_UM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13668\,
            PADOUT => \N__13667\,
            PADIN => \N__13666\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4310\,
            DIN0 => \D_UM_AMIGA_in_3\,
            DOUT0 => \N__6401\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13659\,
            DIN => \N__13658\,
            DOUT => \N__13657\,
            PACKAGEPIN => \A_040_wire\(1)
        );

    \A_040_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13659\,
            PADOUT => \N__13658\,
            PADIN => \N__13657\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13650\,
            DIN => \N__13649\,
            DOUT => \N__13648\,
            PACKAGEPIN => D_LM_AMIGA(4)
        );

    \D_LM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13650\,
            PADOUT => \N__13649\,
            PADIN => \N__13648\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4394\,
            DIN0 => \D_LM_AMIGA_in_4\,
            DOUT0 => \N__9164\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13641\,
            DIN => \N__13640\,
            DOUT => \N__13639\,
            PACKAGEPIN => D_LM_040(7)
        );

    \D_LM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13641\,
            PADOUT => \N__13640\,
            PADIN => \N__13639\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9971\,
            DIN0 => \D_LM_040_in_7\,
            DOUT0 => \N__8339\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13632\,
            DIN => \N__13631\,
            DOUT => \N__13630\,
            PACKAGEPIN => \CLK40B_wire\
        );

    \CLK40B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13632\,
            PADOUT => \N__13631\,
            PADIN => \N__13630\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9617\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13623\,
            DIN => \N__13622\,
            DOUT => \N__13621\,
            PACKAGEPIN => D_UM_040(1)
        );

    \D_UM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13623\,
            PADOUT => \N__13622\,
            PADIN => \N__13621\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9950\,
            DIN0 => \D_UM_040_in_1\,
            DOUT0 => \N__6917\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13614\,
            DIN => \N__13613\,
            DOUT => \N__13612\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13614\,
            PADOUT => \N__13613\,
            PADIN => \N__13612\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TBIn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13605\,
            DIN => \N__13604\,
            DOUT => \N__13603\,
            PACKAGEPIN => D_UU_AMIGA(7)
        );

    \D_UU_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13605\,
            PADOUT => \N__13604\,
            PADIN => \N__13603\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4847\,
            DIN0 => \D_UU_AMIGA_in_7\,
            DOUT0 => \N__8498\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13596\,
            DIN => \N__13595\,
            DOUT => \N__13594\,
            PACKAGEPIN => \BUFDIR_wire\
        );

    \BUFDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13596\,
            PADOUT => \N__13595\,
            PADIN => \N__13594\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10580\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13587\,
            DIN => \N__13586\,
            DOUT => \N__13585\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13587\,
            PADOUT => \N__13586\,
            PADIN => \N__13585\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TS_CPUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13578\,
            DIN => \N__13577\,
            DOUT => \N__13576\,
            PACKAGEPIN => \TS_CPUn_wire\
        );

    \TS_CPUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13578\,
            PADOUT => \N__13577\,
            PADIN => \N__13576\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TS_CPUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13569\,
            DIN => \N__13568\,
            DOUT => \N__13567\,
            PACKAGEPIN => D_LL_040(1)
        );

    \D_LL_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13569\,
            PADOUT => \N__13568\,
            PADIN => \N__13567\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9680\,
            DIN0 => \D_LL_040_in_1\,
            DOUT0 => \N__4922\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13560\,
            DIN => \N__13559\,
            DOUT => \N__13558\,
            PACKAGEPIN => D_UU_040(1)
        );

    \D_UU_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13560\,
            PADOUT => \N__13559\,
            PADIN => \N__13558\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__12278\,
            DIN0 => \D_UU_040_in_1\,
            DOUT0 => \N__6482\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13551\,
            DIN => \N__13550\,
            DOUT => \N__13549\,
            PACKAGEPIN => D_LM_AMIGA(1)
        );

    \D_LM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13551\,
            PADOUT => \N__13550\,
            PADIN => \N__13549\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4226\,
            DIN0 => \D_LM_AMIGA_in_1\,
            DOUT0 => \N__5465\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13542\,
            DIN => \N__13541\,
            DOUT => \N__13540\,
            PACKAGEPIN => D_LM_040(2)
        );

    \D_LM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13542\,
            PADOUT => \N__13541\,
            PADIN => \N__13540\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9791\,
            DIN0 => \D_LM_040_in_2\,
            DOUT0 => \N__5000\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13533\,
            DIN => \N__13532\,
            DOUT => \N__13531\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13533\,
            PADOUT => \N__13532\,
            PADIN => \N__13531\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6818\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__4178\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13524\,
            DIN => \N__13523\,
            DOUT => \N__13522\,
            PACKAGEPIN => D_UM_040(2)
        );

    \D_UM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13524\,
            PADOUT => \N__13523\,
            PADIN => \N__13522\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9860\,
            DIN0 => \D_UM_040_in_2\,
            DOUT0 => \N__9350\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13515\,
            DIN => \N__13514\,
            DOUT => \N__13513\,
            PACKAGEPIN => \CLKRAMB_wire\
        );

    \CLKRAMB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13515\,
            PADOUT => \N__13514\,
            PADIN => \N__13513\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7751\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13506\,
            DIN => \N__13505\,
            DOUT => \N__13504\,
            PACKAGEPIN => D_LL_AMIGA(2)
        );

    \D_LL_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13506\,
            PADOUT => \N__13505\,
            PADIN => \N__13504\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4124\,
            DIN0 => \D_LL_AMIGA_in_2\,
            DOUT0 => \N__4730\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13497\,
            DIN => \N__13496\,
            DOUT => \N__13495\,
            PACKAGEPIN => D_UU_AMIGA(2)
        );

    \D_UU_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13497\,
            PADOUT => \N__13496\,
            PADIN => \N__13495\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5099\,
            DIN0 => \D_UU_AMIGA_in_2\,
            DOUT0 => \N__8117\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEAn_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13488\,
            DIN => \N__13487\,
            DOUT => \N__13486\,
            PACKAGEPIN => \TEAn_wire\
        );

    \TEAn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13488\,
            PADOUT => \N__13487\,
            PADIN => \N__13486\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TEAn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13479\,
            DIN => \N__13478\,
            DOUT => \N__13477\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13479\,
            PADOUT => \N__13478\,
            PADIN => \N__13477\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5123\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMAn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13470\,
            DIN => \N__13469\,
            DOUT => \N__13468\,
            PACKAGEPIN => \DMAn_wire\
        );

    \DMAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13470\,
            PADOUT => \N__13469\,
            PADIN => \N__13468\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5707\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13461\,
            DIN => \N__13460\,
            DOUT => \N__13459\,
            PACKAGEPIN => D_LL_040(6)
        );

    \D_LL_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13461\,
            PADOUT => \N__13460\,
            PADIN => \N__13459\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9632\,
            DIN0 => \D_LL_040_in_6\,
            DOUT0 => \N__5864\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13452\,
            DIN => \N__13451\,
            DOUT => \N__13450\,
            PACKAGEPIN => D_LL_AMIGA(5)
        );

    \D_LL_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13452\,
            PADOUT => \N__13451\,
            PADIN => \N__13450\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4079\,
            DIN0 => \D_LL_AMIGA_in_5\,
            DOUT0 => \N__5396\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13443\,
            DIN => \N__13442\,
            DOUT => \N__13441\,
            PACKAGEPIN => D_UM_AMIGA(0)
        );

    \D_UM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13443\,
            PADOUT => \N__13442\,
            PADIN => \N__13441\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4187\,
            DIN0 => \D_UM_AMIGA_in_0\,
            DOUT0 => \N__5180\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13434\,
            DIN => \N__13433\,
            DOUT => \N__13432\,
            PACKAGEPIN => D_UU_040(2)
        );

    \D_UU_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13434\,
            PADOUT => \N__13433\,
            PADIN => \N__13432\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9482\,
            DIN0 => \D_UU_040_in_2\,
            DOUT0 => \N__7661\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13425\,
            DIN => \N__13424\,
            DOUT => \N__13423\,
            PACKAGEPIN => D_LM_AMIGA(2)
        );

    \D_LM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13425\,
            PADOUT => \N__13424\,
            PADIN => \N__13423\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4565\,
            DIN0 => \D_LM_AMIGA_in_2\,
            DOUT0 => \N__8155\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK80_CPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13416\,
            DIN => \N__13415\,
            DOUT => \N__13414\,
            PACKAGEPIN => \CLK80_CPU_wire\
        );

    \CLK80_CPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13416\,
            PADOUT => \N__13415\,
            PADIN => \N__13414\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7750\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13407\,
            DIN => \N__13406\,
            DOUT => \N__13405\,
            PACKAGEPIN => D_LL_040(3)
        );

    \D_LL_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13407\,
            PADOUT => \N__13406\,
            PADIN => \N__13405\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9665\,
            DIN0 => \D_LL_040_in_3\,
            DOUT0 => \N__5747\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13398\,
            DIN => \N__13397\,
            DOUT => \N__13396\,
            PACKAGEPIN => D_LM_040(1)
        );

    \D_LM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13398\,
            PADOUT => \N__13397\,
            PADIN => \N__13396\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9812\,
            DIN0 => \D_LM_040_in_1\,
            DOUT0 => \N__4769\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13389\,
            DIN => \N__13388\,
            DOUT => \N__13387\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13389\,
            PADOUT => \N__13388\,
            PADIN => \N__13387\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5606\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13380\,
            DIN => \N__13379\,
            DOUT => \N__13378\,
            PACKAGEPIN => D_UM_AMIGA(7)
        );

    \D_UM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13380\,
            PADOUT => \N__13379\,
            PADIN => \N__13378\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4484\,
            DIN0 => \D_UM_AMIGA_in_7\,
            DOUT0 => \N__8843\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13371\,
            DIN => \N__13370\,
            DOUT => \N__13369\,
            PACKAGEPIN => D_LM_AMIGA(7)
        );

    \D_LM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13371\,
            PADOUT => \N__13370\,
            PADIN => \N__13369\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4340\,
            DIN0 => \D_LM_AMIGA_in_7\,
            DOUT0 => \N__8537\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13362\,
            DIN => \N__13361\,
            DOUT => \N__13360\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13362\,
            PADOUT => \N__13361\,
            PADIN => \N__13360\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PORTSIZE_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13353\,
            DIN => \N__13352\,
            DOUT => \N__13351\,
            PACKAGEPIN => \A_AMIGA_wire\(0)
        );

    \A_AMIGA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13353\,
            PADOUT => \N__13352\,
            PADIN => \N__13351\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4613\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13344\,
            DIN => \N__13343\,
            DOUT => \N__13342\,
            PACKAGEPIN => D_LM_040(4)
        );

    \D_LM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13344\,
            PADOUT => \N__13343\,
            PADIN => \N__13342\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9923\,
            DIN0 => \D_LM_040_in_4\,
            DOUT0 => \N__7067\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13335\,
            DIN => \N__13334\,
            DOUT => \N__13333\,
            PACKAGEPIN => D_UM_040(7)
        );

    \D_UM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13335\,
            PADOUT => \N__13334\,
            PADIN => \N__13333\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__12299\,
            DIN0 => \D_UM_040_in_7\,
            DOUT0 => \N__8276\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13326\,
            DIN => \N__13325\,
            DOUT => \N__13324\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13326\,
            PADOUT => \N__13325\,
            PADIN => \N__13324\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13317\,
            DIN => \N__13316\,
            DOUT => \N__13315\,
            PACKAGEPIN => D_UU_AMIGA(1)
        );

    \D_UU_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13317\,
            PADOUT => \N__13316\,
            PADIN => \N__13315\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4499\,
            DIN0 => \D_UU_AMIGA_in_1\,
            DOUT0 => \N__5414\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13308\,
            DIN => \N__13307\,
            DOUT => \N__13306\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13308\,
            PADOUT => \N__13307\,
            PADIN => \N__13306\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9616\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13299\,
            DIN => \N__13298\,
            DOUT => \N__13297\,
            PACKAGEPIN => D_UM_040(0)
        );

    \D_UM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13299\,
            PADOUT => \N__13298\,
            PADIN => \N__13297\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9905\,
            DIN0 => \D_UM_040_in_0\,
            DOUT0 => \N__8927\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13290\,
            DIN => \N__13289\,
            DOUT => \N__13288\,
            PACKAGEPIN => D_LL_AMIGA(0)
        );

    \D_LL_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13290\,
            PADOUT => \N__13289\,
            PADIN => \N__13288\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4139\,
            DIN0 => \D_LL_AMIGA_in_0\,
            DOUT0 => \N__5240\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13281\,
            DIN => \N__13280\,
            DOUT => \N__13279\,
            PACKAGEPIN => D_UU_AMIGA(4)
        );

    \D_UU_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13281\,
            PADOUT => \N__13280\,
            PADIN => \N__13279\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5291\,
            DIN0 => \D_UU_AMIGA_in_4\,
            DOUT0 => \N__9128\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13272\,
            DIN => \N__13271\,
            DOUT => \N__13270\,
            PACKAGEPIN => D_UU_040(7)
        );

    \D_UU_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13272\,
            PADOUT => \N__13271\,
            PADIN => \N__13270\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9437\,
            DIN0 => \D_UU_040_in_7\,
            DOUT0 => \N__7631\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13263\,
            DIN => \N__13262\,
            DOUT => \N__13261\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13263\,
            PADOUT => \N__13262\,
            PADIN => \N__13261\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BGn_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13254\,
            DIN => \N__13253\,
            DOUT => \N__13252\,
            PACKAGEPIN => \BGn_wire\
        );

    \BGn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13254\,
            PADOUT => \N__13253\,
            PADIN => \N__13252\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BGn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13245\,
            DIN => \N__13244\,
            DOUT => \N__13243\,
            PACKAGEPIN => D_LL_040(0)
        );

    \D_LL_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13245\,
            PADOUT => \N__13244\,
            PADIN => \N__13243\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9695\,
            DIN0 => \D_LL_040_in_0\,
            DOUT0 => \N__4793\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13236\,
            DIN => \N__13235\,
            DOUT => \N__13234\,
            PACKAGEPIN => D_UM_AMIGA(2)
        );

    \D_UM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13236\,
            PADOUT => \N__13235\,
            PADIN => \N__13234\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4406\,
            DIN0 => \D_UM_AMIGA_in_2\,
            DOUT0 => \N__4685\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13227\,
            DIN => \N__13226\,
            DOUT => \N__13225\,
            PACKAGEPIN => D_UU_040(0)
        );

    \D_UU_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13227\,
            PADOUT => \N__13226\,
            PADIN => \N__13225\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9461\,
            DIN0 => \D_UU_040_in_0\,
            DOUT0 => \N__6839\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13218\,
            DIN => \N__13217\,
            DOUT => \N__13216\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13218\,
            PADOUT => \N__13217\,
            PADIN => \N__13216\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TCIn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13209\,
            DIN => \N__13208\,
            DOUT => \N__13207\,
            PACKAGEPIN => \A_040_wire\(0)
        );

    \A_040_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13209\,
            PADOUT => \N__13208\,
            PADIN => \N__13207\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13200\,
            DIN => \N__13199\,
            DOUT => \N__13198\,
            PACKAGEPIN => D_LM_AMIGA(0)
        );

    \D_LM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13200\,
            PADOUT => \N__13199\,
            PADIN => \N__13198\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4268\,
            DIN0 => \D_LM_AMIGA_in_0\,
            DOUT0 => \N__5963\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13191\,
            DIN => \N__13190\,
            DOUT => \N__13189\,
            PACKAGEPIN => \TBI_CPUn_wire\
        );

    \TBI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13191\,
            PADOUT => \N__13190\,
            PADIN => \N__13189\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6274\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13182\,
            DIN => \N__13181\,
            DOUT => \N__13180\,
            PACKAGEPIN => \CLK40A_wire\
        );

    \CLK40A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13182\,
            PADOUT => \N__13181\,
            PADIN => \N__13180\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9596\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13173\,
            DIN => \N__13172\,
            DOUT => \N__13171\,
            PACKAGEPIN => D_LM_040(3)
        );

    \D_LM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13173\,
            PADOUT => \N__13172\,
            PADIN => \N__13171\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9743\,
            DIN0 => \D_LM_040_in_3\,
            DOUT0 => \N__5147\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13164\,
            DIN => \N__13163\,
            DOUT => \N__13162\,
            PACKAGEPIN => D_LM_AMIGA(5)
        );

    \D_LM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13164\,
            PADOUT => \N__13163\,
            PADIN => \N__13162\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4373\,
            DIN0 => \D_LM_AMIGA_in_5\,
            DOUT0 => \N__8075\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13155\,
            DIN => \N__13154\,
            DOUT => \N__13153\,
            PACKAGEPIN => D_LM_040(6)
        );

    \D_LM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13155\,
            PADOUT => \N__13154\,
            PADIN => \N__13153\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9992\,
            DIN0 => \D_LM_040_in_6\,
            DOUT0 => \N__5483\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13146\,
            DIN => \N__13145\,
            DOUT => \N__13144\,
            PACKAGEPIN => D_UM_040(5)
        );

    \D_UM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13146\,
            PADOUT => \N__13145\,
            PADIN => \N__13144\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9710\,
            DIN0 => \D_UM_040_in_5\,
            DOUT0 => \N__8201\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13137\,
            DIN => \N__13136\,
            DOUT => \N__13135\,
            PACKAGEPIN => D_LL_AMIGA(3)
        );

    \D_LL_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13137\,
            PADOUT => \N__13136\,
            PADIN => \N__13135\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4154\,
            DIN0 => \D_LL_AMIGA_in_3\,
            DOUT0 => \N__6445\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13128\,
            DIN => \N__13127\,
            DOUT => \N__13126\,
            PACKAGEPIN => D_UU_AMIGA(3)
        );

    \D_UU_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13128\,
            PADOUT => \N__13127\,
            PADIN => \N__13126\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4667\,
            DIN0 => \D_UU_AMIGA_in_3\,
            DOUT0 => \N__6323\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13119\,
            DIN => \N__13118\,
            DOUT => \N__13117\,
            PACKAGEPIN => D_LL_040(5)
        );

    \D_LL_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13119\,
            PADOUT => \N__13118\,
            PADIN => \N__13117\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9875\,
            DIN0 => \D_LL_040_in_5\,
            DOUT0 => \N__7439\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13110\,
            DIN => \N__13109\,
            DOUT => \N__13108\,
            PACKAGEPIN => D_LL_AMIGA(6)
        );

    \D_LL_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13110\,
            PADOUT => \N__13109\,
            PADIN => \N__13108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4283\,
            DIN0 => \D_LL_AMIGA_in_6\,
            DOUT0 => \N__5063\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13101\,
            DIN => \N__13100\,
            DOUT => \N__13099\,
            PACKAGEPIN => D_UU_AMIGA(6)
        );

    \D_UU_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13101\,
            PADOUT => \N__13100\,
            PADIN => \N__13099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4823\,
            DIN0 => \D_UU_AMIGA_in_6\,
            DOUT0 => \N__5780\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13092\,
            DIN => \N__13091\,
            DOUT => \N__13090\,
            PACKAGEPIN => D_UM_AMIGA(1)
        );

    \D_UM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13092\,
            PADOUT => \N__13091\,
            PADIN => \N__13090\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4355\,
            DIN0 => \D_UM_AMIGA_in_1\,
            DOUT0 => \N__5519\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13083\,
            DIN => \N__13082\,
            DOUT => \N__13081\,
            PACKAGEPIN => D_UU_040(5)
        );

    \D_UU_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13083\,
            PADOUT => \N__13082\,
            PADIN => \N__13081\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9545\,
            DIN0 => \D_UU_040_in_5\,
            DOUT0 => \N__6989\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13074\,
            DIN => \N__13073\,
            DOUT => \N__13072\,
            PACKAGEPIN => \CLKRAMA_wire\
        );

    \CLKRAMA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13074\,
            PADOUT => \N__13073\,
            PADIN => \N__13072\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9606\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13065\,
            DIN => \N__13064\,
            DOUT => \N__13063\,
            PACKAGEPIN => D_LL_040(2)
        );

    \D_LL_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13065\,
            PADOUT => \N__13064\,
            PADIN => \N__13063\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9839\,
            DIN0 => \D_LL_040_in_2\,
            DOUT0 => \N__5669\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13056\,
            DIN => \N__13055\,
            DOUT => \N__13054\,
            PACKAGEPIN => \TCI_CPUn_wire\
        );

    \TCI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13056\,
            PADOUT => \N__13055\,
            PADIN => \N__13054\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4064\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13047\,
            DIN => \N__13046\,
            DOUT => \N__13045\,
            PACKAGEPIN => D_UM_AMIGA(4)
        );

    \D_UM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13047\,
            PADOUT => \N__13046\,
            PADIN => \N__13045\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4469\,
            DIN0 => \D_UM_AMIGA_in_4\,
            DOUT0 => \N__9206\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13038\,
            DIN => \N__13037\,
            DOUT => \N__13036\,
            PACKAGEPIN => D_LM_AMIGA(6)
        );

    \D_LM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13038\,
            PADOUT => \N__13037\,
            PADIN => \N__13036\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4325\,
            DIN0 => \D_LM_AMIGA_in_6\,
            DOUT0 => \N__5819\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13029\,
            DIN => \N__13028\,
            DOUT => \N__13027\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13029\,
            PADOUT => \N__13028\,
            PADIN => \N__13027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13020\,
            DIN => \N__13019\,
            DOUT => \N__13018\,
            PACKAGEPIN => D_LM_040(5)
        );

    \D_LM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13020\,
            PADOUT => \N__13019\,
            PADIN => \N__13018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9890\,
            DIN0 => \D_LM_040_in_5\,
            DOUT0 => \N__5984\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13011\,
            DIN => \N__13010\,
            DOUT => \N__13009\,
            PACKAGEPIN => D_UM_040(6)
        );

    \D_UM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13011\,
            PADOUT => \N__13010\,
            PADIN => \N__13009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10016\,
            DIN0 => \D_UM_040_in_6\,
            DOUT0 => \N__9287\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13002\,
            DIN => \N__13001\,
            DOUT => \N__13000\,
            PACKAGEPIN => D_UM_040(3)
        );

    \D_UM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13002\,
            PADOUT => \N__13001\,
            PADIN => \N__13000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__12344\,
            DIN0 => \D_UM_040_in_3\,
            DOUT0 => \N__7478\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12993\,
            DIN => \N__12992\,
            DOUT => \N__12991\,
            PACKAGEPIN => D_UU_AMIGA(5)
        );

    \D_UU_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12993\,
            PADOUT => \N__12992\,
            PADIN => \N__12991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4643\,
            DIN0 => \D_UU_AMIGA_in_5\,
            DOUT0 => \N__8027\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12984\,
            DIN => \N__12983\,
            DOUT => \N__12982\,
            PACKAGEPIN => D_LL_040(7)
        );

    \D_LL_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12984\,
            PADOUT => \N__12983\,
            PADIN => \N__12982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9773\,
            DIN0 => \D_LL_040_in_7\,
            DOUT0 => \N__6791\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12975\,
            DIN => \N__12974\,
            DOUT => \N__12973\,
            PACKAGEPIN => D_LL_AMIGA(4)
        );

    \D_LL_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12975\,
            PADOUT => \N__12974\,
            PADIN => \N__12973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4448\,
            DIN0 => \D_LL_AMIGA_in_4\,
            DOUT0 => \N__9269\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12966\,
            DIN => \N__12965\,
            DOUT => \N__12964\,
            PACKAGEPIN => D_UU_040(3)
        );

    \D_UU_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12966\,
            PADOUT => \N__12965\,
            PADIN => \N__12964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__12323\,
            DIN0 => \D_UU_040_in_3\,
            DOUT0 => \N__7949\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEA_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12957\,
            DIN => \N__12956\,
            DOUT => \N__12955\,
            PACKAGEPIN => \TEA_CPUn_wire\
        );

    \TEA_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12957\,
            PADOUT => \N__12956\,
            PADIN => \N__12955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7340\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12948\,
            DIN => \N__12947\,
            DOUT => \N__12946\,
            PACKAGEPIN => D_LM_AMIGA(3)
        );

    \D_LM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12948\,
            PADOUT => \N__12947\,
            PADIN => \N__12946\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4550\,
            DIN0 => \D_LM_AMIGA_in_3\,
            DOUT0 => \N__6383\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12939\,
            DIN => \N__12938\,
            DOUT => \N__12937\,
            PACKAGEPIN => D_LM_040(0)
        );

    \D_LM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12939\,
            PADOUT => \N__12938\,
            PADIN => \N__12937\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9758\,
            DIN0 => \D_LM_040_in_0\,
            DOUT0 => \N__5630\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12930\,
            DIN => \N__12929\,
            DOUT => \N__12928\,
            PACKAGEPIN => D_UM_AMIGA(6)
        );

    \D_UM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12930\,
            PADOUT => \N__12929\,
            PADIN => \N__12928\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4295\,
            DIN0 => \D_UM_AMIGA_in_6\,
            DOUT0 => \N__5024\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__12921\,
            DIN => \N__12920\,
            DOUT => \N__12919\,
            PACKAGEPIN => \A_AMIGA_wire\(1)
        );

    \A_AMIGA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12921\,
            PADOUT => \N__12920\,
            PADIN => \N__12919\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4598\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12912\,
            DIN => \N__12911\,
            DOUT => \N__12910\,
            PACKAGEPIN => D_UM_040(4)
        );

    \D_UM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12912\,
            PADOUT => \N__12911\,
            PADIN => \N__12910\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9725\,
            DIN0 => \D_UM_040_in_4\,
            DOUT0 => \N__8414\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12903\,
            DIN => \N__12902\,
            DOUT => \N__12901\,
            PACKAGEPIN => D_UU_AMIGA(0)
        );

    \D_UU_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12903\,
            PADOUT => \N__12902\,
            PADIN => \N__12901\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4976\,
            DIN0 => \D_UU_AMIGA_in_0\,
            DOUT0 => \N__5894\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12894\,
            DIN => \N__12893\,
            DOUT => \N__12892\,
            PACKAGEPIN => D_LL_040(4)
        );

    \D_LL_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12894\,
            PADOUT => \N__12893\,
            PADIN => \N__12892\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9422\,
            DIN0 => \D_LL_040_in_4\,
            DOUT0 => \N__5261\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12885\,
            DIN => \N__12884\,
            DOUT => \N__12883\,
            PACKAGEPIN => D_LL_AMIGA(7)
        );

    \D_LL_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12885\,
            PADOUT => \N__12884\,
            PADIN => \N__12883\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4256\,
            DIN0 => \D_LL_AMIGA_in_7\,
            DOUT0 => \N__8894\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12876\,
            DIN => \N__12875\,
            DOUT => \N__12874\,
            PACKAGEPIN => D_UU_040(4)
        );

    \D_UU_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12876\,
            PADOUT => \N__12875\,
            PADIN => \N__12874\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9503\,
            DIN0 => \D_UU_040_in_4\,
            DOUT0 => \N__7562\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12867\,
            DIN => \N__12866\,
            DOUT => \N__12865\,
            PACKAGEPIN => D_UM_AMIGA(5)
        );

    \D_UM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12867\,
            PADOUT => \N__12866\,
            PADIN => \N__12865\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4961\,
            DIN0 => \D_UM_AMIGA_in_5\,
            DOUT0 => \N__5324\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3278\ : InMux
    port map (
            O => \N__12848\,
            I => \N__12845\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__12845\,
            I => \N__12828\
        );

    \I__3276\ : ClkMux
    port map (
            O => \N__12844\,
            I => \N__12659\
        );

    \I__3275\ : ClkMux
    port map (
            O => \N__12843\,
            I => \N__12659\
        );

    \I__3274\ : ClkMux
    port map (
            O => \N__12842\,
            I => \N__12659\
        );

    \I__3273\ : ClkMux
    port map (
            O => \N__12841\,
            I => \N__12659\
        );

    \I__3272\ : ClkMux
    port map (
            O => \N__12840\,
            I => \N__12659\
        );

    \I__3271\ : ClkMux
    port map (
            O => \N__12839\,
            I => \N__12659\
        );

    \I__3270\ : ClkMux
    port map (
            O => \N__12838\,
            I => \N__12659\
        );

    \I__3269\ : ClkMux
    port map (
            O => \N__12837\,
            I => \N__12659\
        );

    \I__3268\ : ClkMux
    port map (
            O => \N__12836\,
            I => \N__12659\
        );

    \I__3267\ : ClkMux
    port map (
            O => \N__12835\,
            I => \N__12659\
        );

    \I__3266\ : ClkMux
    port map (
            O => \N__12834\,
            I => \N__12659\
        );

    \I__3265\ : ClkMux
    port map (
            O => \N__12833\,
            I => \N__12659\
        );

    \I__3264\ : ClkMux
    port map (
            O => \N__12832\,
            I => \N__12659\
        );

    \I__3263\ : ClkMux
    port map (
            O => \N__12831\,
            I => \N__12659\
        );

    \I__3262\ : Glb2LocalMux
    port map (
            O => \N__12828\,
            I => \N__12659\
        );

    \I__3261\ : ClkMux
    port map (
            O => \N__12827\,
            I => \N__12659\
        );

    \I__3260\ : ClkMux
    port map (
            O => \N__12826\,
            I => \N__12659\
        );

    \I__3259\ : ClkMux
    port map (
            O => \N__12825\,
            I => \N__12659\
        );

    \I__3258\ : ClkMux
    port map (
            O => \N__12824\,
            I => \N__12659\
        );

    \I__3257\ : ClkMux
    port map (
            O => \N__12823\,
            I => \N__12659\
        );

    \I__3256\ : ClkMux
    port map (
            O => \N__12822\,
            I => \N__12659\
        );

    \I__3255\ : ClkMux
    port map (
            O => \N__12821\,
            I => \N__12659\
        );

    \I__3254\ : ClkMux
    port map (
            O => \N__12820\,
            I => \N__12659\
        );

    \I__3253\ : ClkMux
    port map (
            O => \N__12819\,
            I => \N__12659\
        );

    \I__3252\ : ClkMux
    port map (
            O => \N__12818\,
            I => \N__12659\
        );

    \I__3251\ : ClkMux
    port map (
            O => \N__12817\,
            I => \N__12659\
        );

    \I__3250\ : ClkMux
    port map (
            O => \N__12816\,
            I => \N__12659\
        );

    \I__3249\ : ClkMux
    port map (
            O => \N__12815\,
            I => \N__12659\
        );

    \I__3248\ : ClkMux
    port map (
            O => \N__12814\,
            I => \N__12659\
        );

    \I__3247\ : ClkMux
    port map (
            O => \N__12813\,
            I => \N__12659\
        );

    \I__3246\ : ClkMux
    port map (
            O => \N__12812\,
            I => \N__12659\
        );

    \I__3245\ : ClkMux
    port map (
            O => \N__12811\,
            I => \N__12659\
        );

    \I__3244\ : ClkMux
    port map (
            O => \N__12810\,
            I => \N__12659\
        );

    \I__3243\ : ClkMux
    port map (
            O => \N__12809\,
            I => \N__12659\
        );

    \I__3242\ : ClkMux
    port map (
            O => \N__12808\,
            I => \N__12659\
        );

    \I__3241\ : ClkMux
    port map (
            O => \N__12807\,
            I => \N__12659\
        );

    \I__3240\ : ClkMux
    port map (
            O => \N__12806\,
            I => \N__12659\
        );

    \I__3239\ : ClkMux
    port map (
            O => \N__12805\,
            I => \N__12659\
        );

    \I__3238\ : ClkMux
    port map (
            O => \N__12804\,
            I => \N__12659\
        );

    \I__3237\ : ClkMux
    port map (
            O => \N__12803\,
            I => \N__12659\
        );

    \I__3236\ : ClkMux
    port map (
            O => \N__12802\,
            I => \N__12659\
        );

    \I__3235\ : ClkMux
    port map (
            O => \N__12801\,
            I => \N__12659\
        );

    \I__3234\ : ClkMux
    port map (
            O => \N__12800\,
            I => \N__12659\
        );

    \I__3233\ : ClkMux
    port map (
            O => \N__12799\,
            I => \N__12659\
        );

    \I__3232\ : ClkMux
    port map (
            O => \N__12798\,
            I => \N__12659\
        );

    \I__3231\ : ClkMux
    port map (
            O => \N__12797\,
            I => \N__12659\
        );

    \I__3230\ : ClkMux
    port map (
            O => \N__12796\,
            I => \N__12659\
        );

    \I__3229\ : ClkMux
    port map (
            O => \N__12795\,
            I => \N__12659\
        );

    \I__3228\ : ClkMux
    port map (
            O => \N__12794\,
            I => \N__12659\
        );

    \I__3227\ : ClkMux
    port map (
            O => \N__12793\,
            I => \N__12659\
        );

    \I__3226\ : ClkMux
    port map (
            O => \N__12792\,
            I => \N__12659\
        );

    \I__3225\ : ClkMux
    port map (
            O => \N__12791\,
            I => \N__12659\
        );

    \I__3224\ : ClkMux
    port map (
            O => \N__12790\,
            I => \N__12659\
        );

    \I__3223\ : ClkMux
    port map (
            O => \N__12789\,
            I => \N__12659\
        );

    \I__3222\ : ClkMux
    port map (
            O => \N__12788\,
            I => \N__12659\
        );

    \I__3221\ : ClkMux
    port map (
            O => \N__12787\,
            I => \N__12659\
        );

    \I__3220\ : ClkMux
    port map (
            O => \N__12786\,
            I => \N__12659\
        );

    \I__3219\ : ClkMux
    port map (
            O => \N__12785\,
            I => \N__12659\
        );

    \I__3218\ : ClkMux
    port map (
            O => \N__12784\,
            I => \N__12659\
        );

    \I__3217\ : ClkMux
    port map (
            O => \N__12783\,
            I => \N__12659\
        );

    \I__3216\ : ClkMux
    port map (
            O => \N__12782\,
            I => \N__12659\
        );

    \I__3215\ : GlobalMux
    port map (
            O => \N__12659\,
            I => \CLK40\
        );

    \I__3214\ : CEMux
    port map (
            O => \N__12656\,
            I => \N__12521\
        );

    \I__3213\ : CEMux
    port map (
            O => \N__12655\,
            I => \N__12521\
        );

    \I__3212\ : CEMux
    port map (
            O => \N__12654\,
            I => \N__12521\
        );

    \I__3211\ : CEMux
    port map (
            O => \N__12653\,
            I => \N__12521\
        );

    \I__3210\ : CEMux
    port map (
            O => \N__12652\,
            I => \N__12521\
        );

    \I__3209\ : CEMux
    port map (
            O => \N__12651\,
            I => \N__12521\
        );

    \I__3208\ : CEMux
    port map (
            O => \N__12650\,
            I => \N__12521\
        );

    \I__3207\ : CEMux
    port map (
            O => \N__12649\,
            I => \N__12521\
        );

    \I__3206\ : CEMux
    port map (
            O => \N__12648\,
            I => \N__12521\
        );

    \I__3205\ : CEMux
    port map (
            O => \N__12647\,
            I => \N__12521\
        );

    \I__3204\ : CEMux
    port map (
            O => \N__12646\,
            I => \N__12521\
        );

    \I__3203\ : CEMux
    port map (
            O => \N__12645\,
            I => \N__12521\
        );

    \I__3202\ : CEMux
    port map (
            O => \N__12644\,
            I => \N__12521\
        );

    \I__3201\ : CEMux
    port map (
            O => \N__12643\,
            I => \N__12521\
        );

    \I__3200\ : CEMux
    port map (
            O => \N__12642\,
            I => \N__12521\
        );

    \I__3199\ : CEMux
    port map (
            O => \N__12641\,
            I => \N__12521\
        );

    \I__3198\ : CEMux
    port map (
            O => \N__12640\,
            I => \N__12521\
        );

    \I__3197\ : CEMux
    port map (
            O => \N__12639\,
            I => \N__12521\
        );

    \I__3196\ : CEMux
    port map (
            O => \N__12638\,
            I => \N__12521\
        );

    \I__3195\ : CEMux
    port map (
            O => \N__12637\,
            I => \N__12521\
        );

    \I__3194\ : CEMux
    port map (
            O => \N__12636\,
            I => \N__12521\
        );

    \I__3193\ : CEMux
    port map (
            O => \N__12635\,
            I => \N__12521\
        );

    \I__3192\ : CEMux
    port map (
            O => \N__12634\,
            I => \N__12521\
        );

    \I__3191\ : CEMux
    port map (
            O => \N__12633\,
            I => \N__12521\
        );

    \I__3190\ : CEMux
    port map (
            O => \N__12632\,
            I => \N__12521\
        );

    \I__3189\ : CEMux
    port map (
            O => \N__12631\,
            I => \N__12521\
        );

    \I__3188\ : CEMux
    port map (
            O => \N__12630\,
            I => \N__12521\
        );

    \I__3187\ : CEMux
    port map (
            O => \N__12629\,
            I => \N__12521\
        );

    \I__3186\ : CEMux
    port map (
            O => \N__12628\,
            I => \N__12521\
        );

    \I__3185\ : CEMux
    port map (
            O => \N__12627\,
            I => \N__12521\
        );

    \I__3184\ : CEMux
    port map (
            O => \N__12626\,
            I => \N__12521\
        );

    \I__3183\ : CEMux
    port map (
            O => \N__12625\,
            I => \N__12521\
        );

    \I__3182\ : CEMux
    port map (
            O => \N__12624\,
            I => \N__12521\
        );

    \I__3181\ : CEMux
    port map (
            O => \N__12623\,
            I => \N__12521\
        );

    \I__3180\ : CEMux
    port map (
            O => \N__12622\,
            I => \N__12521\
        );

    \I__3179\ : CEMux
    port map (
            O => \N__12621\,
            I => \N__12521\
        );

    \I__3178\ : CEMux
    port map (
            O => \N__12620\,
            I => \N__12521\
        );

    \I__3177\ : CEMux
    port map (
            O => \N__12619\,
            I => \N__12521\
        );

    \I__3176\ : CEMux
    port map (
            O => \N__12618\,
            I => \N__12521\
        );

    \I__3175\ : CEMux
    port map (
            O => \N__12617\,
            I => \N__12521\
        );

    \I__3174\ : CEMux
    port map (
            O => \N__12616\,
            I => \N__12521\
        );

    \I__3173\ : CEMux
    port map (
            O => \N__12615\,
            I => \N__12521\
        );

    \I__3172\ : CEMux
    port map (
            O => \N__12614\,
            I => \N__12521\
        );

    \I__3171\ : CEMux
    port map (
            O => \N__12613\,
            I => \N__12521\
        );

    \I__3170\ : CEMux
    port map (
            O => \N__12612\,
            I => \N__12521\
        );

    \I__3169\ : GlobalMux
    port map (
            O => \N__12521\,
            I => \N__12518\
        );

    \I__3168\ : gio2CtrlBuf
    port map (
            O => \N__12518\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_g_0\
        );

    \I__3167\ : InMux
    port map (
            O => \N__12515\,
            I => \N__12512\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__12512\,
            I => \N__12459\
        );

    \I__3165\ : SRMux
    port map (
            O => \N__12511\,
            I => \N__12356\
        );

    \I__3164\ : SRMux
    port map (
            O => \N__12510\,
            I => \N__12356\
        );

    \I__3163\ : SRMux
    port map (
            O => \N__12509\,
            I => \N__12356\
        );

    \I__3162\ : SRMux
    port map (
            O => \N__12508\,
            I => \N__12356\
        );

    \I__3161\ : SRMux
    port map (
            O => \N__12507\,
            I => \N__12356\
        );

    \I__3160\ : SRMux
    port map (
            O => \N__12506\,
            I => \N__12356\
        );

    \I__3159\ : SRMux
    port map (
            O => \N__12505\,
            I => \N__12356\
        );

    \I__3158\ : SRMux
    port map (
            O => \N__12504\,
            I => \N__12356\
        );

    \I__3157\ : SRMux
    port map (
            O => \N__12503\,
            I => \N__12356\
        );

    \I__3156\ : SRMux
    port map (
            O => \N__12502\,
            I => \N__12356\
        );

    \I__3155\ : SRMux
    port map (
            O => \N__12501\,
            I => \N__12356\
        );

    \I__3154\ : SRMux
    port map (
            O => \N__12500\,
            I => \N__12356\
        );

    \I__3153\ : SRMux
    port map (
            O => \N__12499\,
            I => \N__12356\
        );

    \I__3152\ : SRMux
    port map (
            O => \N__12498\,
            I => \N__12356\
        );

    \I__3151\ : SRMux
    port map (
            O => \N__12497\,
            I => \N__12356\
        );

    \I__3150\ : SRMux
    port map (
            O => \N__12496\,
            I => \N__12356\
        );

    \I__3149\ : SRMux
    port map (
            O => \N__12495\,
            I => \N__12356\
        );

    \I__3148\ : SRMux
    port map (
            O => \N__12494\,
            I => \N__12356\
        );

    \I__3147\ : SRMux
    port map (
            O => \N__12493\,
            I => \N__12356\
        );

    \I__3146\ : SRMux
    port map (
            O => \N__12492\,
            I => \N__12356\
        );

    \I__3145\ : SRMux
    port map (
            O => \N__12491\,
            I => \N__12356\
        );

    \I__3144\ : SRMux
    port map (
            O => \N__12490\,
            I => \N__12356\
        );

    \I__3143\ : SRMux
    port map (
            O => \N__12489\,
            I => \N__12356\
        );

    \I__3142\ : SRMux
    port map (
            O => \N__12488\,
            I => \N__12356\
        );

    \I__3141\ : SRMux
    port map (
            O => \N__12487\,
            I => \N__12356\
        );

    \I__3140\ : SRMux
    port map (
            O => \N__12486\,
            I => \N__12356\
        );

    \I__3139\ : SRMux
    port map (
            O => \N__12485\,
            I => \N__12356\
        );

    \I__3138\ : SRMux
    port map (
            O => \N__12484\,
            I => \N__12356\
        );

    \I__3137\ : SRMux
    port map (
            O => \N__12483\,
            I => \N__12356\
        );

    \I__3136\ : SRMux
    port map (
            O => \N__12482\,
            I => \N__12356\
        );

    \I__3135\ : SRMux
    port map (
            O => \N__12481\,
            I => \N__12356\
        );

    \I__3134\ : SRMux
    port map (
            O => \N__12480\,
            I => \N__12356\
        );

    \I__3133\ : SRMux
    port map (
            O => \N__12479\,
            I => \N__12356\
        );

    \I__3132\ : SRMux
    port map (
            O => \N__12478\,
            I => \N__12356\
        );

    \I__3131\ : SRMux
    port map (
            O => \N__12477\,
            I => \N__12356\
        );

    \I__3130\ : SRMux
    port map (
            O => \N__12476\,
            I => \N__12356\
        );

    \I__3129\ : SRMux
    port map (
            O => \N__12475\,
            I => \N__12356\
        );

    \I__3128\ : SRMux
    port map (
            O => \N__12474\,
            I => \N__12356\
        );

    \I__3127\ : SRMux
    port map (
            O => \N__12473\,
            I => \N__12356\
        );

    \I__3126\ : SRMux
    port map (
            O => \N__12472\,
            I => \N__12356\
        );

    \I__3125\ : SRMux
    port map (
            O => \N__12471\,
            I => \N__12356\
        );

    \I__3124\ : SRMux
    port map (
            O => \N__12470\,
            I => \N__12356\
        );

    \I__3123\ : SRMux
    port map (
            O => \N__12469\,
            I => \N__12356\
        );

    \I__3122\ : SRMux
    port map (
            O => \N__12468\,
            I => \N__12356\
        );

    \I__3121\ : SRMux
    port map (
            O => \N__12467\,
            I => \N__12356\
        );

    \I__3120\ : SRMux
    port map (
            O => \N__12466\,
            I => \N__12356\
        );

    \I__3119\ : SRMux
    port map (
            O => \N__12465\,
            I => \N__12356\
        );

    \I__3118\ : SRMux
    port map (
            O => \N__12464\,
            I => \N__12356\
        );

    \I__3117\ : SRMux
    port map (
            O => \N__12463\,
            I => \N__12356\
        );

    \I__3116\ : SRMux
    port map (
            O => \N__12462\,
            I => \N__12356\
        );

    \I__3115\ : Glb2LocalMux
    port map (
            O => \N__12459\,
            I => \N__12356\
        );

    \I__3114\ : GlobalMux
    port map (
            O => \N__12356\,
            I => \N__12353\
        );

    \I__3113\ : gio2CtrlBuf
    port map (
            O => \N__12353\,
            I => \RESETn_c_i_g\
        );

    \I__3112\ : InMux
    port map (
            O => \N__12350\,
            I => \N__12347\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__12347\,
            I => \READ_CYCLE_ACTIVE_rep11_i_ess\
        );

    \I__3110\ : IoInMux
    port map (
            O => \N__12344\,
            I => \N__12341\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__12341\,
            I => \N__12338\
        );

    \I__3108\ : Span4Mux_s3_h
    port map (
            O => \N__12338\,
            I => \N__12335\
        );

    \I__3107\ : Span4Mux_v
    port map (
            O => \N__12335\,
            I => \N__12332\
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__12332\,
            I => \N_192_i\
        );

    \I__3105\ : InMux
    port map (
            O => \N__12329\,
            I => \N__12326\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__12326\,
            I => \READ_CYCLE_ACTIVE_rep3_i_ess\
        );

    \I__3103\ : IoInMux
    port map (
            O => \N__12323\,
            I => \N__12320\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__12320\,
            I => \N__12317\
        );

    \I__3101\ : IoSpan4Mux
    port map (
            O => \N__12317\,
            I => \N__12314\
        );

    \I__3100\ : Span4Mux_s3_v
    port map (
            O => \N__12314\,
            I => \N__12311\
        );

    \I__3099\ : Span4Mux_v
    port map (
            O => \N__12311\,
            I => \N__12308\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__12308\,
            I => \N_184_i\
        );

    \I__3097\ : InMux
    port map (
            O => \N__12305\,
            I => \N__12302\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__12302\,
            I => \READ_CYCLE_ACTIVE_rep15_i_ess\
        );

    \I__3095\ : IoInMux
    port map (
            O => \N__12299\,
            I => \N__12296\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__12296\,
            I => \N__12293\
        );

    \I__3093\ : IoSpan4Mux
    port map (
            O => \N__12293\,
            I => \N__12290\
        );

    \I__3092\ : Span4Mux_s3_h
    port map (
            O => \N__12290\,
            I => \N__12287\
        );

    \I__3091\ : Odrv4
    port map (
            O => \N__12287\,
            I => \N_196_i\
        );

    \I__3090\ : InMux
    port map (
            O => \N__12284\,
            I => \N__12281\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__12281\,
            I => \READ_CYCLE_ACTIVE_rep1_i_ess\
        );

    \I__3088\ : IoInMux
    port map (
            O => \N__12278\,
            I => \N__12275\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__12275\,
            I => \N__12272\
        );

    \I__3086\ : Span12Mux_s4_h
    port map (
            O => \N__12272\,
            I => \N__12269\
        );

    \I__3085\ : Odrv12
    port map (
            O => \N__12269\,
            I => \N_182_i\
        );

    \I__3084\ : InMux
    port map (
            O => \N__12266\,
            I => \N__12263\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__12263\,
            I => \READ_CYCLE_ACTIVE_rep13_i_ess\
        );

    \I__3082\ : CascadeMux
    port map (
            O => \N__12260\,
            I => \N__12253\
        );

    \I__3081\ : InMux
    port map (
            O => \N__12259\,
            I => \N__12248\
        );

    \I__3080\ : InMux
    port map (
            O => \N__12258\,
            I => \N__12245\
        );

    \I__3079\ : InMux
    port map (
            O => \N__12257\,
            I => \N__12239\
        );

    \I__3078\ : InMux
    port map (
            O => \N__12256\,
            I => \N__12236\
        );

    \I__3077\ : InMux
    port map (
            O => \N__12253\,
            I => \N__12231\
        );

    \I__3076\ : InMux
    port map (
            O => \N__12252\,
            I => \N__12231\
        );

    \I__3075\ : InMux
    port map (
            O => \N__12251\,
            I => \N__12223\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__12248\,
            I => \N__12218\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__12245\,
            I => \N__12218\
        );

    \I__3072\ : InMux
    port map (
            O => \N__12244\,
            I => \N__12213\
        );

    \I__3071\ : InMux
    port map (
            O => \N__12243\,
            I => \N__12210\
        );

    \I__3070\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12207\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__12239\,
            I => \N__12197\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__12236\,
            I => \N__12197\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__12231\,
            I => \N__12194\
        );

    \I__3066\ : InMux
    port map (
            O => \N__12230\,
            I => \N__12189\
        );

    \I__3065\ : InMux
    port map (
            O => \N__12229\,
            I => \N__12189\
        );

    \I__3064\ : InMux
    port map (
            O => \N__12228\,
            I => \N__12186\
        );

    \I__3063\ : InMux
    port map (
            O => \N__12227\,
            I => \N__12183\
        );

    \I__3062\ : InMux
    port map (
            O => \N__12226\,
            I => \N__12180\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__12223\,
            I => \N__12175\
        );

    \I__3060\ : Span4Mux_v
    port map (
            O => \N__12218\,
            I => \N__12175\
        );

    \I__3059\ : InMux
    port map (
            O => \N__12217\,
            I => \N__12172\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__12216\,
            I => \N__12168\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__12213\,
            I => \N__12159\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__12210\,
            I => \N__12159\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__12207\,
            I => \N__12159\
        );

    \I__3054\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12156\
        );

    \I__3053\ : InMux
    port map (
            O => \N__12205\,
            I => \N__12153\
        );

    \I__3052\ : InMux
    port map (
            O => \N__12204\,
            I => \N__12150\
        );

    \I__3051\ : InMux
    port map (
            O => \N__12203\,
            I => \N__12147\
        );

    \I__3050\ : InMux
    port map (
            O => \N__12202\,
            I => \N__12144\
        );

    \I__3049\ : Span4Mux_v
    port map (
            O => \N__12197\,
            I => \N__12127\
        );

    \I__3048\ : Span4Mux_h
    port map (
            O => \N__12194\,
            I => \N__12127\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__12189\,
            I => \N__12127\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__12186\,
            I => \N__12127\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__12183\,
            I => \N__12127\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__12180\,
            I => \N__12127\
        );

    \I__3043\ : Span4Mux_h
    port map (
            O => \N__12175\,
            I => \N__12127\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__12172\,
            I => \N__12127\
        );

    \I__3041\ : InMux
    port map (
            O => \N__12171\,
            I => \N__12124\
        );

    \I__3040\ : InMux
    port map (
            O => \N__12168\,
            I => \N__12121\
        );

    \I__3039\ : InMux
    port map (
            O => \N__12167\,
            I => \N__12118\
        );

    \I__3038\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12113\
        );

    \I__3037\ : Span4Mux_v
    port map (
            O => \N__12159\,
            I => \N__12106\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__12156\,
            I => \N__12106\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__12153\,
            I => \N__12106\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__12150\,
            I => \N__12095\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__12147\,
            I => \N__12095\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__12144\,
            I => \N__12095\
        );

    \I__3031\ : Span4Mux_v
    port map (
            O => \N__12127\,
            I => \N__12095\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__12124\,
            I => \N__12095\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__12121\,
            I => \N__12084\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__12118\,
            I => \N__12084\
        );

    \I__3027\ : InMux
    port map (
            O => \N__12117\,
            I => \N__12081\
        );

    \I__3026\ : InMux
    port map (
            O => \N__12116\,
            I => \N__12078\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__12113\,
            I => \N__12075\
        );

    \I__3024\ : Span4Mux_v
    port map (
            O => \N__12106\,
            I => \N__12068\
        );

    \I__3023\ : Span4Mux_v
    port map (
            O => \N__12095\,
            I => \N__12068\
        );

    \I__3022\ : InMux
    port map (
            O => \N__12094\,
            I => \N__12065\
        );

    \I__3021\ : InMux
    port map (
            O => \N__12093\,
            I => \N__12062\
        );

    \I__3020\ : InMux
    port map (
            O => \N__12092\,
            I => \N__12059\
        );

    \I__3019\ : InMux
    port map (
            O => \N__12091\,
            I => \N__12056\
        );

    \I__3018\ : InMux
    port map (
            O => \N__12090\,
            I => \N__12053\
        );

    \I__3017\ : InMux
    port map (
            O => \N__12089\,
            I => \N__12039\
        );

    \I__3016\ : Span4Mux_v
    port map (
            O => \N__12084\,
            I => \N__12032\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__12081\,
            I => \N__12032\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__12078\,
            I => \N__12032\
        );

    \I__3013\ : Span4Mux_v
    port map (
            O => \N__12075\,
            I => \N__12029\
        );

    \I__3012\ : InMux
    port map (
            O => \N__12074\,
            I => \N__12024\
        );

    \I__3011\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12024\
        );

    \I__3010\ : Span4Mux_h
    port map (
            O => \N__12068\,
            I => \N__12017\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__12065\,
            I => \N__12017\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__12062\,
            I => \N__12014\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__12059\,
            I => \N__12008\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__12056\,
            I => \N__12008\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__12053\,
            I => \N__12005\
        );

    \I__3004\ : InMux
    port map (
            O => \N__12052\,
            I => \N__11998\
        );

    \I__3003\ : InMux
    port map (
            O => \N__12051\,
            I => \N__11998\
        );

    \I__3002\ : InMux
    port map (
            O => \N__12050\,
            I => \N__11998\
        );

    \I__3001\ : InMux
    port map (
            O => \N__12049\,
            I => \N__11995\
        );

    \I__3000\ : InMux
    port map (
            O => \N__12048\,
            I => \N__11986\
        );

    \I__2999\ : InMux
    port map (
            O => \N__12047\,
            I => \N__11986\
        );

    \I__2998\ : InMux
    port map (
            O => \N__12046\,
            I => \N__11986\
        );

    \I__2997\ : InMux
    port map (
            O => \N__12045\,
            I => \N__11981\
        );

    \I__2996\ : InMux
    port map (
            O => \N__12044\,
            I => \N__11981\
        );

    \I__2995\ : InMux
    port map (
            O => \N__12043\,
            I => \N__11976\
        );

    \I__2994\ : InMux
    port map (
            O => \N__12042\,
            I => \N__11976\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__12039\,
            I => \N__11966\
        );

    \I__2992\ : Sp12to4
    port map (
            O => \N__12032\,
            I => \N__11966\
        );

    \I__2991\ : Span4Mux_h
    port map (
            O => \N__12029\,
            I => \N__11961\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__12024\,
            I => \N__11961\
        );

    \I__2989\ : InMux
    port map (
            O => \N__12023\,
            I => \N__11956\
        );

    \I__2988\ : InMux
    port map (
            O => \N__12022\,
            I => \N__11956\
        );

    \I__2987\ : Span4Mux_h
    port map (
            O => \N__12017\,
            I => \N__11951\
        );

    \I__2986\ : Span4Mux_v
    port map (
            O => \N__12014\,
            I => \N__11951\
        );

    \I__2985\ : InMux
    port map (
            O => \N__12013\,
            I => \N__11948\
        );

    \I__2984\ : Span4Mux_v
    port map (
            O => \N__12008\,
            I => \N__11945\
        );

    \I__2983\ : Span4Mux_v
    port map (
            O => \N__12005\,
            I => \N__11942\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__11998\,
            I => \N__11939\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__11995\,
            I => \N__11934\
        );

    \I__2980\ : InMux
    port map (
            O => \N__11994\,
            I => \N__11929\
        );

    \I__2979\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11929\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__11986\,
            I => \N__11920\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__11981\,
            I => \N__11920\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__11976\,
            I => \N__11917\
        );

    \I__2975\ : InMux
    port map (
            O => \N__11975\,
            I => \N__11908\
        );

    \I__2974\ : InMux
    port map (
            O => \N__11974\,
            I => \N__11908\
        );

    \I__2973\ : InMux
    port map (
            O => \N__11973\,
            I => \N__11908\
        );

    \I__2972\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11908\
        );

    \I__2971\ : InMux
    port map (
            O => \N__11971\,
            I => \N__11905\
        );

    \I__2970\ : Span12Mux_v
    port map (
            O => \N__11966\,
            I => \N__11897\
        );

    \I__2969\ : Sp12to4
    port map (
            O => \N__11961\,
            I => \N__11894\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__11956\,
            I => \N__11891\
        );

    \I__2967\ : Span4Mux_v
    port map (
            O => \N__11951\,
            I => \N__11888\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__11948\,
            I => \N__11885\
        );

    \I__2965\ : Span4Mux_v
    port map (
            O => \N__11945\,
            I => \N__11882\
        );

    \I__2964\ : Span4Mux_h
    port map (
            O => \N__11942\,
            I => \N__11877\
        );

    \I__2963\ : Span4Mux_v
    port map (
            O => \N__11939\,
            I => \N__11877\
        );

    \I__2962\ : InMux
    port map (
            O => \N__11938\,
            I => \N__11874\
        );

    \I__2961\ : InMux
    port map (
            O => \N__11937\,
            I => \N__11871\
        );

    \I__2960\ : Span4Mux_v
    port map (
            O => \N__11934\,
            I => \N__11868\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__11929\,
            I => \N__11865\
        );

    \I__2958\ : InMux
    port map (
            O => \N__11928\,
            I => \N__11858\
        );

    \I__2957\ : InMux
    port map (
            O => \N__11927\,
            I => \N__11858\
        );

    \I__2956\ : InMux
    port map (
            O => \N__11926\,
            I => \N__11858\
        );

    \I__2955\ : InMux
    port map (
            O => \N__11925\,
            I => \N__11855\
        );

    \I__2954\ : Span4Mux_v
    port map (
            O => \N__11920\,
            I => \N__11848\
        );

    \I__2953\ : Span4Mux_h
    port map (
            O => \N__11917\,
            I => \N__11848\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__11908\,
            I => \N__11848\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__11905\,
            I => \N__11845\
        );

    \I__2950\ : InMux
    port map (
            O => \N__11904\,
            I => \N__11840\
        );

    \I__2949\ : InMux
    port map (
            O => \N__11903\,
            I => \N__11840\
        );

    \I__2948\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11833\
        );

    \I__2947\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11833\
        );

    \I__2946\ : InMux
    port map (
            O => \N__11900\,
            I => \N__11833\
        );

    \I__2945\ : Span12Mux_h
    port map (
            O => \N__11897\,
            I => \N__11830\
        );

    \I__2944\ : Span12Mux_v
    port map (
            O => \N__11894\,
            I => \N__11825\
        );

    \I__2943\ : Span12Mux_s9_h
    port map (
            O => \N__11891\,
            I => \N__11825\
        );

    \I__2942\ : Sp12to4
    port map (
            O => \N__11888\,
            I => \N__11820\
        );

    \I__2941\ : Span12Mux_v
    port map (
            O => \N__11885\,
            I => \N__11820\
        );

    \I__2940\ : Span4Mux_v
    port map (
            O => \N__11882\,
            I => \N__11815\
        );

    \I__2939\ : Span4Mux_v
    port map (
            O => \N__11877\,
            I => \N__11815\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__11874\,
            I => \N__11810\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__11871\,
            I => \N__11810\
        );

    \I__2936\ : Span4Mux_h
    port map (
            O => \N__11868\,
            I => \N__11801\
        );

    \I__2935\ : Span4Mux_v
    port map (
            O => \N__11865\,
            I => \N__11801\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__11858\,
            I => \N__11801\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__11855\,
            I => \N__11801\
        );

    \I__2932\ : Span4Mux_v
    port map (
            O => \N__11848\,
            I => \N__11792\
        );

    \I__2931\ : Span4Mux_h
    port map (
            O => \N__11845\,
            I => \N__11792\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__11840\,
            I => \N__11792\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__11833\,
            I => \N__11792\
        );

    \I__2928\ : Span12Mux_h
    port map (
            O => \N__11830\,
            I => \N__11789\
        );

    \I__2927\ : Span12Mux_h
    port map (
            O => \N__11825\,
            I => \N__11786\
        );

    \I__2926\ : Span12Mux_h
    port map (
            O => \N__11820\,
            I => \N__11779\
        );

    \I__2925\ : Sp12to4
    port map (
            O => \N__11815\,
            I => \N__11779\
        );

    \I__2924\ : Span12Mux_v
    port map (
            O => \N__11810\,
            I => \N__11779\
        );

    \I__2923\ : Span4Mux_v
    port map (
            O => \N__11801\,
            I => \N__11774\
        );

    \I__2922\ : Span4Mux_v
    port map (
            O => \N__11792\,
            I => \N__11774\
        );

    \I__2921\ : Odrv12
    port map (
            O => \N__11789\,
            I => \BGn_c\
        );

    \I__2920\ : Odrv12
    port map (
            O => \N__11786\,
            I => \BGn_c\
        );

    \I__2919\ : Odrv12
    port map (
            O => \N__11779\,
            I => \BGn_c\
        );

    \I__2918\ : Odrv4
    port map (
            O => \N__11774\,
            I => \BGn_c\
        );

    \I__2917\ : CascadeMux
    port map (
            O => \N__11765\,
            I => \N__11761\
        );

    \I__2916\ : InMux
    port map (
            O => \N__11764\,
            I => \N__11755\
        );

    \I__2915\ : InMux
    port map (
            O => \N__11761\,
            I => \N__11752\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__11760\,
            I => \N__11749\
        );

    \I__2913\ : CascadeMux
    port map (
            O => \N__11759\,
            I => \N__11745\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__11758\,
            I => \N__11741\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__11755\,
            I => \N__11734\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__11752\,
            I => \N__11734\
        );

    \I__2909\ : InMux
    port map (
            O => \N__11749\,
            I => \N__11731\
        );

    \I__2908\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11726\
        );

    \I__2907\ : InMux
    port map (
            O => \N__11745\,
            I => \N__11726\
        );

    \I__2906\ : InMux
    port map (
            O => \N__11744\,
            I => \N__11723\
        );

    \I__2905\ : InMux
    port map (
            O => \N__11741\,
            I => \N__11720\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__11740\,
            I => \N__11717\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__11739\,
            I => \N__11712\
        );

    \I__2902\ : Span4Mux_v
    port map (
            O => \N__11734\,
            I => \N__11692\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__11731\,
            I => \N__11692\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__11726\,
            I => \N__11692\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__11723\,
            I => \N__11692\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__11720\,
            I => \N__11692\
        );

    \I__2897\ : InMux
    port map (
            O => \N__11717\,
            I => \N__11689\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__11716\,
            I => \N__11685\
        );

    \I__2895\ : InMux
    port map (
            O => \N__11715\,
            I => \N__11677\
        );

    \I__2894\ : InMux
    port map (
            O => \N__11712\,
            I => \N__11677\
        );

    \I__2893\ : InMux
    port map (
            O => \N__11711\,
            I => \N__11677\
        );

    \I__2892\ : InMux
    port map (
            O => \N__11710\,
            I => \N__11674\
        );

    \I__2891\ : InMux
    port map (
            O => \N__11709\,
            I => \N__11671\
        );

    \I__2890\ : CascadeMux
    port map (
            O => \N__11708\,
            I => \N__11668\
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__11707\,
            I => \N__11663\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__11706\,
            I => \N__11659\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__11705\,
            I => \N__11656\
        );

    \I__2886\ : InMux
    port map (
            O => \N__11704\,
            I => \N__11651\
        );

    \I__2885\ : CascadeMux
    port map (
            O => \N__11703\,
            I => \N__11646\
        );

    \I__2884\ : Span4Mux_v
    port map (
            O => \N__11692\,
            I => \N__11641\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__11689\,
            I => \N__11641\
        );

    \I__2882\ : InMux
    port map (
            O => \N__11688\,
            I => \N__11636\
        );

    \I__2881\ : InMux
    port map (
            O => \N__11685\,
            I => \N__11636\
        );

    \I__2880\ : InMux
    port map (
            O => \N__11684\,
            I => \N__11633\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__11677\,
            I => \N__11623\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__11674\,
            I => \N__11623\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__11671\,
            I => \N__11623\
        );

    \I__2876\ : InMux
    port map (
            O => \N__11668\,
            I => \N__11618\
        );

    \I__2875\ : InMux
    port map (
            O => \N__11667\,
            I => \N__11618\
        );

    \I__2874\ : InMux
    port map (
            O => \N__11666\,
            I => \N__11609\
        );

    \I__2873\ : InMux
    port map (
            O => \N__11663\,
            I => \N__11609\
        );

    \I__2872\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11609\
        );

    \I__2871\ : InMux
    port map (
            O => \N__11659\,
            I => \N__11609\
        );

    \I__2870\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11602\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__11655\,
            I => \N__11598\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__11654\,
            I => \N__11590\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__11651\,
            I => \N__11581\
        );

    \I__2866\ : InMux
    port map (
            O => \N__11650\,
            I => \N__11576\
        );

    \I__2865\ : InMux
    port map (
            O => \N__11649\,
            I => \N__11576\
        );

    \I__2864\ : InMux
    port map (
            O => \N__11646\,
            I => \N__11573\
        );

    \I__2863\ : Span4Mux_v
    port map (
            O => \N__11641\,
            I => \N__11566\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__11636\,
            I => \N__11566\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__11633\,
            I => \N__11566\
        );

    \I__2860\ : InMux
    port map (
            O => \N__11632\,
            I => \N__11561\
        );

    \I__2859\ : InMux
    port map (
            O => \N__11631\,
            I => \N__11561\
        );

    \I__2858\ : CascadeMux
    port map (
            O => \N__11630\,
            I => \N__11555\
        );

    \I__2857\ : Span4Mux_v
    port map (
            O => \N__11623\,
            I => \N__11547\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__11618\,
            I => \N__11547\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__11609\,
            I => \N__11547\
        );

    \I__2854\ : InMux
    port map (
            O => \N__11608\,
            I => \N__11544\
        );

    \I__2853\ : InMux
    port map (
            O => \N__11607\,
            I => \N__11539\
        );

    \I__2852\ : InMux
    port map (
            O => \N__11606\,
            I => \N__11539\
        );

    \I__2851\ : InMux
    port map (
            O => \N__11605\,
            I => \N__11532\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__11602\,
            I => \N__11529\
        );

    \I__2849\ : InMux
    port map (
            O => \N__11601\,
            I => \N__11526\
        );

    \I__2848\ : InMux
    port map (
            O => \N__11598\,
            I => \N__11523\
        );

    \I__2847\ : InMux
    port map (
            O => \N__11597\,
            I => \N__11515\
        );

    \I__2846\ : InMux
    port map (
            O => \N__11596\,
            I => \N__11515\
        );

    \I__2845\ : InMux
    port map (
            O => \N__11595\,
            I => \N__11515\
        );

    \I__2844\ : InMux
    port map (
            O => \N__11594\,
            I => \N__11508\
        );

    \I__2843\ : InMux
    port map (
            O => \N__11593\,
            I => \N__11508\
        );

    \I__2842\ : InMux
    port map (
            O => \N__11590\,
            I => \N__11502\
        );

    \I__2841\ : InMux
    port map (
            O => \N__11589\,
            I => \N__11499\
        );

    \I__2840\ : InMux
    port map (
            O => \N__11588\,
            I => \N__11496\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__11587\,
            I => \N__11493\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__11586\,
            I => \N__11490\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__11585\,
            I => \N__11485\
        );

    \I__2836\ : CascadeMux
    port map (
            O => \N__11584\,
            I => \N__11482\
        );

    \I__2835\ : Span4Mux_v
    port map (
            O => \N__11581\,
            I => \N__11479\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__11576\,
            I => \N__11474\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__11573\,
            I => \N__11474\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__11566\,
            I => \N__11469\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__11561\,
            I => \N__11469\
        );

    \I__2830\ : InMux
    port map (
            O => \N__11560\,
            I => \N__11466\
        );

    \I__2829\ : InMux
    port map (
            O => \N__11559\,
            I => \N__11461\
        );

    \I__2828\ : InMux
    port map (
            O => \N__11558\,
            I => \N__11461\
        );

    \I__2827\ : InMux
    port map (
            O => \N__11555\,
            I => \N__11458\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__11554\,
            I => \N__11454\
        );

    \I__2825\ : Span4Mux_v
    port map (
            O => \N__11547\,
            I => \N__11448\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__11544\,
            I => \N__11448\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__11539\,
            I => \N__11445\
        );

    \I__2822\ : InMux
    port map (
            O => \N__11538\,
            I => \N__11442\
        );

    \I__2821\ : InMux
    port map (
            O => \N__11537\,
            I => \N__11435\
        );

    \I__2820\ : InMux
    port map (
            O => \N__11536\,
            I => \N__11435\
        );

    \I__2819\ : InMux
    port map (
            O => \N__11535\,
            I => \N__11435\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__11532\,
            I => \N__11432\
        );

    \I__2817\ : Span4Mux_h
    port map (
            O => \N__11529\,
            I => \N__11425\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__11526\,
            I => \N__11425\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__11523\,
            I => \N__11425\
        );

    \I__2814\ : InMux
    port map (
            O => \N__11522\,
            I => \N__11422\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__11515\,
            I => \N__11419\
        );

    \I__2812\ : InMux
    port map (
            O => \N__11514\,
            I => \N__11416\
        );

    \I__2811\ : InMux
    port map (
            O => \N__11513\,
            I => \N__11413\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__11508\,
            I => \N__11410\
        );

    \I__2809\ : InMux
    port map (
            O => \N__11507\,
            I => \N__11407\
        );

    \I__2808\ : InMux
    port map (
            O => \N__11506\,
            I => \N__11404\
        );

    \I__2807\ : InMux
    port map (
            O => \N__11505\,
            I => \N__11401\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__11502\,
            I => \N__11396\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__11499\,
            I => \N__11396\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__11496\,
            I => \N__11393\
        );

    \I__2803\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11390\
        );

    \I__2802\ : InMux
    port map (
            O => \N__11490\,
            I => \N__11383\
        );

    \I__2801\ : InMux
    port map (
            O => \N__11489\,
            I => \N__11383\
        );

    \I__2800\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11383\
        );

    \I__2799\ : InMux
    port map (
            O => \N__11485\,
            I => \N__11380\
        );

    \I__2798\ : InMux
    port map (
            O => \N__11482\,
            I => \N__11377\
        );

    \I__2797\ : Span4Mux_v
    port map (
            O => \N__11479\,
            I => \N__11374\
        );

    \I__2796\ : Span4Mux_v
    port map (
            O => \N__11474\,
            I => \N__11371\
        );

    \I__2795\ : Span4Mux_h
    port map (
            O => \N__11469\,
            I => \N__11364\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__11466\,
            I => \N__11364\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__11461\,
            I => \N__11364\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__11458\,
            I => \N__11361\
        );

    \I__2791\ : InMux
    port map (
            O => \N__11457\,
            I => \N__11356\
        );

    \I__2790\ : InMux
    port map (
            O => \N__11454\,
            I => \N__11356\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__11453\,
            I => \N__11353\
        );

    \I__2788\ : Span4Mux_v
    port map (
            O => \N__11448\,
            I => \N__11346\
        );

    \I__2787\ : Span4Mux_v
    port map (
            O => \N__11445\,
            I => \N__11346\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__11442\,
            I => \N__11346\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__11435\,
            I => \N__11343\
        );

    \I__2784\ : Span4Mux_v
    port map (
            O => \N__11432\,
            I => \N__11339\
        );

    \I__2783\ : Span4Mux_h
    port map (
            O => \N__11425\,
            I => \N__11334\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__11422\,
            I => \N__11334\
        );

    \I__2781\ : Span4Mux_h
    port map (
            O => \N__11419\,
            I => \N__11327\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__11416\,
            I => \N__11327\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__11413\,
            I => \N__11327\
        );

    \I__2778\ : Span4Mux_h
    port map (
            O => \N__11410\,
            I => \N__11324\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__11407\,
            I => \N__11321\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__11404\,
            I => \N__11316\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__11401\,
            I => \N__11316\
        );

    \I__2774\ : Span12Mux_v
    port map (
            O => \N__11396\,
            I => \N__11309\
        );

    \I__2773\ : Span12Mux_s6_h
    port map (
            O => \N__11393\,
            I => \N__11309\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__11390\,
            I => \N__11309\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__11383\,
            I => \N__11306\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__11380\,
            I => \N__11303\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__11377\,
            I => \N__11300\
        );

    \I__2768\ : Span4Mux_v
    port map (
            O => \N__11374\,
            I => \N__11293\
        );

    \I__2767\ : Span4Mux_h
    port map (
            O => \N__11371\,
            I => \N__11293\
        );

    \I__2766\ : Span4Mux_v
    port map (
            O => \N__11364\,
            I => \N__11293\
        );

    \I__2765\ : Span12Mux_s6_h
    port map (
            O => \N__11361\,
            I => \N__11290\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__11356\,
            I => \N__11287\
        );

    \I__2763\ : InMux
    port map (
            O => \N__11353\,
            I => \N__11284\
        );

    \I__2762\ : Span4Mux_v
    port map (
            O => \N__11346\,
            I => \N__11279\
        );

    \I__2761\ : Span4Mux_v
    port map (
            O => \N__11343\,
            I => \N__11279\
        );

    \I__2760\ : InMux
    port map (
            O => \N__11342\,
            I => \N__11276\
        );

    \I__2759\ : Span4Mux_v
    port map (
            O => \N__11339\,
            I => \N__11271\
        );

    \I__2758\ : Span4Mux_h
    port map (
            O => \N__11334\,
            I => \N__11271\
        );

    \I__2757\ : Span4Mux_h
    port map (
            O => \N__11327\,
            I => \N__11268\
        );

    \I__2756\ : Span4Mux_v
    port map (
            O => \N__11324\,
            I => \N__11265\
        );

    \I__2755\ : Span4Mux_v
    port map (
            O => \N__11321\,
            I => \N__11262\
        );

    \I__2754\ : Span12Mux_v
    port map (
            O => \N__11316\,
            I => \N__11259\
        );

    \I__2753\ : Span12Mux_h
    port map (
            O => \N__11309\,
            I => \N__11254\
        );

    \I__2752\ : Span12Mux_h
    port map (
            O => \N__11306\,
            I => \N__11254\
        );

    \I__2751\ : Span12Mux_h
    port map (
            O => \N__11303\,
            I => \N__11251\
        );

    \I__2750\ : Span12Mux_v
    port map (
            O => \N__11300\,
            I => \N__11246\
        );

    \I__2749\ : Sp12to4
    port map (
            O => \N__11293\,
            I => \N__11246\
        );

    \I__2748\ : Span12Mux_h
    port map (
            O => \N__11290\,
            I => \N__11241\
        );

    \I__2747\ : Span12Mux_h
    port map (
            O => \N__11287\,
            I => \N__11241\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__11284\,
            I => \N__11238\
        );

    \I__2745\ : Sp12to4
    port map (
            O => \N__11279\,
            I => \N__11233\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__11276\,
            I => \N__11233\
        );

    \I__2743\ : Span4Mux_v
    port map (
            O => \N__11271\,
            I => \N__11230\
        );

    \I__2742\ : Span4Mux_v
    port map (
            O => \N__11268\,
            I => \N__11227\
        );

    \I__2741\ : IoSpan4Mux
    port map (
            O => \N__11265\,
            I => \N__11224\
        );

    \I__2740\ : Span4Mux_v
    port map (
            O => \N__11262\,
            I => \N__11221\
        );

    \I__2739\ : Span12Mux_h
    port map (
            O => \N__11259\,
            I => \N__11216\
        );

    \I__2738\ : Span12Mux_v
    port map (
            O => \N__11254\,
            I => \N__11216\
        );

    \I__2737\ : Span12Mux_v
    port map (
            O => \N__11251\,
            I => \N__11211\
        );

    \I__2736\ : Span12Mux_h
    port map (
            O => \N__11246\,
            I => \N__11211\
        );

    \I__2735\ : Span12Mux_v
    port map (
            O => \N__11241\,
            I => \N__11204\
        );

    \I__2734\ : Span12Mux_h
    port map (
            O => \N__11238\,
            I => \N__11204\
        );

    \I__2733\ : Span12Mux_h
    port map (
            O => \N__11233\,
            I => \N__11204\
        );

    \I__2732\ : Span4Mux_h
    port map (
            O => \N__11230\,
            I => \N__11199\
        );

    \I__2731\ : Span4Mux_h
    port map (
            O => \N__11227\,
            I => \N__11199\
        );

    \I__2730\ : IoSpan4Mux
    port map (
            O => \N__11224\,
            I => \N__11194\
        );

    \I__2729\ : IoSpan4Mux
    port map (
            O => \N__11221\,
            I => \N__11194\
        );

    \I__2728\ : Odrv12
    port map (
            O => \N__11216\,
            I => \TS_CPUn_c\
        );

    \I__2727\ : Odrv12
    port map (
            O => \N__11211\,
            I => \TS_CPUn_c\
        );

    \I__2726\ : Odrv12
    port map (
            O => \N__11204\,
            I => \TS_CPUn_c\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__11199\,
            I => \TS_CPUn_c\
        );

    \I__2724\ : Odrv4
    port map (
            O => \N__11194\,
            I => \TS_CPUn_c\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__11183\,
            I => \N__11178\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__11182\,
            I => \N__11175\
        );

    \I__2721\ : InMux
    port map (
            O => \N__11181\,
            I => \N__11169\
        );

    \I__2720\ : InMux
    port map (
            O => \N__11178\,
            I => \N__11169\
        );

    \I__2719\ : InMux
    port map (
            O => \N__11175\,
            I => \N__11163\
        );

    \I__2718\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11158\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__11169\,
            I => \N__11154\
        );

    \I__2716\ : InMux
    port map (
            O => \N__11168\,
            I => \N__11151\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__11167\,
            I => \N__11145\
        );

    \I__2714\ : CascadeMux
    port map (
            O => \N__11166\,
            I => \N__11139\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__11163\,
            I => \N__11134\
        );

    \I__2712\ : InMux
    port map (
            O => \N__11162\,
            I => \N__11127\
        );

    \I__2711\ : InMux
    port map (
            O => \N__11161\,
            I => \N__11123\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__11158\,
            I => \N__11120\
        );

    \I__2709\ : InMux
    port map (
            O => \N__11157\,
            I => \N__11117\
        );

    \I__2708\ : Span4Mux_v
    port map (
            O => \N__11154\,
            I => \N__11114\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__11151\,
            I => \N__11110\
        );

    \I__2706\ : InMux
    port map (
            O => \N__11150\,
            I => \N__11104\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11104\
        );

    \I__2704\ : InMux
    port map (
            O => \N__11148\,
            I => \N__11101\
        );

    \I__2703\ : InMux
    port map (
            O => \N__11145\,
            I => \N__11098\
        );

    \I__2702\ : InMux
    port map (
            O => \N__11144\,
            I => \N__11095\
        );

    \I__2701\ : InMux
    port map (
            O => \N__11143\,
            I => \N__11092\
        );

    \I__2700\ : InMux
    port map (
            O => \N__11142\,
            I => \N__11087\
        );

    \I__2699\ : InMux
    port map (
            O => \N__11139\,
            I => \N__11087\
        );

    \I__2698\ : InMux
    port map (
            O => \N__11138\,
            I => \N__11084\
        );

    \I__2697\ : CascadeMux
    port map (
            O => \N__11137\,
            I => \N__11080\
        );

    \I__2696\ : Span4Mux_h
    port map (
            O => \N__11134\,
            I => \N__11073\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__11133\,
            I => \N__11070\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__11132\,
            I => \N__11061\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__11131\,
            I => \N__11058\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__11130\,
            I => \N__11055\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__11127\,
            I => \N__11050\
        );

    \I__2690\ : InMux
    port map (
            O => \N__11126\,
            I => \N__11047\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__11123\,
            I => \N__11044\
        );

    \I__2688\ : Span4Mux_v
    port map (
            O => \N__11120\,
            I => \N__11039\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__11117\,
            I => \N__11039\
        );

    \I__2686\ : Span4Mux_v
    port map (
            O => \N__11114\,
            I => \N__11034\
        );

    \I__2685\ : InMux
    port map (
            O => \N__11113\,
            I => \N__11031\
        );

    \I__2684\ : Span4Mux_v
    port map (
            O => \N__11110\,
            I => \N__11028\
        );

    \I__2683\ : InMux
    port map (
            O => \N__11109\,
            I => \N__11025\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__11104\,
            I => \N__11016\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__11101\,
            I => \N__11016\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__11098\,
            I => \N__11016\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__11095\,
            I => \N__11007\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__11092\,
            I => \N__11007\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11087\,
            I => \N__11007\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__11084\,
            I => \N__11007\
        );

    \I__2675\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11004\
        );

    \I__2674\ : InMux
    port map (
            O => \N__11080\,
            I => \N__11001\
        );

    \I__2673\ : InMux
    port map (
            O => \N__11079\,
            I => \N__10998\
        );

    \I__2672\ : InMux
    port map (
            O => \N__11078\,
            I => \N__10995\
        );

    \I__2671\ : InMux
    port map (
            O => \N__11077\,
            I => \N__10989\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__11076\,
            I => \N__10986\
        );

    \I__2669\ : Span4Mux_v
    port map (
            O => \N__11073\,
            I => \N__10983\
        );

    \I__2668\ : InMux
    port map (
            O => \N__11070\,
            I => \N__10980\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__11069\,
            I => \N__10977\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__11068\,
            I => \N__10974\
        );

    \I__2665\ : CascadeMux
    port map (
            O => \N__11067\,
            I => \N__10970\
        );

    \I__2664\ : InMux
    port map (
            O => \N__11066\,
            I => \N__10962\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__11065\,
            I => \N__10958\
        );

    \I__2662\ : CascadeMux
    port map (
            O => \N__11064\,
            I => \N__10955\
        );

    \I__2661\ : InMux
    port map (
            O => \N__11061\,
            I => \N__10946\
        );

    \I__2660\ : InMux
    port map (
            O => \N__11058\,
            I => \N__10946\
        );

    \I__2659\ : InMux
    port map (
            O => \N__11055\,
            I => \N__10946\
        );

    \I__2658\ : InMux
    port map (
            O => \N__11054\,
            I => \N__10943\
        );

    \I__2657\ : InMux
    port map (
            O => \N__11053\,
            I => \N__10940\
        );

    \I__2656\ : Span4Mux_h
    port map (
            O => \N__11050\,
            I => \N__10935\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__11047\,
            I => \N__10935\
        );

    \I__2654\ : Span4Mux_v
    port map (
            O => \N__11044\,
            I => \N__10932\
        );

    \I__2653\ : Span4Mux_h
    port map (
            O => \N__11039\,
            I => \N__10929\
        );

    \I__2652\ : InMux
    port map (
            O => \N__11038\,
            I => \N__10926\
        );

    \I__2651\ : InMux
    port map (
            O => \N__11037\,
            I => \N__10923\
        );

    \I__2650\ : Span4Mux_h
    port map (
            O => \N__11034\,
            I => \N__10918\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__11031\,
            I => \N__10918\
        );

    \I__2648\ : Span4Mux_v
    port map (
            O => \N__11028\,
            I => \N__10913\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__11025\,
            I => \N__10913\
        );

    \I__2646\ : InMux
    port map (
            O => \N__11024\,
            I => \N__10908\
        );

    \I__2645\ : InMux
    port map (
            O => \N__11023\,
            I => \N__10908\
        );

    \I__2644\ : Span4Mux_v
    port map (
            O => \N__11016\,
            I => \N__10905\
        );

    \I__2643\ : Span4Mux_v
    port map (
            O => \N__11007\,
            I => \N__10894\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__11004\,
            I => \N__10894\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__11001\,
            I => \N__10894\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__10998\,
            I => \N__10894\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__10995\,
            I => \N__10894\
        );

    \I__2638\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10891\
        );

    \I__2637\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10888\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__10992\,
            I => \N__10885\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__10989\,
            I => \N__10880\
        );

    \I__2634\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10877\
        );

    \I__2633\ : Span4Mux_v
    port map (
            O => \N__10983\,
            I => \N__10871\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__10980\,
            I => \N__10871\
        );

    \I__2631\ : InMux
    port map (
            O => \N__10977\,
            I => \N__10866\
        );

    \I__2630\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10866\
        );

    \I__2629\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10859\
        );

    \I__2628\ : InMux
    port map (
            O => \N__10970\,
            I => \N__10859\
        );

    \I__2627\ : InMux
    port map (
            O => \N__10969\,
            I => \N__10859\
        );

    \I__2626\ : InMux
    port map (
            O => \N__10968\,
            I => \N__10856\
        );

    \I__2625\ : CascadeMux
    port map (
            O => \N__10967\,
            I => \N__10848\
        );

    \I__2624\ : CascadeMux
    port map (
            O => \N__10966\,
            I => \N__10844\
        );

    \I__2623\ : CascadeMux
    port map (
            O => \N__10965\,
            I => \N__10840\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__10962\,
            I => \N__10836\
        );

    \I__2621\ : InMux
    port map (
            O => \N__10961\,
            I => \N__10831\
        );

    \I__2620\ : InMux
    port map (
            O => \N__10958\,
            I => \N__10831\
        );

    \I__2619\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10828\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__10954\,
            I => \N__10825\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__10953\,
            I => \N__10821\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__10946\,
            I => \N__10813\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__10943\,
            I => \N__10813\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__10940\,
            I => \N__10813\
        );

    \I__2613\ : Span4Mux_v
    port map (
            O => \N__10935\,
            I => \N__10810\
        );

    \I__2612\ : Span4Mux_h
    port map (
            O => \N__10932\,
            I => \N__10801\
        );

    \I__2611\ : Span4Mux_v
    port map (
            O => \N__10929\,
            I => \N__10801\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__10926\,
            I => \N__10801\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__10923\,
            I => \N__10801\
        );

    \I__2608\ : Span4Mux_v
    port map (
            O => \N__10918\,
            I => \N__10794\
        );

    \I__2607\ : Span4Mux_v
    port map (
            O => \N__10913\,
            I => \N__10794\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__10908\,
            I => \N__10794\
        );

    \I__2605\ : Span4Mux_v
    port map (
            O => \N__10905\,
            I => \N__10785\
        );

    \I__2604\ : Span4Mux_v
    port map (
            O => \N__10894\,
            I => \N__10785\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__10891\,
            I => \N__10785\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__10888\,
            I => \N__10785\
        );

    \I__2601\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10782\
        );

    \I__2600\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10779\
        );

    \I__2599\ : InMux
    port map (
            O => \N__10883\,
            I => \N__10776\
        );

    \I__2598\ : Span4Mux_h
    port map (
            O => \N__10880\,
            I => \N__10771\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__10877\,
            I => \N__10771\
        );

    \I__2596\ : InMux
    port map (
            O => \N__10876\,
            I => \N__10768\
        );

    \I__2595\ : Span4Mux_h
    port map (
            O => \N__10871\,
            I => \N__10765\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__10866\,
            I => \N__10758\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__10859\,
            I => \N__10758\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__10856\,
            I => \N__10758\
        );

    \I__2591\ : InMux
    port map (
            O => \N__10855\,
            I => \N__10751\
        );

    \I__2590\ : InMux
    port map (
            O => \N__10854\,
            I => \N__10751\
        );

    \I__2589\ : InMux
    port map (
            O => \N__10853\,
            I => \N__10751\
        );

    \I__2588\ : InMux
    port map (
            O => \N__10852\,
            I => \N__10746\
        );

    \I__2587\ : InMux
    port map (
            O => \N__10851\,
            I => \N__10746\
        );

    \I__2586\ : InMux
    port map (
            O => \N__10848\,
            I => \N__10737\
        );

    \I__2585\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10737\
        );

    \I__2584\ : InMux
    port map (
            O => \N__10844\,
            I => \N__10737\
        );

    \I__2583\ : InMux
    port map (
            O => \N__10843\,
            I => \N__10737\
        );

    \I__2582\ : InMux
    port map (
            O => \N__10840\,
            I => \N__10732\
        );

    \I__2581\ : InMux
    port map (
            O => \N__10839\,
            I => \N__10732\
        );

    \I__2580\ : Span4Mux_v
    port map (
            O => \N__10836\,
            I => \N__10725\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__10831\,
            I => \N__10725\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__10828\,
            I => \N__10725\
        );

    \I__2577\ : InMux
    port map (
            O => \N__10825\,
            I => \N__10718\
        );

    \I__2576\ : InMux
    port map (
            O => \N__10824\,
            I => \N__10718\
        );

    \I__2575\ : InMux
    port map (
            O => \N__10821\,
            I => \N__10718\
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__10820\,
            I => \N__10715\
        );

    \I__2573\ : Span4Mux_v
    port map (
            O => \N__10813\,
            I => \N__10712\
        );

    \I__2572\ : Span4Mux_h
    port map (
            O => \N__10810\,
            I => \N__10707\
        );

    \I__2571\ : Span4Mux_v
    port map (
            O => \N__10801\,
            I => \N__10707\
        );

    \I__2570\ : Span4Mux_v
    port map (
            O => \N__10794\,
            I => \N__10704\
        );

    \I__2569\ : Span4Mux_v
    port map (
            O => \N__10785\,
            I => \N__10694\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__10782\,
            I => \N__10694\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__10779\,
            I => \N__10694\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__10776\,
            I => \N__10694\
        );

    \I__2565\ : Span4Mux_v
    port map (
            O => \N__10771\,
            I => \N__10690\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__10768\,
            I => \N__10687\
        );

    \I__2563\ : Span4Mux_v
    port map (
            O => \N__10765\,
            I => \N__10683\
        );

    \I__2562\ : Span12Mux_s11_v
    port map (
            O => \N__10758\,
            I => \N__10672\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__10751\,
            I => \N__10672\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__10746\,
            I => \N__10672\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__10737\,
            I => \N__10672\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__10732\,
            I => \N__10672\
        );

    \I__2557\ : Span4Mux_v
    port map (
            O => \N__10725\,
            I => \N__10669\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__10718\,
            I => \N__10666\
        );

    \I__2555\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10663\
        );

    \I__2554\ : Sp12to4
    port map (
            O => \N__10712\,
            I => \N__10658\
        );

    \I__2553\ : Sp12to4
    port map (
            O => \N__10707\,
            I => \N__10658\
        );

    \I__2552\ : Span4Mux_v
    port map (
            O => \N__10704\,
            I => \N__10655\
        );

    \I__2551\ : InMux
    port map (
            O => \N__10703\,
            I => \N__10652\
        );

    \I__2550\ : Span4Mux_v
    port map (
            O => \N__10694\,
            I => \N__10649\
        );

    \I__2549\ : InMux
    port map (
            O => \N__10693\,
            I => \N__10646\
        );

    \I__2548\ : Span4Mux_h
    port map (
            O => \N__10690\,
            I => \N__10643\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__10687\,
            I => \N__10640\
        );

    \I__2546\ : InMux
    port map (
            O => \N__10686\,
            I => \N__10637\
        );

    \I__2545\ : Span4Mux_v
    port map (
            O => \N__10683\,
            I => \N__10634\
        );

    \I__2544\ : Span12Mux_v
    port map (
            O => \N__10672\,
            I => \N__10625\
        );

    \I__2543\ : Sp12to4
    port map (
            O => \N__10669\,
            I => \N__10625\
        );

    \I__2542\ : Span12Mux_s8_v
    port map (
            O => \N__10666\,
            I => \N__10625\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__10663\,
            I => \N__10625\
        );

    \I__2540\ : Span12Mux_h
    port map (
            O => \N__10658\,
            I => \N__10622\
        );

    \I__2539\ : Sp12to4
    port map (
            O => \N__10655\,
            I => \N__10613\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__10652\,
            I => \N__10613\
        );

    \I__2537\ : Sp12to4
    port map (
            O => \N__10649\,
            I => \N__10613\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10646\,
            I => \N__10613\
        );

    \I__2535\ : Span4Mux_h
    port map (
            O => \N__10643\,
            I => \N__10606\
        );

    \I__2534\ : Span4Mux_v
    port map (
            O => \N__10640\,
            I => \N__10606\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__10637\,
            I => \N__10606\
        );

    \I__2532\ : Span4Mux_v
    port map (
            O => \N__10634\,
            I => \N__10603\
        );

    \I__2531\ : Span12Mux_h
    port map (
            O => \N__10625\,
            I => \N__10596\
        );

    \I__2530\ : Span12Mux_v
    port map (
            O => \N__10622\,
            I => \N__10596\
        );

    \I__2529\ : Span12Mux_h
    port map (
            O => \N__10613\,
            I => \N__10596\
        );

    \I__2528\ : Span4Mux_v
    port map (
            O => \N__10606\,
            I => \N__10593\
        );

    \I__2527\ : Odrv4
    port map (
            O => \N__10603\,
            I => \LBENn_c\
        );

    \I__2526\ : Odrv12
    port map (
            O => \N__10596\,
            I => \LBENn_c\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__10593\,
            I => \LBENn_c\
        );

    \I__2524\ : InMux
    port map (
            O => \N__10586\,
            I => \N__10577\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__10585\,
            I => \N__10574\
        );

    \I__2522\ : InMux
    port map (
            O => \N__10584\,
            I => \N__10564\
        );

    \I__2521\ : InMux
    port map (
            O => \N__10583\,
            I => \N__10561\
        );

    \I__2520\ : InMux
    port map (
            O => \N__10582\,
            I => \N__10558\
        );

    \I__2519\ : InMux
    port map (
            O => \N__10581\,
            I => \N__10555\
        );

    \I__2518\ : IoInMux
    port map (
            O => \N__10580\,
            I => \N__10551\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__10577\,
            I => \N__10545\
        );

    \I__2516\ : InMux
    port map (
            O => \N__10574\,
            I => \N__10542\
        );

    \I__2515\ : InMux
    port map (
            O => \N__10573\,
            I => \N__10539\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__10572\,
            I => \N__10536\
        );

    \I__2513\ : InMux
    port map (
            O => \N__10571\,
            I => \N__10532\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__10570\,
            I => \N__10529\
        );

    \I__2511\ : InMux
    port map (
            O => \N__10569\,
            I => \N__10524\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__10568\,
            I => \N__10521\
        );

    \I__2509\ : InMux
    port map (
            O => \N__10567\,
            I => \N__10518\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10564\,
            I => \N__10511\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__10561\,
            I => \N__10511\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__10558\,
            I => \N__10511\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__10555\,
            I => \N__10508\
        );

    \I__2504\ : InMux
    port map (
            O => \N__10554\,
            I => \N__10505\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10551\,
            I => \N__10499\
        );

    \I__2502\ : CascadeMux
    port map (
            O => \N__10550\,
            I => \N__10495\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__10549\,
            I => \N__10490\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__10548\,
            I => \N__10487\
        );

    \I__2499\ : Span4Mux_v
    port map (
            O => \N__10545\,
            I => \N__10478\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__10542\,
            I => \N__10478\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__10539\,
            I => \N__10478\
        );

    \I__2496\ : InMux
    port map (
            O => \N__10536\,
            I => \N__10473\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10535\,
            I => \N__10473\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__10532\,
            I => \N__10470\
        );

    \I__2493\ : InMux
    port map (
            O => \N__10529\,
            I => \N__10465\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10528\,
            I => \N__10465\
        );

    \I__2491\ : InMux
    port map (
            O => \N__10527\,
            I => \N__10462\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10524\,
            I => \N__10458\
        );

    \I__2489\ : InMux
    port map (
            O => \N__10521\,
            I => \N__10455\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__10518\,
            I => \N__10451\
        );

    \I__2487\ : Span4Mux_v
    port map (
            O => \N__10511\,
            I => \N__10434\
        );

    \I__2486\ : Span4Mux_h
    port map (
            O => \N__10508\,
            I => \N__10434\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__10505\,
            I => \N__10434\
        );

    \I__2484\ : InMux
    port map (
            O => \N__10504\,
            I => \N__10431\
        );

    \I__2483\ : InMux
    port map (
            O => \N__10503\,
            I => \N__10428\
        );

    \I__2482\ : InMux
    port map (
            O => \N__10502\,
            I => \N__10425\
        );

    \I__2481\ : Span4Mux_s3_v
    port map (
            O => \N__10499\,
            I => \N__10422\
        );

    \I__2480\ : InMux
    port map (
            O => \N__10498\,
            I => \N__10419\
        );

    \I__2479\ : InMux
    port map (
            O => \N__10495\,
            I => \N__10416\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10494\,
            I => \N__10411\
        );

    \I__2477\ : InMux
    port map (
            O => \N__10493\,
            I => \N__10411\
        );

    \I__2476\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10406\
        );

    \I__2475\ : InMux
    port map (
            O => \N__10487\,
            I => \N__10406\
        );

    \I__2474\ : InMux
    port map (
            O => \N__10486\,
            I => \N__10403\
        );

    \I__2473\ : InMux
    port map (
            O => \N__10485\,
            I => \N__10400\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__10478\,
            I => \N__10395\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__10473\,
            I => \N__10395\
        );

    \I__2470\ : Span4Mux_v
    port map (
            O => \N__10470\,
            I => \N__10392\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__10465\,
            I => \N__10389\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__10462\,
            I => \N__10386\
        );

    \I__2467\ : InMux
    port map (
            O => \N__10461\,
            I => \N__10383\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__10458\,
            I => \N__10376\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__10455\,
            I => \N__10376\
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__10454\,
            I => \N__10373\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__10451\,
            I => \N__10369\
        );

    \I__2462\ : InMux
    port map (
            O => \N__10450\,
            I => \N__10366\
        );

    \I__2461\ : InMux
    port map (
            O => \N__10449\,
            I => \N__10361\
        );

    \I__2460\ : InMux
    port map (
            O => \N__10448\,
            I => \N__10361\
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__10447\,
            I => \N__10358\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__10446\,
            I => \N__10355\
        );

    \I__2457\ : CascadeMux
    port map (
            O => \N__10445\,
            I => \N__10352\
        );

    \I__2456\ : InMux
    port map (
            O => \N__10444\,
            I => \N__10347\
        );

    \I__2455\ : InMux
    port map (
            O => \N__10443\,
            I => \N__10340\
        );

    \I__2454\ : InMux
    port map (
            O => \N__10442\,
            I => \N__10340\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10441\,
            I => \N__10340\
        );

    \I__2452\ : Span4Mux_v
    port map (
            O => \N__10434\,
            I => \N__10327\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__10431\,
            I => \N__10327\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10428\,
            I => \N__10327\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__10425\,
            I => \N__10327\
        );

    \I__2448\ : Span4Mux_v
    port map (
            O => \N__10422\,
            I => \N__10312\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__10419\,
            I => \N__10312\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__10416\,
            I => \N__10312\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__10411\,
            I => \N__10312\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__10406\,
            I => \N__10312\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__10403\,
            I => \N__10312\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__10400\,
            I => \N__10312\
        );

    \I__2441\ : Span4Mux_v
    port map (
            O => \N__10395\,
            I => \N__10309\
        );

    \I__2440\ : Span4Mux_h
    port map (
            O => \N__10392\,
            I => \N__10300\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__10389\,
            I => \N__10300\
        );

    \I__2438\ : Span4Mux_h
    port map (
            O => \N__10386\,
            I => \N__10300\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__10383\,
            I => \N__10300\
        );

    \I__2436\ : InMux
    port map (
            O => \N__10382\,
            I => \N__10297\
        );

    \I__2435\ : InMux
    port map (
            O => \N__10381\,
            I => \N__10294\
        );

    \I__2434\ : Span4Mux_v
    port map (
            O => \N__10376\,
            I => \N__10291\
        );

    \I__2433\ : InMux
    port map (
            O => \N__10373\,
            I => \N__10288\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__10372\,
            I => \N__10285\
        );

    \I__2431\ : Span4Mux_h
    port map (
            O => \N__10369\,
            I => \N__10282\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__10366\,
            I => \N__10277\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__10361\,
            I => \N__10277\
        );

    \I__2428\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10274\
        );

    \I__2427\ : InMux
    port map (
            O => \N__10355\,
            I => \N__10271\
        );

    \I__2426\ : InMux
    port map (
            O => \N__10352\,
            I => \N__10268\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__10351\,
            I => \N__10265\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__10350\,
            I => \N__10262\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__10347\,
            I => \N__10257\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__10340\,
            I => \N__10257\
        );

    \I__2421\ : InMux
    port map (
            O => \N__10339\,
            I => \N__10252\
        );

    \I__2420\ : InMux
    port map (
            O => \N__10338\,
            I => \N__10252\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__10337\,
            I => \N__10245\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__10336\,
            I => \N__10242\
        );

    \I__2417\ : Span4Mux_v
    port map (
            O => \N__10327\,
            I => \N__10227\
        );

    \I__2416\ : Span4Mux_v
    port map (
            O => \N__10312\,
            I => \N__10227\
        );

    \I__2415\ : Span4Mux_h
    port map (
            O => \N__10309\,
            I => \N__10222\
        );

    \I__2414\ : Span4Mux_v
    port map (
            O => \N__10300\,
            I => \N__10222\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__10297\,
            I => \N__10217\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__10294\,
            I => \N__10217\
        );

    \I__2411\ : Span4Mux_h
    port map (
            O => \N__10291\,
            I => \N__10212\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__10288\,
            I => \N__10212\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10285\,
            I => \N__10209\
        );

    \I__2408\ : Span4Mux_h
    port map (
            O => \N__10282\,
            I => \N__10206\
        );

    \I__2407\ : Span4Mux_v
    port map (
            O => \N__10277\,
            I => \N__10201\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__10274\,
            I => \N__10201\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__10271\,
            I => \N__10196\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10268\,
            I => \N__10196\
        );

    \I__2403\ : InMux
    port map (
            O => \N__10265\,
            I => \N__10193\
        );

    \I__2402\ : InMux
    port map (
            O => \N__10262\,
            I => \N__10190\
        );

    \I__2401\ : Span4Mux_h
    port map (
            O => \N__10257\,
            I => \N__10185\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__10252\,
            I => \N__10185\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10251\,
            I => \N__10176\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10250\,
            I => \N__10176\
        );

    \I__2397\ : InMux
    port map (
            O => \N__10249\,
            I => \N__10176\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10248\,
            I => \N__10176\
        );

    \I__2395\ : InMux
    port map (
            O => \N__10245\,
            I => \N__10171\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10242\,
            I => \N__10171\
        );

    \I__2393\ : CascadeMux
    port map (
            O => \N__10241\,
            I => \N__10167\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__10240\,
            I => \N__10164\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10239\,
            I => \N__10157\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10238\,
            I => \N__10157\
        );

    \I__2389\ : InMux
    port map (
            O => \N__10237\,
            I => \N__10157\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10236\,
            I => \N__10152\
        );

    \I__2387\ : InMux
    port map (
            O => \N__10235\,
            I => \N__10152\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__10234\,
            I => \N__10149\
        );

    \I__2385\ : CascadeMux
    port map (
            O => \N__10233\,
            I => \N__10145\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__10232\,
            I => \N__10142\
        );

    \I__2383\ : Sp12to4
    port map (
            O => \N__10227\,
            I => \N__10137\
        );

    \I__2382\ : Sp12to4
    port map (
            O => \N__10222\,
            I => \N__10137\
        );

    \I__2381\ : Span12Mux_s11_h
    port map (
            O => \N__10217\,
            I => \N__10134\
        );

    \I__2380\ : Sp12to4
    port map (
            O => \N__10212\,
            I => \N__10131\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__10209\,
            I => \N__10128\
        );

    \I__2378\ : Span4Mux_h
    port map (
            O => \N__10206\,
            I => \N__10123\
        );

    \I__2377\ : Span4Mux_v
    port map (
            O => \N__10201\,
            I => \N__10123\
        );

    \I__2376\ : Span4Mux_h
    port map (
            O => \N__10196\,
            I => \N__10116\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__10193\,
            I => \N__10116\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__10190\,
            I => \N__10116\
        );

    \I__2373\ : Span4Mux_v
    port map (
            O => \N__10185\,
            I => \N__10111\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10176\,
            I => \N__10111\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10171\,
            I => \N__10108\
        );

    \I__2370\ : InMux
    port map (
            O => \N__10170\,
            I => \N__10101\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10167\,
            I => \N__10101\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10101\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10157\,
            I => \N__10098\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__10152\,
            I => \N__10095\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10149\,
            I => \N__10088\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10088\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10145\,
            I => \N__10088\
        );

    \I__2362\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10085\
        );

    \I__2361\ : Span12Mux_h
    port map (
            O => \N__10137\,
            I => \N__10082\
        );

    \I__2360\ : Span12Mux_h
    port map (
            O => \N__10134\,
            I => \N__10079\
        );

    \I__2359\ : Span12Mux_s11_v
    port map (
            O => \N__10131\,
            I => \N__10074\
        );

    \I__2358\ : Span12Mux_s11_h
    port map (
            O => \N__10128\,
            I => \N__10074\
        );

    \I__2357\ : Span4Mux_v
    port map (
            O => \N__10123\,
            I => \N__10069\
        );

    \I__2356\ : Span4Mux_v
    port map (
            O => \N__10116\,
            I => \N__10069\
        );

    \I__2355\ : Span4Mux_v
    port map (
            O => \N__10111\,
            I => \N__10062\
        );

    \I__2354\ : Span4Mux_h
    port map (
            O => \N__10108\,
            I => \N__10062\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__10101\,
            I => \N__10062\
        );

    \I__2352\ : Span4Mux_h
    port map (
            O => \N__10098\,
            I => \N__10053\
        );

    \I__2351\ : Span4Mux_v
    port map (
            O => \N__10095\,
            I => \N__10053\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__10088\,
            I => \N__10053\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__10085\,
            I => \N__10053\
        );

    \I__2348\ : Span12Mux_h
    port map (
            O => \N__10082\,
            I => \N__10050\
        );

    \I__2347\ : Span12Mux_v
    port map (
            O => \N__10079\,
            I => \N__10045\
        );

    \I__2346\ : Span12Mux_h
    port map (
            O => \N__10074\,
            I => \N__10045\
        );

    \I__2345\ : Span4Mux_h
    port map (
            O => \N__10069\,
            I => \N__10042\
        );

    \I__2344\ : Span4Mux_v
    port map (
            O => \N__10062\,
            I => \N__10037\
        );

    \I__2343\ : Span4Mux_v
    port map (
            O => \N__10053\,
            I => \N__10037\
        );

    \I__2342\ : Odrv12
    port map (
            O => \N__10050\,
            I => \RnW_c\
        );

    \I__2341\ : Odrv12
    port map (
            O => \N__10045\,
            I => \RnW_c\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__10042\,
            I => \RnW_c\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__10037\,
            I => \RnW_c\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10028\,
            I => \N__10025\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__10025\,
            I => \READ_CYCLE_ACTIVE_rep12_i_ess\
        );

    \I__2336\ : InMux
    port map (
            O => \N__10022\,
            I => \N__10019\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__10019\,
            I => \READ_CYCLE_ACTIVE_rep29_i_ess\
        );

    \I__2334\ : IoInMux
    port map (
            O => \N__10016\,
            I => \N__10013\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__10013\,
            I => \N__10010\
        );

    \I__2332\ : Span4Mux_s3_h
    port map (
            O => \N__10010\,
            I => \N__10007\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__10007\,
            I => \N_195_i\
        );

    \I__2330\ : InMux
    port map (
            O => \N__10004\,
            I => \N__10001\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10001\,
            I => \READ_CYCLE_ACTIVE_rep14_i_ess\
        );

    \I__2328\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9995\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__9995\,
            I => \READ_CYCLE_ACTIVE_rep22_i_ess\
        );

    \I__2326\ : IoInMux
    port map (
            O => \N__9992\,
            I => \N__9989\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__9989\,
            I => \N__9986\
        );

    \I__2324\ : Span4Mux_s3_h
    port map (
            O => \N__9986\,
            I => \N__9983\
        );

    \I__2323\ : Odrv4
    port map (
            O => \N__9983\,
            I => \N_203_i\
        );

    \I__2322\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9977\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__9977\,
            I => \N__9974\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__9974\,
            I => \READ_CYCLE_ACTIVE_rep23_i_ess\
        );

    \I__2319\ : IoInMux
    port map (
            O => \N__9971\,
            I => \N__9968\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__9968\,
            I => \N__9965\
        );

    \I__2317\ : IoSpan4Mux
    port map (
            O => \N__9965\,
            I => \N__9962\
        );

    \I__2316\ : Span4Mux_s3_h
    port map (
            O => \N__9962\,
            I => \N__9959\
        );

    \I__2315\ : Odrv4
    port map (
            O => \N__9959\,
            I => \N_204_i\
        );

    \I__2314\ : InMux
    port map (
            O => \N__9956\,
            I => \N__9953\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__9953\,
            I => \READ_CYCLE_ACTIVE_rep9_i_ess\
        );

    \I__2312\ : IoInMux
    port map (
            O => \N__9950\,
            I => \N__9947\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__9947\,
            I => \N__9944\
        );

    \I__2310\ : Span4Mux_s3_h
    port map (
            O => \N__9944\,
            I => \N__9941\
        );

    \I__2309\ : Span4Mux_v
    port map (
            O => \N__9941\,
            I => \N__9938\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__9938\,
            I => \N_190_i\
        );

    \I__2307\ : InMux
    port map (
            O => \N__9935\,
            I => \N__9932\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__9932\,
            I => \READ_CYCLE_ACTIVE_rep16_i_ess\
        );

    \I__2305\ : InMux
    port map (
            O => \N__9929\,
            I => \N__9926\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__9926\,
            I => \READ_CYCLE_ACTIVE_rep20_i_ess\
        );

    \I__2303\ : IoInMux
    port map (
            O => \N__9923\,
            I => \N__9920\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__9920\,
            I => \N__9917\
        );

    \I__2301\ : Span4Mux_s3_h
    port map (
            O => \N__9917\,
            I => \N__9914\
        );

    \I__2300\ : Odrv4
    port map (
            O => \N__9914\,
            I => \N_201_i\
        );

    \I__2299\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9908\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__9908\,
            I => \READ_CYCLE_ACTIVE_rep8_i_ess\
        );

    \I__2297\ : IoInMux
    port map (
            O => \N__9905\,
            I => \N__9902\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__9902\,
            I => \N__9899\
        );

    \I__2295\ : Odrv12
    port map (
            O => \N__9899\,
            I => \N_189_i\
        );

    \I__2294\ : InMux
    port map (
            O => \N__9896\,
            I => \N__9893\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__9893\,
            I => \READ_CYCLE_ACTIVE_rep21_i_ess\
        );

    \I__2292\ : IoInMux
    port map (
            O => \N__9890\,
            I => \N__9887\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__9887\,
            I => \N__9884\
        );

    \I__2290\ : IoSpan4Mux
    port map (
            O => \N__9884\,
            I => \N__9881\
        );

    \I__2289\ : Span4Mux_s3_h
    port map (
            O => \N__9881\,
            I => \N__9878\
        );

    \I__2288\ : Odrv4
    port map (
            O => \N__9878\,
            I => \N_202_i\
        );

    \I__2287\ : IoInMux
    port map (
            O => \N__9875\,
            I => \N__9872\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__9872\,
            I => \N__9869\
        );

    \I__2285\ : Span12Mux_s11_h
    port map (
            O => \N__9869\,
            I => \N__9866\
        );

    \I__2284\ : Span12Mux_v
    port map (
            O => \N__9866\,
            I => \N__9863\
        );

    \I__2283\ : Odrv12
    port map (
            O => \N__9863\,
            I => \N_210_i\
        );

    \I__2282\ : IoInMux
    port map (
            O => \N__9860\,
            I => \N__9857\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__9857\,
            I => \N__9854\
        );

    \I__2280\ : Odrv12
    port map (
            O => \N__9854\,
            I => \N_191_i\
        );

    \I__2279\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9848\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__9848\,
            I => \READ_CYCLE_ACTIVE_rep10_i_ess\
        );

    \I__2277\ : InMux
    port map (
            O => \N__9845\,
            I => \N__9842\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__9842\,
            I => \READ_CYCLE_ACTIVE_rep26_i_ess\
        );

    \I__2275\ : IoInMux
    port map (
            O => \N__9839\,
            I => \N__9836\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__9836\,
            I => \N__9833\
        );

    \I__2273\ : Span4Mux_s3_h
    port map (
            O => \N__9833\,
            I => \N__9830\
        );

    \I__2272\ : Span4Mux_v
    port map (
            O => \N__9830\,
            I => \N__9827\
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__9827\,
            I => \N_207_i\
        );

    \I__2270\ : InMux
    port map (
            O => \N__9824\,
            I => \N__9821\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__9821\,
            I => \READ_CYCLE_ACTIVE_rep30_i_ess\
        );

    \I__2268\ : InMux
    port map (
            O => \N__9818\,
            I => \N__9815\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__9815\,
            I => \READ_CYCLE_ACTIVE_rep17_i_ess\
        );

    \I__2266\ : IoInMux
    port map (
            O => \N__9812\,
            I => \N__9809\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__9809\,
            I => \N__9806\
        );

    \I__2264\ : Span4Mux_s3_h
    port map (
            O => \N__9806\,
            I => \N__9803\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__9803\,
            I => \N__9800\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__9800\,
            I => \N_198_i\
        );

    \I__2261\ : InMux
    port map (
            O => \N__9797\,
            I => \N__9794\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__9794\,
            I => \READ_CYCLE_ACTIVE_rep18_i_ess\
        );

    \I__2259\ : IoInMux
    port map (
            O => \N__9791\,
            I => \N__9788\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__9788\,
            I => \N__9785\
        );

    \I__2257\ : Span12Mux_s4_h
    port map (
            O => \N__9785\,
            I => \N__9782\
        );

    \I__2256\ : Odrv12
    port map (
            O => \N__9782\,
            I => \N_199_i\
        );

    \I__2255\ : InMux
    port map (
            O => \N__9779\,
            I => \N__9776\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__9776\,
            I => \READ_CYCLE_ACTIVE_rep31_i_ess\
        );

    \I__2253\ : IoInMux
    port map (
            O => \N__9773\,
            I => \N__9770\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__9770\,
            I => \N__9767\
        );

    \I__2251\ : Span4Mux_s3_h
    port map (
            O => \N__9767\,
            I => \N__9764\
        );

    \I__2250\ : Span4Mux_v
    port map (
            O => \N__9764\,
            I => \N__9761\
        );

    \I__2249\ : Odrv4
    port map (
            O => \N__9761\,
            I => \N_212_i\
        );

    \I__2248\ : IoInMux
    port map (
            O => \N__9758\,
            I => \N__9755\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__9755\,
            I => \N__9752\
        );

    \I__2246\ : Span4Mux_s3_h
    port map (
            O => \N__9752\,
            I => \N__9749\
        );

    \I__2245\ : Span4Mux_v
    port map (
            O => \N__9749\,
            I => \N__9746\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__9746\,
            I => \N_197_i\
        );

    \I__2243\ : IoInMux
    port map (
            O => \N__9743\,
            I => \N__9740\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__9740\,
            I => \N__9737\
        );

    \I__2241\ : Span4Mux_s3_h
    port map (
            O => \N__9737\,
            I => \N__9734\
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__9734\,
            I => \N_200_i\
        );

    \I__2239\ : InMux
    port map (
            O => \N__9731\,
            I => \N__9728\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__9728\,
            I => \READ_CYCLE_ACTIVE_rep19_i_ess\
        );

    \I__2237\ : IoInMux
    port map (
            O => \N__9725\,
            I => \N__9722\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__9722\,
            I => \N__9719\
        );

    \I__2235\ : Span4Mux_s3_v
    port map (
            O => \N__9719\,
            I => \N__9716\
        );

    \I__2234\ : Span4Mux_h
    port map (
            O => \N__9716\,
            I => \N__9713\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__9713\,
            I => \N_193_i\
        );

    \I__2232\ : IoInMux
    port map (
            O => \N__9710\,
            I => \N__9707\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9707\,
            I => \N__9704\
        );

    \I__2230\ : Span4Mux_s2_v
    port map (
            O => \N__9704\,
            I => \N__9701\
        );

    \I__2229\ : Span4Mux_v
    port map (
            O => \N__9701\,
            I => \N__9698\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__9698\,
            I => \N_194_i\
        );

    \I__2227\ : IoInMux
    port map (
            O => \N__9695\,
            I => \N__9692\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__9692\,
            I => \N__9689\
        );

    \I__2225\ : Span4Mux_s3_h
    port map (
            O => \N__9689\,
            I => \N__9686\
        );

    \I__2224\ : Span4Mux_v
    port map (
            O => \N__9686\,
            I => \N__9683\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__9683\,
            I => \N_205_i\
        );

    \I__2222\ : IoInMux
    port map (
            O => \N__9680\,
            I => \N__9677\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__9677\,
            I => \N__9674\
        );

    \I__2220\ : IoSpan4Mux
    port map (
            O => \N__9674\,
            I => \N__9671\
        );

    \I__2219\ : Span4Mux_s3_h
    port map (
            O => \N__9671\,
            I => \N__9668\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__9668\,
            I => \N_206_i\
        );

    \I__2217\ : IoInMux
    port map (
            O => \N__9665\,
            I => \N__9662\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__9662\,
            I => \N__9659\
        );

    \I__2215\ : Span4Mux_s3_h
    port map (
            O => \N__9659\,
            I => \N__9656\
        );

    \I__2214\ : Span4Mux_v
    port map (
            O => \N__9656\,
            I => \N__9653\
        );

    \I__2213\ : Odrv4
    port map (
            O => \N__9653\,
            I => \N_208_i\
        );

    \I__2212\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9647\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__9647\,
            I => \READ_CYCLE_ACTIVE_rep25_i_ess\
        );

    \I__2210\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9641\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__9641\,
            I => \READ_CYCLE_ACTIVE_rep24_i_ess\
        );

    \I__2208\ : InMux
    port map (
            O => \N__9638\,
            I => \N__9635\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__9635\,
            I => \READ_CYCLE_ACTIVE_rep27_i_ess\
        );

    \I__2206\ : IoInMux
    port map (
            O => \N__9632\,
            I => \N__9629\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__9629\,
            I => \N__9626\
        );

    \I__2204\ : Span4Mux_s3_h
    port map (
            O => \N__9626\,
            I => \N__9623\
        );

    \I__2203\ : Span4Mux_v
    port map (
            O => \N__9623\,
            I => \N__9620\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__9620\,
            I => \N_211_i\
        );

    \I__2201\ : IoInMux
    port map (
            O => \N__9617\,
            I => \N__9613\
        );

    \I__2200\ : IoInMux
    port map (
            O => \N__9616\,
            I => \N__9610\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__9613\,
            I => \N__9607\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__9610\,
            I => \N__9603\
        );

    \I__2197\ : IoSpan4Mux
    port map (
            O => \N__9607\,
            I => \N__9600\
        );

    \I__2196\ : IoInMux
    port map (
            O => \N__9606\,
            I => \N__9597\
        );

    \I__2195\ : IoSpan4Mux
    port map (
            O => \N__9603\,
            I => \N__9593\
        );

    \I__2194\ : IoSpan4Mux
    port map (
            O => \N__9600\,
            I => \N__9588\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__9597\,
            I => \N__9588\
        );

    \I__2192\ : IoInMux
    port map (
            O => \N__9596\,
            I => \N__9585\
        );

    \I__2191\ : Sp12to4
    port map (
            O => \N__9593\,
            I => \N__9582\
        );

    \I__2190\ : IoSpan4Mux
    port map (
            O => \N__9588\,
            I => \N__9579\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__9585\,
            I => \N__9576\
        );

    \I__2188\ : Span12Mux_s6_h
    port map (
            O => \N__9582\,
            I => \N__9573\
        );

    \I__2187\ : Span4Mux_s3_v
    port map (
            O => \N__9579\,
            I => \N__9570\
        );

    \I__2186\ : IoSpan4Mux
    port map (
            O => \N__9576\,
            I => \N__9567\
        );

    \I__2185\ : Span12Mux_h
    port map (
            O => \N__9573\,
            I => \N__9564\
        );

    \I__2184\ : Sp12to4
    port map (
            O => \N__9570\,
            I => \N__9561\
        );

    \I__2183\ : Span4Mux_s3_h
    port map (
            O => \N__9567\,
            I => \N__9558\
        );

    \I__2182\ : Odrv12
    port map (
            O => \N__9564\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__2181\ : Odrv12
    port map (
            O => \N__9561\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__2180\ : Odrv4
    port map (
            O => \N__9558\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9551\,
            I => \N__9548\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9548\,
            I => \READ_CYCLE_ACTIVE_rep5_i_ess\
        );

    \I__2177\ : IoInMux
    port map (
            O => \N__9545\,
            I => \N__9542\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9542\,
            I => \N__9539\
        );

    \I__2175\ : Span4Mux_s2_v
    port map (
            O => \N__9539\,
            I => \N__9536\
        );

    \I__2174\ : Span4Mux_v
    port map (
            O => \N__9536\,
            I => \N__9533\
        );

    \I__2173\ : Odrv4
    port map (
            O => \N__9533\,
            I => \N_186_i\
        );

    \I__2172\ : InMux
    port map (
            O => \N__9530\,
            I => \N__9527\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9527\,
            I => \READ_CYCLE_ACTIVE_rep6_i_ess\
        );

    \I__2170\ : IoInMux
    port map (
            O => \N__9524\,
            I => \N__9521\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__9521\,
            I => \N__9518\
        );

    \I__2168\ : Span4Mux_s2_v
    port map (
            O => \N__9518\,
            I => \N__9515\
        );

    \I__2167\ : Span4Mux_v
    port map (
            O => \N__9515\,
            I => \N__9512\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__9512\,
            I => \N_187_i\
        );

    \I__2165\ : InMux
    port map (
            O => \N__9509\,
            I => \N__9506\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9506\,
            I => \READ_CYCLE_ACTIVE_rep4_i_ess\
        );

    \I__2163\ : IoInMux
    port map (
            O => \N__9503\,
            I => \N__9500\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__9500\,
            I => \N__9497\
        );

    \I__2161\ : Span4Mux_s2_v
    port map (
            O => \N__9497\,
            I => \N__9494\
        );

    \I__2160\ : Span4Mux_v
    port map (
            O => \N__9494\,
            I => \N__9491\
        );

    \I__2159\ : Odrv4
    port map (
            O => \N__9491\,
            I => \N_185_i\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9485\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9485\,
            I => \READ_CYCLE_ACTIVE_rep2_i_ess\
        );

    \I__2156\ : IoInMux
    port map (
            O => \N__9482\,
            I => \N__9479\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9479\,
            I => \N__9476\
        );

    \I__2154\ : Span4Mux_s2_v
    port map (
            O => \N__9476\,
            I => \N__9473\
        );

    \I__2153\ : Span4Mux_v
    port map (
            O => \N__9473\,
            I => \N__9470\
        );

    \I__2152\ : Odrv4
    port map (
            O => \N__9470\,
            I => \N_183_i\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9467\,
            I => \N__9464\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__9464\,
            I => \READ_CYCLE_ACTIVE_rep0_i_ess\
        );

    \I__2149\ : IoInMux
    port map (
            O => \N__9461\,
            I => \N__9458\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__2147\ : Span4Mux_s0_v
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__2146\ : Span4Mux_v
    port map (
            O => \N__9452\,
            I => \N__9449\
        );

    \I__2145\ : Span4Mux_v
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__2144\ : Odrv4
    port map (
            O => \N__9446\,
            I => \N_181_i\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9443\,
            I => \N__9440\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9440\,
            I => \READ_CYCLE_ACTIVE_rep7_i_ess\
        );

    \I__2141\ : IoInMux
    port map (
            O => \N__9437\,
            I => \N__9434\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__9434\,
            I => \N__9431\
        );

    \I__2139\ : Span4Mux_s2_v
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__2138\ : Span4Mux_v
    port map (
            O => \N__9428\,
            I => \N__9425\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__9425\,
            I => \N_188_i\
        );

    \I__2136\ : IoInMux
    port map (
            O => \N__9422\,
            I => \N__9419\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__9419\,
            I => \N__9416\
        );

    \I__2134\ : IoSpan4Mux
    port map (
            O => \N__9416\,
            I => \N__9413\
        );

    \I__2133\ : IoSpan4Mux
    port map (
            O => \N__9413\,
            I => \N__9410\
        );

    \I__2132\ : Span4Mux_s2_h
    port map (
            O => \N__9410\,
            I => \N__9407\
        );

    \I__2131\ : Odrv4
    port map (
            O => \N__9407\,
            I => \N_209_i\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9404\,
            I => \N__9401\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__9401\,
            I => \READ_CYCLE_ACTIVE_rep28_i_ess\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9395\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__9395\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9388\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9385\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9388\,
            I => \N__9381\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__9385\,
            I => \N__9378\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9384\,
            I => \N__9375\
        );

    \I__2121\ : Span4Mux_v
    port map (
            O => \N__9381\,
            I => \N__9372\
        );

    \I__2120\ : Span4Mux_h
    port map (
            O => \N__9378\,
            I => \N__9367\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__9375\,
            I => \N__9367\
        );

    \I__2118\ : Span4Mux_v
    port map (
            O => \N__9372\,
            I => \N__9362\
        );

    \I__2117\ : Span4Mux_h
    port map (
            O => \N__9367\,
            I => \N__9362\
        );

    \I__2116\ : Span4Mux_v
    port map (
            O => \N__9362\,
            I => \N__9359\
        );

    \I__2115\ : Sp12to4
    port map (
            O => \N__9359\,
            I => \N__9356\
        );

    \I__2114\ : Span12Mux_h
    port map (
            O => \N__9356\,
            I => \N__9353\
        );

    \I__2113\ : Odrv12
    port map (
            O => \N__9353\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__2112\ : IoInMux
    port map (
            O => \N__9350\,
            I => \N__9347\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__9347\,
            I => \N__9344\
        );

    \I__2110\ : Span12Mux_s6_h
    port map (
            O => \N__9344\,
            I => \N__9341\
        );

    \I__2109\ : Odrv12
    port map (
            O => \N__9341\,
            I => \un1_D_UM_AMIGA_2\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9335\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__9335\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9329\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__9329\,
            I => \N__9325\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9322\
        );

    \I__2103\ : Span4Mux_v
    port map (
            O => \N__9325\,
            I => \N__9318\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__9322\,
            I => \N__9315\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9321\,
            I => \N__9312\
        );

    \I__2100\ : Span4Mux_v
    port map (
            O => \N__9318\,
            I => \N__9309\
        );

    \I__2099\ : Span4Mux_v
    port map (
            O => \N__9315\,
            I => \N__9306\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__9312\,
            I => \N__9303\
        );

    \I__2097\ : Sp12to4
    port map (
            O => \N__9309\,
            I => \N__9296\
        );

    \I__2096\ : Sp12to4
    port map (
            O => \N__9306\,
            I => \N__9296\
        );

    \I__2095\ : Span12Mux_v
    port map (
            O => \N__9303\,
            I => \N__9296\
        );

    \I__2094\ : Span12Mux_h
    port map (
            O => \N__9296\,
            I => \N__9293\
        );

    \I__2093\ : Span12Mux_v
    port map (
            O => \N__9293\,
            I => \N__9290\
        );

    \I__2092\ : Odrv12
    port map (
            O => \N__9290\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__2091\ : IoInMux
    port map (
            O => \N__9287\,
            I => \N__9284\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9284\,
            I => \N__9281\
        );

    \I__2089\ : IoSpan4Mux
    port map (
            O => \N__9281\,
            I => \N__9278\
        );

    \I__2088\ : Span4Mux_s2_h
    port map (
            O => \N__9278\,
            I => \N__9275\
        );

    \I__2087\ : Sp12to4
    port map (
            O => \N__9275\,
            I => \N__9272\
        );

    \I__2086\ : Odrv12
    port map (
            O => \N__9272\,
            I => \un1_D_UM_AMIGA_6\
        );

    \I__2085\ : IoInMux
    port map (
            O => \N__9269\,
            I => \N__9265\
        );

    \I__2084\ : InMux
    port map (
            O => \N__9268\,
            I => \N__9262\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__9265\,
            I => \N__9259\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__9262\,
            I => \N__9256\
        );

    \I__2081\ : Span4Mux_s2_h
    port map (
            O => \N__9259\,
            I => \N__9253\
        );

    \I__2080\ : Sp12to4
    port map (
            O => \N__9256\,
            I => \N__9250\
        );

    \I__2079\ : Span4Mux_v
    port map (
            O => \N__9253\,
            I => \N__9247\
        );

    \I__2078\ : Span12Mux_v
    port map (
            O => \N__9250\,
            I => \N__9244\
        );

    \I__2077\ : Sp12to4
    port map (
            O => \N__9247\,
            I => \N__9241\
        );

    \I__2076\ : Span12Mux_v
    port map (
            O => \N__9244\,
            I => \N__9238\
        );

    \I__2075\ : Span12Mux_h
    port map (
            O => \N__9241\,
            I => \N__9235\
        );

    \I__2074\ : Span12Mux_h
    port map (
            O => \N__9238\,
            I => \N__9232\
        );

    \I__2073\ : Span12Mux_h
    port map (
            O => \N__9235\,
            I => \N__9229\
        );

    \I__2072\ : Odrv12
    port map (
            O => \N__9232\,
            I => \D_LL_040_in_4\
        );

    \I__2071\ : Odrv12
    port map (
            O => \N__9229\,
            I => \D_LL_040_in_4\
        );

    \I__2070\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9221\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__9221\,
            I => \N__9218\
        );

    \I__2068\ : Span4Mux_v
    port map (
            O => \N__9218\,
            I => \N__9215\
        );

    \I__2067\ : Sp12to4
    port map (
            O => \N__9215\,
            I => \N__9212\
        );

    \I__2066\ : Span12Mux_h
    port map (
            O => \N__9212\,
            I => \N__9209\
        );

    \I__2065\ : Odrv12
    port map (
            O => \N__9209\,
            I => \D_UM_040_in_4\
        );

    \I__2064\ : IoInMux
    port map (
            O => \N__9206\,
            I => \N__9203\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__2062\ : IoSpan4Mux
    port map (
            O => \N__9200\,
            I => \N__9197\
        );

    \I__2061\ : Span4Mux_s3_h
    port map (
            O => \N__9197\,
            I => \N__9194\
        );

    \I__2060\ : Span4Mux_h
    port map (
            O => \N__9194\,
            I => \N__9191\
        );

    \I__2059\ : Span4Mux_h
    port map (
            O => \N__9191\,
            I => \N__9188\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__9188\,
            I => \N__9185\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__9185\,
            I => \un1_D_UM_040_4\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9179\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__9179\,
            I => \N__9176\
        );

    \I__2054\ : Span4Mux_v
    port map (
            O => \N__9176\,
            I => \N__9173\
        );

    \I__2053\ : Span4Mux_h
    port map (
            O => \N__9173\,
            I => \N__9170\
        );

    \I__2052\ : Span4Mux_h
    port map (
            O => \N__9170\,
            I => \N__9167\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__9167\,
            I => \D_UU_040_in_4\
        );

    \I__2050\ : IoInMux
    port map (
            O => \N__9164\,
            I => \N__9161\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9161\,
            I => \N__9158\
        );

    \I__2048\ : Span4Mux_s1_h
    port map (
            O => \N__9158\,
            I => \N__9155\
        );

    \I__2047\ : Sp12to4
    port map (
            O => \N__9155\,
            I => \N__9151\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9154\,
            I => \N__9148\
        );

    \I__2045\ : Span12Mux_v
    port map (
            O => \N__9151\,
            I => \N__9145\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__9148\,
            I => \N__9142\
        );

    \I__2043\ : Span12Mux_h
    port map (
            O => \N__9145\,
            I => \N__9139\
        );

    \I__2042\ : Span12Mux_h
    port map (
            O => \N__9142\,
            I => \N__9136\
        );

    \I__2041\ : Span12Mux_h
    port map (
            O => \N__9139\,
            I => \N__9131\
        );

    \I__2040\ : Span12Mux_v
    port map (
            O => \N__9136\,
            I => \N__9131\
        );

    \I__2039\ : Odrv12
    port map (
            O => \N__9131\,
            I => \D_LM_040_in_4\
        );

    \I__2038\ : IoInMux
    port map (
            O => \N__9128\,
            I => \N__9125\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__9125\,
            I => \N__9122\
        );

    \I__2036\ : IoSpan4Mux
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__2035\ : Sp12to4
    port map (
            O => \N__9119\,
            I => \N__9116\
        );

    \I__2034\ : Span12Mux_s6_v
    port map (
            O => \N__9116\,
            I => \N__9113\
        );

    \I__2033\ : Odrv12
    port map (
            O => \N__9113\,
            I => \un1_D_UU_040_4\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9110\,
            I => \N__9097\
        );

    \I__2031\ : InMux
    port map (
            O => \N__9109\,
            I => \N__9097\
        );

    \I__2030\ : InMux
    port map (
            O => \N__9108\,
            I => \N__9097\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9107\,
            I => \N__9092\
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__9106\,
            I => \N__9086\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9105\,
            I => \N__9080\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9104\,
            I => \N__9080\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__9097\,
            I => \N__9077\
        );

    \I__2024\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9074\
        );

    \I__2023\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9071\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__9092\,
            I => \N__9068\
        );

    \I__2021\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9063\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9063\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9056\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9056\
        );

    \I__2017\ : InMux
    port map (
            O => \N__9085\,
            I => \N__9056\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9080\,
            I => \N__9053\
        );

    \I__2015\ : Span4Mux_h
    port map (
            O => \N__9077\,
            I => \N__9046\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__9074\,
            I => \N__9046\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__9071\,
            I => \N__9043\
        );

    \I__2012\ : Span4Mux_h
    port map (
            O => \N__9068\,
            I => \N__9038\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__9063\,
            I => \N__9038\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__9056\,
            I => \N__9033\
        );

    \I__2009\ : Span4Mux_h
    port map (
            O => \N__9053\,
            I => \N__9033\
        );

    \I__2008\ : InMux
    port map (
            O => \N__9052\,
            I => \N__9030\
        );

    \I__2007\ : InMux
    port map (
            O => \N__9051\,
            I => \N__9027\
        );

    \I__2006\ : Span4Mux_v
    port map (
            O => \N__9046\,
            I => \N__9022\
        );

    \I__2005\ : Sp12to4
    port map (
            O => \N__9043\,
            I => \N__9011\
        );

    \I__2004\ : Sp12to4
    port map (
            O => \N__9038\,
            I => \N__9011\
        );

    \I__2003\ : Sp12to4
    port map (
            O => \N__9033\,
            I => \N__9011\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9030\,
            I => \N__9011\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__9027\,
            I => \N__9011\
        );

    \I__2000\ : InMux
    port map (
            O => \N__9026\,
            I => \N__9008\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__9025\,
            I => \N__9005\
        );

    \I__1998\ : Span4Mux_v
    port map (
            O => \N__9022\,
            I => \N__9002\
        );

    \I__1997\ : Span12Mux_v
    port map (
            O => \N__9011\,
            I => \N__8999\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__9008\,
            I => \N__8996\
        );

    \I__1995\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8993\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__9002\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1993\ : Odrv12
    port map (
            O => \N__8999\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1992\ : Odrv12
    port map (
            O => \N__8996\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__8993\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1990\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__8981\,
            I => \N__8978\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__8978\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\
        );

    \I__1987\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8972\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__8972\,
            I => \N__8968\
        );

    \I__1985\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8964\
        );

    \I__1984\ : Span4Mux_v
    port map (
            O => \N__8968\,
            I => \N__8961\
        );

    \I__1983\ : InMux
    port map (
            O => \N__8967\,
            I => \N__8958\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__8964\,
            I => \N__8955\
        );

    \I__1981\ : Span4Mux_v
    port map (
            O => \N__8961\,
            I => \N__8952\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__8958\,
            I => \N__8949\
        );

    \I__1979\ : Span4Mux_v
    port map (
            O => \N__8955\,
            I => \N__8946\
        );

    \I__1978\ : Span4Mux_v
    port map (
            O => \N__8952\,
            I => \N__8943\
        );

    \I__1977\ : Span4Mux_v
    port map (
            O => \N__8949\,
            I => \N__8940\
        );

    \I__1976\ : Sp12to4
    port map (
            O => \N__8946\,
            I => \N__8933\
        );

    \I__1975\ : Sp12to4
    port map (
            O => \N__8943\,
            I => \N__8933\
        );

    \I__1974\ : Sp12to4
    port map (
            O => \N__8940\,
            I => \N__8933\
        );

    \I__1973\ : Span12Mux_h
    port map (
            O => \N__8933\,
            I => \N__8930\
        );

    \I__1972\ : Odrv12
    port map (
            O => \N__8930\,
            I => \D_UM_AMIGA_in_0\
        );

    \I__1971\ : IoInMux
    port map (
            O => \N__8927\,
            I => \N__8924\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__1969\ : Span12Mux_s8_h
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__1968\ : Odrv12
    port map (
            O => \N__8918\,
            I => \un1_D_UM_AMIGA_0\
        );

    \I__1967\ : InMux
    port map (
            O => \N__8915\,
            I => \N__8912\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__8912\,
            I => \N__8909\
        );

    \I__1965\ : Span4Mux_v
    port map (
            O => \N__8909\,
            I => \N__8906\
        );

    \I__1964\ : Span4Mux_v
    port map (
            O => \N__8906\,
            I => \N__8903\
        );

    \I__1963\ : Sp12to4
    port map (
            O => \N__8903\,
            I => \N__8900\
        );

    \I__1962\ : Span12Mux_h
    port map (
            O => \N__8900\,
            I => \N__8897\
        );

    \I__1961\ : Odrv12
    port map (
            O => \N__8897\,
            I => \D_UM_040_in_7\
        );

    \I__1960\ : IoInMux
    port map (
            O => \N__8894\,
            I => \N__8891\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__8891\,
            I => \N__8887\
        );

    \I__1958\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8884\
        );

    \I__1957\ : IoSpan4Mux
    port map (
            O => \N__8887\,
            I => \N__8881\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__8884\,
            I => \N__8878\
        );

    \I__1955\ : Span4Mux_s3_h
    port map (
            O => \N__8881\,
            I => \N__8875\
        );

    \I__1954\ : Span4Mux_h
    port map (
            O => \N__8878\,
            I => \N__8872\
        );

    \I__1953\ : Sp12to4
    port map (
            O => \N__8875\,
            I => \N__8869\
        );

    \I__1952\ : Sp12to4
    port map (
            O => \N__8872\,
            I => \N__8866\
        );

    \I__1951\ : Span12Mux_v
    port map (
            O => \N__8869\,
            I => \N__8863\
        );

    \I__1950\ : Span12Mux_v
    port map (
            O => \N__8866\,
            I => \N__8860\
        );

    \I__1949\ : Span12Mux_h
    port map (
            O => \N__8863\,
            I => \N__8857\
        );

    \I__1948\ : Span12Mux_v
    port map (
            O => \N__8860\,
            I => \N__8854\
        );

    \I__1947\ : Span12Mux_h
    port map (
            O => \N__8857\,
            I => \N__8851\
        );

    \I__1946\ : Span12Mux_h
    port map (
            O => \N__8854\,
            I => \N__8848\
        );

    \I__1945\ : Odrv12
    port map (
            O => \N__8851\,
            I => \D_LL_040_in_7\
        );

    \I__1944\ : Odrv12
    port map (
            O => \N__8848\,
            I => \D_LL_040_in_7\
        );

    \I__1943\ : IoInMux
    port map (
            O => \N__8843\,
            I => \N__8840\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__8840\,
            I => \N__8837\
        );

    \I__1941\ : Span12Mux_s5_h
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__1940\ : Span12Mux_h
    port map (
            O => \N__8834\,
            I => \N__8831\
        );

    \I__1939\ : Odrv12
    port map (
            O => \N__8831\,
            I => \un1_D_UM_040_7\
        );

    \I__1938\ : InMux
    port map (
            O => \N__8828\,
            I => \N__8824\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8827\,
            I => \N__8818\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8824\,
            I => \N__8812\
        );

    \I__1935\ : InMux
    port map (
            O => \N__8823\,
            I => \N__8809\
        );

    \I__1934\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8804\
        );

    \I__1933\ : InMux
    port map (
            O => \N__8821\,
            I => \N__8801\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__8818\,
            I => \N__8793\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8817\,
            I => \N__8788\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8785\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8815\,
            I => \N__8782\
        );

    \I__1928\ : Span4Mux_h
    port map (
            O => \N__8812\,
            I => \N__8776\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__8809\,
            I => \N__8776\
        );

    \I__1926\ : InMux
    port map (
            O => \N__8808\,
            I => \N__8773\
        );

    \I__1925\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8770\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8804\,
            I => \N__8763\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__8801\,
            I => \N__8763\
        );

    \I__1922\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8758\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8799\,
            I => \N__8758\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8798\,
            I => \N__8751\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8797\,
            I => \N__8751\
        );

    \I__1918\ : InMux
    port map (
            O => \N__8796\,
            I => \N__8748\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__8793\,
            I => \N__8742\
        );

    \I__1916\ : InMux
    port map (
            O => \N__8792\,
            I => \N__8736\
        );

    \I__1915\ : InMux
    port map (
            O => \N__8791\,
            I => \N__8736\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__8788\,
            I => \N__8731\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__8785\,
            I => \N__8728\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__8782\,
            I => \N__8725\
        );

    \I__1911\ : InMux
    port map (
            O => \N__8781\,
            I => \N__8722\
        );

    \I__1910\ : Span4Mux_h
    port map (
            O => \N__8776\,
            I => \N__8714\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__8773\,
            I => \N__8714\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8770\,
            I => \N__8714\
        );

    \I__1907\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8711\
        );

    \I__1906\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8707\
        );

    \I__1905\ : Span4Mux_h
    port map (
            O => \N__8763\,
            I => \N__8702\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8758\,
            I => \N__8702\
        );

    \I__1903\ : InMux
    port map (
            O => \N__8757\,
            I => \N__8699\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8696\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__8751\,
            I => \N__8691\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__8748\,
            I => \N__8691\
        );

    \I__1899\ : InMux
    port map (
            O => \N__8747\,
            I => \N__8688\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8746\,
            I => \N__8685\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8745\,
            I => \N__8682\
        );

    \I__1896\ : Span4Mux_v
    port map (
            O => \N__8742\,
            I => \N__8679\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8676\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__8736\,
            I => \N__8673\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8735\,
            I => \N__8670\
        );

    \I__1892\ : InMux
    port map (
            O => \N__8734\,
            I => \N__8667\
        );

    \I__1891\ : Span4Mux_h
    port map (
            O => \N__8731\,
            I => \N__8657\
        );

    \I__1890\ : Span4Mux_h
    port map (
            O => \N__8728\,
            I => \N__8657\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__8725\,
            I => \N__8657\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8722\,
            I => \N__8657\
        );

    \I__1887\ : InMux
    port map (
            O => \N__8721\,
            I => \N__8654\
        );

    \I__1886\ : Span4Mux_v
    port map (
            O => \N__8714\,
            I => \N__8649\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8711\,
            I => \N__8649\
        );

    \I__1884\ : InMux
    port map (
            O => \N__8710\,
            I => \N__8646\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__8707\,
            I => \N__8642\
        );

    \I__1882\ : Sp12to4
    port map (
            O => \N__8702\,
            I => \N__8637\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__8699\,
            I => \N__8637\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__8696\,
            I => \N__8634\
        );

    \I__1879\ : Span4Mux_v
    port map (
            O => \N__8691\,
            I => \N__8625\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8688\,
            I => \N__8625\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8685\,
            I => \N__8625\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8682\,
            I => \N__8625\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__8679\,
            I => \N__8616\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__8676\,
            I => \N__8616\
        );

    \I__1873\ : Span4Mux_v
    port map (
            O => \N__8673\,
            I => \N__8616\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8670\,
            I => \N__8616\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8667\,
            I => \N__8613\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8610\
        );

    \I__1869\ : Span4Mux_v
    port map (
            O => \N__8657\,
            I => \N__8605\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8654\,
            I => \N__8605\
        );

    \I__1867\ : Span4Mux_h
    port map (
            O => \N__8649\,
            I => \N__8600\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__8646\,
            I => \N__8600\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8597\
        );

    \I__1864\ : Span12Mux_v
    port map (
            O => \N__8642\,
            I => \N__8593\
        );

    \I__1863\ : Span12Mux_v
    port map (
            O => \N__8637\,
            I => \N__8588\
        );

    \I__1862\ : Span12Mux_v
    port map (
            O => \N__8634\,
            I => \N__8588\
        );

    \I__1861\ : Span4Mux_v
    port map (
            O => \N__8625\,
            I => \N__8583\
        );

    \I__1860\ : Span4Mux_h
    port map (
            O => \N__8616\,
            I => \N__8583\
        );

    \I__1859\ : Span12Mux_s9_v
    port map (
            O => \N__8613\,
            I => \N__8578\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__8610\,
            I => \N__8578\
        );

    \I__1857\ : Span4Mux_v
    port map (
            O => \N__8605\,
            I => \N__8571\
        );

    \I__1856\ : Span4Mux_v
    port map (
            O => \N__8600\,
            I => \N__8571\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__8597\,
            I => \N__8571\
        );

    \I__1854\ : InMux
    port map (
            O => \N__8596\,
            I => \N__8568\
        );

    \I__1853\ : Odrv12
    port map (
            O => \N__8593\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1852\ : Odrv12
    port map (
            O => \N__8588\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__8583\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1850\ : Odrv12
    port map (
            O => \N__8578\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__8571\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8568\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8555\,
            I => \N__8552\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__8552\,
            I => \N__8549\
        );

    \I__1845\ : Span4Mux_v
    port map (
            O => \N__8549\,
            I => \N__8546\
        );

    \I__1844\ : Sp12to4
    port map (
            O => \N__8546\,
            I => \N__8543\
        );

    \I__1843\ : Span12Mux_h
    port map (
            O => \N__8543\,
            I => \N__8540\
        );

    \I__1842\ : Odrv12
    port map (
            O => \N__8540\,
            I => \D_UU_040_in_7\
        );

    \I__1841\ : IoInMux
    port map (
            O => \N__8537\,
            I => \N__8534\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__1839\ : IoSpan4Mux
    port map (
            O => \N__8531\,
            I => \N__8528\
        );

    \I__1838\ : Span4Mux_s2_h
    port map (
            O => \N__8528\,
            I => \N__8524\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8521\
        );

    \I__1836\ : Sp12to4
    port map (
            O => \N__8524\,
            I => \N__8518\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8521\,
            I => \N__8515\
        );

    \I__1834\ : Span12Mux_h
    port map (
            O => \N__8518\,
            I => \N__8512\
        );

    \I__1833\ : Span12Mux_s9_v
    port map (
            O => \N__8515\,
            I => \N__8509\
        );

    \I__1832\ : Span12Mux_h
    port map (
            O => \N__8512\,
            I => \N__8506\
        );

    \I__1831\ : Span12Mux_h
    port map (
            O => \N__8509\,
            I => \N__8503\
        );

    \I__1830\ : Odrv12
    port map (
            O => \N__8506\,
            I => \D_LM_040_in_7\
        );

    \I__1829\ : Odrv12
    port map (
            O => \N__8503\,
            I => \D_LM_040_in_7\
        );

    \I__1828\ : IoInMux
    port map (
            O => \N__8498\,
            I => \N__8495\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8495\,
            I => \N__8492\
        );

    \I__1826\ : IoSpan4Mux
    port map (
            O => \N__8492\,
            I => \N__8489\
        );

    \I__1825\ : Span4Mux_s3_v
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__1824\ : Span4Mux_h
    port map (
            O => \N__8486\,
            I => \N__8483\
        );

    \I__1823\ : Span4Mux_h
    port map (
            O => \N__8483\,
            I => \N__8480\
        );

    \I__1822\ : Span4Mux_h
    port map (
            O => \N__8480\,
            I => \N__8477\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__8477\,
            I => \un1_D_UU_040_7\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8471\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8471\,
            I => \N__8468\
        );

    \I__1818\ : Odrv12
    port map (
            O => \N__8468\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8461\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8464\,
            I => \N__8458\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__8461\,
            I => \N__8454\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8458\,
            I => \N__8451\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8457\,
            I => \N__8448\
        );

    \I__1812\ : Span4Mux_v
    port map (
            O => \N__8454\,
            I => \N__8445\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__8451\,
            I => \N__8440\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8448\,
            I => \N__8440\
        );

    \I__1809\ : Span4Mux_v
    port map (
            O => \N__8445\,
            I => \N__8437\
        );

    \I__1808\ : Span4Mux_v
    port map (
            O => \N__8440\,
            I => \N__8434\
        );

    \I__1807\ : Sp12to4
    port map (
            O => \N__8437\,
            I => \N__8431\
        );

    \I__1806\ : Span4Mux_v
    port map (
            O => \N__8434\,
            I => \N__8428\
        );

    \I__1805\ : Span12Mux_h
    port map (
            O => \N__8431\,
            I => \N__8425\
        );

    \I__1804\ : Sp12to4
    port map (
            O => \N__8428\,
            I => \N__8422\
        );

    \I__1803\ : Span12Mux_v
    port map (
            O => \N__8425\,
            I => \N__8417\
        );

    \I__1802\ : Span12Mux_h
    port map (
            O => \N__8422\,
            I => \N__8417\
        );

    \I__1801\ : Odrv12
    port map (
            O => \N__8417\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__1800\ : IoInMux
    port map (
            O => \N__8414\,
            I => \N__8411\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8411\,
            I => \N__8408\
        );

    \I__1798\ : IoSpan4Mux
    port map (
            O => \N__8408\,
            I => \N__8405\
        );

    \I__1797\ : Span4Mux_s2_v
    port map (
            O => \N__8405\,
            I => \N__8402\
        );

    \I__1796\ : Sp12to4
    port map (
            O => \N__8402\,
            I => \N__8399\
        );

    \I__1795\ : Span12Mux_s10_v
    port map (
            O => \N__8399\,
            I => \N__8396\
        );

    \I__1794\ : Odrv12
    port map (
            O => \N__8396\,
            I => \un1_D_UM_AMIGA_4\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__8390\,
            I => \N__8387\
        );

    \I__1791\ : Span4Mux_v
    port map (
            O => \N__8387\,
            I => \N__8384\
        );

    \I__1790\ : Sp12to4
    port map (
            O => \N__8384\,
            I => \N__8381\
        );

    \I__1789\ : Span12Mux_h
    port map (
            O => \N__8381\,
            I => \N__8378\
        );

    \I__1788\ : Odrv12
    port map (
            O => \N__8378\,
            I => \D_LM_AMIGA_in_7\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8375\,
            I => \N__8372\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8372\,
            I => \N__8367\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8371\,
            I => \N__8364\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8361\
        );

    \I__1783\ : Sp12to4
    port map (
            O => \N__8367\,
            I => \N__8358\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8364\,
            I => \N__8353\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__8361\,
            I => \N__8353\
        );

    \I__1780\ : Span12Mux_h
    port map (
            O => \N__8358\,
            I => \N__8350\
        );

    \I__1779\ : Span12Mux_v
    port map (
            O => \N__8353\,
            I => \N__8347\
        );

    \I__1778\ : Span12Mux_v
    port map (
            O => \N__8350\,
            I => \N__8342\
        );

    \I__1777\ : Span12Mux_h
    port map (
            O => \N__8347\,
            I => \N__8342\
        );

    \I__1776\ : Odrv12
    port map (
            O => \N__8342\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__1775\ : IoInMux
    port map (
            O => \N__8339\,
            I => \N__8336\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__8336\,
            I => \N__8333\
        );

    \I__1773\ : Span12Mux_s7_h
    port map (
            O => \N__8333\,
            I => \N__8330\
        );

    \I__1772\ : Odrv12
    port map (
            O => \N__8330\,
            I => \un2_D_LM_AMIGA_7\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8327\,
            I => \N__8324\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8324\,
            I => \N__8321\
        );

    \I__1769\ : Odrv12
    port map (
            O => \N__8321\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\
        );

    \I__1768\ : InMux
    port map (
            O => \N__8318\,
            I => \N__8315\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__8315\,
            I => \N__8312\
        );

    \I__1766\ : Span4Mux_v
    port map (
            O => \N__8312\,
            I => \N__8307\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8311\,
            I => \N__8304\
        );

    \I__1764\ : InMux
    port map (
            O => \N__8310\,
            I => \N__8301\
        );

    \I__1763\ : Sp12to4
    port map (
            O => \N__8307\,
            I => \N__8296\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__8304\,
            I => \N__8296\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8301\,
            I => \N__8293\
        );

    \I__1760\ : Span12Mux_h
    port map (
            O => \N__8296\,
            I => \N__8290\
        );

    \I__1759\ : Span12Mux_v
    port map (
            O => \N__8293\,
            I => \N__8287\
        );

    \I__1758\ : Span12Mux_v
    port map (
            O => \N__8290\,
            I => \N__8284\
        );

    \I__1757\ : Span12Mux_h
    port map (
            O => \N__8287\,
            I => \N__8281\
        );

    \I__1756\ : Odrv12
    port map (
            O => \N__8284\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1755\ : Odrv12
    port map (
            O => \N__8281\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1754\ : IoInMux
    port map (
            O => \N__8276\,
            I => \N__8273\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__8273\,
            I => \N__8270\
        );

    \I__1752\ : Span12Mux_s4_h
    port map (
            O => \N__8270\,
            I => \N__8267\
        );

    \I__1751\ : Span12Mux_h
    port map (
            O => \N__8267\,
            I => \N__8264\
        );

    \I__1750\ : Odrv12
    port map (
            O => \N__8264\,
            I => \un1_D_UM_AMIGA_7\
        );

    \I__1749\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8257\
        );

    \I__1748\ : InMux
    port map (
            O => \N__8260\,
            I => \N__8253\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8257\,
            I => \N__8250\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8256\,
            I => \N__8247\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8253\,
            I => \N__8244\
        );

    \I__1744\ : Sp12to4
    port map (
            O => \N__8250\,
            I => \N__8241\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8247\,
            I => \N__8238\
        );

    \I__1742\ : Span4Mux_v
    port map (
            O => \N__8244\,
            I => \N__8235\
        );

    \I__1741\ : Span12Mux_v
    port map (
            O => \N__8241\,
            I => \N__8232\
        );

    \I__1740\ : Span12Mux_h
    port map (
            O => \N__8238\,
            I => \N__8229\
        );

    \I__1739\ : Sp12to4
    port map (
            O => \N__8235\,
            I => \N__8226\
        );

    \I__1738\ : Span12Mux_h
    port map (
            O => \N__8232\,
            I => \N__8223\
        );

    \I__1737\ : Span12Mux_v
    port map (
            O => \N__8229\,
            I => \N__8218\
        );

    \I__1736\ : Span12Mux_h
    port map (
            O => \N__8226\,
            I => \N__8218\
        );

    \I__1735\ : Odrv12
    port map (
            O => \N__8223\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1734\ : Odrv12
    port map (
            O => \N__8218\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1733\ : InMux
    port map (
            O => \N__8213\,
            I => \N__8210\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__8210\,
            I => \N__8207\
        );

    \I__1731\ : Span12Mux_s8_v
    port map (
            O => \N__8207\,
            I => \N__8204\
        );

    \I__1730\ : Odrv12
    port map (
            O => \N__8204\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\
        );

    \I__1729\ : IoInMux
    port map (
            O => \N__8201\,
            I => \N__8198\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__8198\,
            I => \N__8195\
        );

    \I__1727\ : IoSpan4Mux
    port map (
            O => \N__8195\,
            I => \N__8192\
        );

    \I__1726\ : IoSpan4Mux
    port map (
            O => \N__8192\,
            I => \N__8189\
        );

    \I__1725\ : IoSpan4Mux
    port map (
            O => \N__8189\,
            I => \N__8186\
        );

    \I__1724\ : Span4Mux_s2_v
    port map (
            O => \N__8186\,
            I => \N__8183\
        );

    \I__1723\ : Span4Mux_v
    port map (
            O => \N__8183\,
            I => \N__8180\
        );

    \I__1722\ : Odrv4
    port map (
            O => \N__8180\,
            I => \un1_D_UM_AMIGA_5\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8177\,
            I => \N__8174\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8174\,
            I => \N__8171\
        );

    \I__1719\ : Span4Mux_v
    port map (
            O => \N__8171\,
            I => \N__8168\
        );

    \I__1718\ : Sp12to4
    port map (
            O => \N__8168\,
            I => \N__8165\
        );

    \I__1717\ : Span12Mux_h
    port map (
            O => \N__8165\,
            I => \N__8162\
        );

    \I__1716\ : Odrv12
    port map (
            O => \N__8162\,
            I => \D_UU_040_in_2\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8159\,
            I => \N__8156\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8156\,
            I => \N__8152\
        );

    \I__1713\ : IoInMux
    port map (
            O => \N__8155\,
            I => \N__8149\
        );

    \I__1712\ : Span4Mux_h
    port map (
            O => \N__8152\,
            I => \N__8146\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8149\,
            I => \N__8143\
        );

    \I__1710\ : Sp12to4
    port map (
            O => \N__8146\,
            I => \N__8140\
        );

    \I__1709\ : Span12Mux_s9_h
    port map (
            O => \N__8143\,
            I => \N__8137\
        );

    \I__1708\ : Span12Mux_v
    port map (
            O => \N__8140\,
            I => \N__8134\
        );

    \I__1707\ : Span12Mux_h
    port map (
            O => \N__8137\,
            I => \N__8131\
        );

    \I__1706\ : Span12Mux_v
    port map (
            O => \N__8134\,
            I => \N__8128\
        );

    \I__1705\ : Span12Mux_v
    port map (
            O => \N__8131\,
            I => \N__8125\
        );

    \I__1704\ : Span12Mux_h
    port map (
            O => \N__8128\,
            I => \N__8122\
        );

    \I__1703\ : Odrv12
    port map (
            O => \N__8125\,
            I => \D_LM_040_in_2\
        );

    \I__1702\ : Odrv12
    port map (
            O => \N__8122\,
            I => \D_LM_040_in_2\
        );

    \I__1701\ : IoInMux
    port map (
            O => \N__8117\,
            I => \N__8114\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8114\,
            I => \N__8111\
        );

    \I__1699\ : IoSpan4Mux
    port map (
            O => \N__8111\,
            I => \N__8108\
        );

    \I__1698\ : IoSpan4Mux
    port map (
            O => \N__8108\,
            I => \N__8105\
        );

    \I__1697\ : Span4Mux_s3_v
    port map (
            O => \N__8105\,
            I => \N__8102\
        );

    \I__1696\ : Span4Mux_h
    port map (
            O => \N__8102\,
            I => \N__8099\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__8099\,
            I => \un1_D_UU_040_2\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8096\,
            I => \N__8093\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8093\,
            I => \N__8090\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__8090\,
            I => \N__8087\
        );

    \I__1691\ : Span4Mux_v
    port map (
            O => \N__8087\,
            I => \N__8084\
        );

    \I__1690\ : Sp12to4
    port map (
            O => \N__8084\,
            I => \N__8081\
        );

    \I__1689\ : Span12Mux_h
    port map (
            O => \N__8081\,
            I => \N__8078\
        );

    \I__1688\ : Odrv12
    port map (
            O => \N__8078\,
            I => \D_UU_040_in_5\
        );

    \I__1687\ : IoInMux
    port map (
            O => \N__8075\,
            I => \N__8072\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8072\,
            I => \N__8069\
        );

    \I__1685\ : IoSpan4Mux
    port map (
            O => \N__8069\,
            I => \N__8065\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8068\,
            I => \N__8062\
        );

    \I__1683\ : IoSpan4Mux
    port map (
            O => \N__8065\,
            I => \N__8059\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__8062\,
            I => \N__8056\
        );

    \I__1681\ : Span4Mux_s2_h
    port map (
            O => \N__8059\,
            I => \N__8053\
        );

    \I__1680\ : Span4Mux_v
    port map (
            O => \N__8056\,
            I => \N__8050\
        );

    \I__1679\ : Sp12to4
    port map (
            O => \N__8053\,
            I => \N__8047\
        );

    \I__1678\ : Sp12to4
    port map (
            O => \N__8050\,
            I => \N__8044\
        );

    \I__1677\ : Span12Mux_h
    port map (
            O => \N__8047\,
            I => \N__8041\
        );

    \I__1676\ : Span12Mux_h
    port map (
            O => \N__8044\,
            I => \N__8038\
        );

    \I__1675\ : Span12Mux_h
    port map (
            O => \N__8041\,
            I => \N__8035\
        );

    \I__1674\ : Span12Mux_v
    port map (
            O => \N__8038\,
            I => \N__8032\
        );

    \I__1673\ : Odrv12
    port map (
            O => \N__8035\,
            I => \D_LM_040_in_5\
        );

    \I__1672\ : Odrv12
    port map (
            O => \N__8032\,
            I => \D_LM_040_in_5\
        );

    \I__1671\ : IoInMux
    port map (
            O => \N__8027\,
            I => \N__8024\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8024\,
            I => \N__8021\
        );

    \I__1669\ : Span4Mux_s3_h
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__1668\ : Sp12to4
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__1667\ : Span12Mux_s7_v
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__1666\ : Span12Mux_h
    port map (
            O => \N__8012\,
            I => \N__8009\
        );

    \I__1665\ : Odrv12
    port map (
            O => \N__8009\,
            I => \un1_D_UU_040_5\
        );

    \I__1664\ : InMux
    port map (
            O => \N__8006\,
            I => \N__8002\
        );

    \I__1663\ : InMux
    port map (
            O => \N__8005\,
            I => \N__7999\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__8002\,
            I => \N__7996\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__7999\,
            I => \N__7993\
        );

    \I__1660\ : Span4Mux_v
    port map (
            O => \N__7996\,
            I => \N__7989\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__7993\,
            I => \N__7986\
        );

    \I__1658\ : InMux
    port map (
            O => \N__7992\,
            I => \N__7983\
        );

    \I__1657\ : Span4Mux_v
    port map (
            O => \N__7989\,
            I => \N__7980\
        );

    \I__1656\ : Span4Mux_v
    port map (
            O => \N__7986\,
            I => \N__7975\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__7983\,
            I => \N__7975\
        );

    \I__1654\ : Span4Mux_v
    port map (
            O => \N__7980\,
            I => \N__7970\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__7975\,
            I => \N__7970\
        );

    \I__1652\ : Sp12to4
    port map (
            O => \N__7970\,
            I => \N__7967\
        );

    \I__1651\ : Span12Mux_h
    port map (
            O => \N__7967\,
            I => \N__7964\
        );

    \I__1650\ : Odrv12
    port map (
            O => \N__7964\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__1649\ : InMux
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__7958\,
            I => \N__7955\
        );

    \I__1647\ : Span12Mux_s7_v
    port map (
            O => \N__7955\,
            I => \N__7952\
        );

    \I__1646\ : Odrv12
    port map (
            O => \N__7952\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__1645\ : IoInMux
    port map (
            O => \N__7949\,
            I => \N__7946\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7946\,
            I => \N__7943\
        );

    \I__1643\ : Span4Mux_s2_v
    port map (
            O => \N__7943\,
            I => \N__7940\
        );

    \I__1642\ : Span4Mux_h
    port map (
            O => \N__7940\,
            I => \N__7937\
        );

    \I__1641\ : Span4Mux_v
    port map (
            O => \N__7937\,
            I => \N__7934\
        );

    \I__1640\ : Sp12to4
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__1639\ : Odrv12
    port map (
            O => \N__7931\,
            I => \un1_D_UU_AMIGA_3\
        );

    \I__1638\ : InMux
    port map (
            O => \N__7928\,
            I => \N__7924\
        );

    \I__1637\ : InMux
    port map (
            O => \N__7927\,
            I => \N__7921\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__7924\,
            I => \N__7917\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__7921\,
            I => \N__7914\
        );

    \I__1634\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7911\
        );

    \I__1633\ : Span12Mux_v
    port map (
            O => \N__7917\,
            I => \N__7904\
        );

    \I__1632\ : Span12Mux_s9_v
    port map (
            O => \N__7914\,
            I => \N__7904\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__7911\,
            I => \N__7904\
        );

    \I__1630\ : Span12Mux_h
    port map (
            O => \N__7904\,
            I => \N__7901\
        );

    \I__1629\ : Odrv12
    port map (
            O => \N__7901\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7895\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__7895\,
            I => \N__7892\
        );

    \I__1626\ : Span12Mux_s11_v
    port map (
            O => \N__7892\,
            I => \N__7889\
        );

    \I__1625\ : Odrv12
    port map (
            O => \N__7889\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__1624\ : IoInMux
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7883\,
            I => \N__7880\
        );

    \I__1622\ : Span4Mux_s0_v
    port map (
            O => \N__7880\,
            I => \N__7877\
        );

    \I__1621\ : Sp12to4
    port map (
            O => \N__7877\,
            I => \N__7874\
        );

    \I__1620\ : Span12Mux_h
    port map (
            O => \N__7874\,
            I => \N__7871\
        );

    \I__1619\ : Odrv12
    port map (
            O => \N__7871\,
            I => \un1_D_UU_AMIGA_6\
        );

    \I__1618\ : CEMux
    port map (
            O => \N__7868\,
            I => \N__7862\
        );

    \I__1617\ : CEMux
    port map (
            O => \N__7867\,
            I => \N__7859\
        );

    \I__1616\ : CEMux
    port map (
            O => \N__7866\,
            I => \N__7854\
        );

    \I__1615\ : CEMux
    port map (
            O => \N__7865\,
            I => \N__7851\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__7862\,
            I => \N__7848\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__7859\,
            I => \N__7845\
        );

    \I__1612\ : CEMux
    port map (
            O => \N__7858\,
            I => \N__7842\
        );

    \I__1611\ : CEMux
    port map (
            O => \N__7857\,
            I => \N__7839\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__7854\,
            I => \N__7836\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__7851\,
            I => \N__7833\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__7848\,
            I => \N__7826\
        );

    \I__1607\ : Span4Mux_h
    port map (
            O => \N__7845\,
            I => \N__7826\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__7842\,
            I => \N__7826\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__7839\,
            I => \N__7823\
        );

    \I__1604\ : Span4Mux_v
    port map (
            O => \N__7836\,
            I => \N__7820\
        );

    \I__1603\ : Span4Mux_h
    port map (
            O => \N__7833\,
            I => \N__7817\
        );

    \I__1602\ : Span4Mux_v
    port map (
            O => \N__7826\,
            I => \N__7814\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__7823\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0\
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__7820\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0\
        );

    \I__1599\ : Odrv4
    port map (
            O => \N__7817\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0\
        );

    \I__1598\ : Odrv4
    port map (
            O => \N__7814\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0\
        );

    \I__1597\ : SRMux
    port map (
            O => \N__7805\,
            I => \N__7802\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__7802\,
            I => \N__7799\
        );

    \I__1595\ : Span4Mux_h
    port map (
            O => \N__7799\,
            I => \N__7791\
        );

    \I__1594\ : SRMux
    port map (
            O => \N__7798\,
            I => \N__7788\
        );

    \I__1593\ : SRMux
    port map (
            O => \N__7797\,
            I => \N__7785\
        );

    \I__1592\ : SRMux
    port map (
            O => \N__7796\,
            I => \N__7782\
        );

    \I__1591\ : SRMux
    port map (
            O => \N__7795\,
            I => \N__7779\
        );

    \I__1590\ : SRMux
    port map (
            O => \N__7794\,
            I => \N__7776\
        );

    \I__1589\ : Odrv4
    port map (
            O => \N__7791\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__7788\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__7785\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__7782\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7779\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7776\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7763\,
            I => \N__7760\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7760\,
            I => \N__7757\
        );

    \I__1581\ : Glb2LocalMux
    port map (
            O => \N__7757\,
            I => \N__7754\
        );

    \I__1580\ : GlobalMux
    port map (
            O => \N__7754\,
            I => \CLK80\
        );

    \I__1579\ : IoInMux
    port map (
            O => \N__7751\,
            I => \N__7747\
        );

    \I__1578\ : IoInMux
    port map (
            O => \N__7750\,
            I => \N__7744\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7747\,
            I => \N__7741\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__7744\,
            I => \N__7738\
        );

    \I__1575\ : Span4Mux_s3_v
    port map (
            O => \N__7741\,
            I => \N__7735\
        );

    \I__1574\ : IoSpan4Mux
    port map (
            O => \N__7738\,
            I => \N__7732\
        );

    \I__1573\ : Span4Mux_v
    port map (
            O => \N__7735\,
            I => \N__7729\
        );

    \I__1572\ : Span4Mux_s3_h
    port map (
            O => \N__7732\,
            I => \N__7726\
        );

    \I__1571\ : Span4Mux_v
    port map (
            O => \N__7729\,
            I => \N__7723\
        );

    \I__1570\ : Span4Mux_h
    port map (
            O => \N__7726\,
            I => \N__7720\
        );

    \I__1569\ : Span4Mux_v
    port map (
            O => \N__7723\,
            I => \N__7717\
        );

    \I__1568\ : Sp12to4
    port map (
            O => \N__7720\,
            I => \N__7714\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__7717\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1566\ : Odrv12
    port map (
            O => \N__7714\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7709\,
            I => \N__7706\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__7706\,
            I => \N__7703\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__7703\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7700\,
            I => \N__7695\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7699\,
            I => \N__7692\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7698\,
            I => \N__7689\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7695\,
            I => \N__7684\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7692\,
            I => \N__7684\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7689\,
            I => \N__7681\
        );

    \I__1556\ : Span4Mux_v
    port map (
            O => \N__7684\,
            I => \N__7678\
        );

    \I__1555\ : Span4Mux_v
    port map (
            O => \N__7681\,
            I => \N__7675\
        );

    \I__1554\ : Sp12to4
    port map (
            O => \N__7678\,
            I => \N__7672\
        );

    \I__1553\ : Span4Mux_h
    port map (
            O => \N__7675\,
            I => \N__7669\
        );

    \I__1552\ : Span12Mux_h
    port map (
            O => \N__7672\,
            I => \N__7664\
        );

    \I__1551\ : Sp12to4
    port map (
            O => \N__7669\,
            I => \N__7664\
        );

    \I__1550\ : Odrv12
    port map (
            O => \N__7664\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__1549\ : IoInMux
    port map (
            O => \N__7661\,
            I => \N__7658\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7658\,
            I => \N__7655\
        );

    \I__1547\ : IoSpan4Mux
    port map (
            O => \N__7655\,
            I => \N__7652\
        );

    \I__1546\ : Span4Mux_s0_v
    port map (
            O => \N__7652\,
            I => \N__7649\
        );

    \I__1545\ : Sp12to4
    port map (
            O => \N__7649\,
            I => \N__7646\
        );

    \I__1544\ : Span12Mux_v
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__1543\ : Odrv12
    port map (
            O => \N__7643\,
            I => \un1_D_UU_AMIGA_2\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7637\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__7637\,
            I => \N__7634\
        );

    \I__1540\ : Odrv12
    port map (
            O => \N__7634\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__1539\ : IoInMux
    port map (
            O => \N__7631\,
            I => \N__7628\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7628\,
            I => \N__7625\
        );

    \I__1537\ : Span4Mux_s0_v
    port map (
            O => \N__7625\,
            I => \N__7622\
        );

    \I__1536\ : Sp12to4
    port map (
            O => \N__7622\,
            I => \N__7619\
        );

    \I__1535\ : Span12Mux_s9_h
    port map (
            O => \N__7619\,
            I => \N__7616\
        );

    \I__1534\ : Span12Mux_v
    port map (
            O => \N__7616\,
            I => \N__7613\
        );

    \I__1533\ : Odrv12
    port map (
            O => \N__7613\,
            I => \un1_D_UU_AMIGA_7\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7610\,
            I => \N__7607\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__7607\,
            I => \N__7604\
        );

    \I__1530\ : Odrv4
    port map (
            O => \N__7604\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7601\,
            I => \N__7596\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7600\,
            I => \N__7593\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7599\,
            I => \N__7590\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__7596\,
            I => \N__7585\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7593\,
            I => \N__7585\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7590\,
            I => \N__7582\
        );

    \I__1523\ : Span4Mux_v
    port map (
            O => \N__7585\,
            I => \N__7579\
        );

    \I__1522\ : Span12Mux_h
    port map (
            O => \N__7582\,
            I => \N__7576\
        );

    \I__1521\ : Sp12to4
    port map (
            O => \N__7579\,
            I => \N__7573\
        );

    \I__1520\ : Span12Mux_v
    port map (
            O => \N__7576\,
            I => \N__7570\
        );

    \I__1519\ : Span12Mux_h
    port map (
            O => \N__7573\,
            I => \N__7567\
        );

    \I__1518\ : Odrv12
    port map (
            O => \N__7570\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__1517\ : Odrv12
    port map (
            O => \N__7567\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__1516\ : IoInMux
    port map (
            O => \N__7562\,
            I => \N__7559\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__7559\,
            I => \N__7556\
        );

    \I__1514\ : IoSpan4Mux
    port map (
            O => \N__7556\,
            I => \N__7553\
        );

    \I__1513\ : Span4Mux_s2_v
    port map (
            O => \N__7553\,
            I => \N__7550\
        );

    \I__1512\ : Sp12to4
    port map (
            O => \N__7550\,
            I => \N__7547\
        );

    \I__1511\ : Span12Mux_h
    port map (
            O => \N__7547\,
            I => \N__7544\
        );

    \I__1510\ : Odrv12
    port map (
            O => \N__7544\,
            I => \un1_D_UU_AMIGA_4\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7541\,
            I => \N__7537\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7540\,
            I => \N__7533\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7537\,
            I => \N__7530\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7536\,
            I => \N__7527\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7533\,
            I => \N__7524\
        );

    \I__1504\ : Span4Mux_v
    port map (
            O => \N__7530\,
            I => \N__7519\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7527\,
            I => \N__7519\
        );

    \I__1502\ : Sp12to4
    port map (
            O => \N__7524\,
            I => \N__7516\
        );

    \I__1501\ : Span4Mux_v
    port map (
            O => \N__7519\,
            I => \N__7513\
        );

    \I__1500\ : Span12Mux_v
    port map (
            O => \N__7516\,
            I => \N__7510\
        );

    \I__1499\ : Span4Mux_v
    port map (
            O => \N__7513\,
            I => \N__7507\
        );

    \I__1498\ : Span12Mux_v
    port map (
            O => \N__7510\,
            I => \N__7504\
        );

    \I__1497\ : Sp12to4
    port map (
            O => \N__7507\,
            I => \N__7501\
        );

    \I__1496\ : Span12Mux_h
    port map (
            O => \N__7504\,
            I => \N__7498\
        );

    \I__1495\ : Span12Mux_h
    port map (
            O => \N__7501\,
            I => \N__7495\
        );

    \I__1494\ : Odrv12
    port map (
            O => \N__7498\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1493\ : Odrv12
    port map (
            O => \N__7495\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7490\,
            I => \N__7487\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7487\,
            I => \N__7484\
        );

    \I__1490\ : Span4Mux_v
    port map (
            O => \N__7484\,
            I => \N__7481\
        );

    \I__1489\ : Odrv4
    port map (
            O => \N__7481\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\
        );

    \I__1488\ : IoInMux
    port map (
            O => \N__7478\,
            I => \N__7475\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7475\,
            I => \N__7472\
        );

    \I__1486\ : IoSpan4Mux
    port map (
            O => \N__7472\,
            I => \N__7469\
        );

    \I__1485\ : Span4Mux_s2_h
    port map (
            O => \N__7469\,
            I => \N__7466\
        );

    \I__1484\ : Sp12to4
    port map (
            O => \N__7466\,
            I => \N__7463\
        );

    \I__1483\ : Span12Mux_h
    port map (
            O => \N__7463\,
            I => \N__7460\
        );

    \I__1482\ : Odrv12
    port map (
            O => \N__7460\,
            I => \un1_D_UM_AMIGA_3\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7457\,
            I => \N__7454\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__7454\,
            I => \N__7451\
        );

    \I__1479\ : Span4Mux_v
    port map (
            O => \N__7451\,
            I => \N__7448\
        );

    \I__1478\ : Sp12to4
    port map (
            O => \N__7448\,
            I => \N__7445\
        );

    \I__1477\ : Span12Mux_h
    port map (
            O => \N__7445\,
            I => \N__7442\
        );

    \I__1476\ : Odrv12
    port map (
            O => \N__7442\,
            I => \D_LL_AMIGA_in_5\
        );

    \I__1475\ : IoInMux
    port map (
            O => \N__7439\,
            I => \N__7436\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7436\,
            I => \N__7433\
        );

    \I__1473\ : IoSpan4Mux
    port map (
            O => \N__7433\,
            I => \N__7430\
        );

    \I__1472\ : Span4Mux_s2_h
    port map (
            O => \N__7430\,
            I => \N__7427\
        );

    \I__1471\ : Sp12to4
    port map (
            O => \N__7427\,
            I => \N__7424\
        );

    \I__1470\ : Span12Mux_h
    port map (
            O => \N__7424\,
            I => \N__7421\
        );

    \I__1469\ : Odrv12
    port map (
            O => \N__7421\,
            I => \un2_D_LL_AMIGA_5\
        );

    \I__1468\ : IoInMux
    port map (
            O => \N__7418\,
            I => \N__7415\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__7415\,
            I => \N__7411\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__7414\,
            I => \N__7406\
        );

    \I__1465\ : Span4Mux_s1_v
    port map (
            O => \N__7411\,
            I => \N__7402\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7410\,
            I => \N__7399\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7409\,
            I => \N__7396\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7406\,
            I => \N__7391\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7405\,
            I => \N__7391\
        );

    \I__1460\ : Span4Mux_v
    port map (
            O => \N__7402\,
            I => \N__7388\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7399\,
            I => \N__7383\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7396\,
            I => \N__7378\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7391\,
            I => \N__7378\
        );

    \I__1456\ : Sp12to4
    port map (
            O => \N__7388\,
            I => \N__7375\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7387\,
            I => \N__7372\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7369\
        );

    \I__1453\ : Span4Mux_v
    port map (
            O => \N__7383\,
            I => \N__7363\
        );

    \I__1452\ : Span4Mux_v
    port map (
            O => \N__7378\,
            I => \N__7363\
        );

    \I__1451\ : Span12Mux_h
    port map (
            O => \N__7375\,
            I => \N__7356\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7372\,
            I => \N__7356\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7369\,
            I => \N__7356\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7368\,
            I => \N__7353\
        );

    \I__1447\ : Sp12to4
    port map (
            O => \N__7363\,
            I => \N__7346\
        );

    \I__1446\ : Span12Mux_v
    port map (
            O => \N__7356\,
            I => \N__7346\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7353\,
            I => \N__7346\
        );

    \I__1444\ : Span12Mux_v
    port map (
            O => \N__7346\,
            I => \N__7343\
        );

    \I__1443\ : Odrv12
    port map (
            O => \N__7343\,
            I => \TACKn_in\
        );

    \I__1442\ : IoInMux
    port map (
            O => \N__7340\,
            I => \N__7337\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7337\,
            I => \N__7334\
        );

    \I__1440\ : Span4Mux_s1_v
    port map (
            O => \N__7334\,
            I => \N__7326\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7323\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7320\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7331\,
            I => \N__7317\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7330\,
            I => \N__7312\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7329\,
            I => \N__7312\
        );

    \I__1434\ : Span4Mux_v
    port map (
            O => \N__7326\,
            I => \N__7308\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7323\,
            I => \N__7299\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7320\,
            I => \N__7299\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__7317\,
            I => \N__7299\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__7312\,
            I => \N__7299\
        );

    \I__1429\ : InMux
    port map (
            O => \N__7311\,
            I => \N__7296\
        );

    \I__1428\ : Span4Mux_v
    port map (
            O => \N__7308\,
            I => \N__7293\
        );

    \I__1427\ : Span4Mux_v
    port map (
            O => \N__7299\,
            I => \N__7288\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__7296\,
            I => \N__7288\
        );

    \I__1425\ : Sp12to4
    port map (
            O => \N__7293\,
            I => \N__7285\
        );

    \I__1424\ : Span4Mux_v
    port map (
            O => \N__7288\,
            I => \N__7282\
        );

    \I__1423\ : Span12Mux_h
    port map (
            O => \N__7285\,
            I => \N__7279\
        );

    \I__1422\ : Span4Mux_h
    port map (
            O => \N__7282\,
            I => \N__7276\
        );

    \I__1421\ : Span12Mux_v
    port map (
            O => \N__7279\,
            I => \N__7271\
        );

    \I__1420\ : Sp12to4
    port map (
            O => \N__7276\,
            I => \N__7271\
        );

    \I__1419\ : Odrv12
    port map (
            O => \N__7271\,
            I => \TEAn_c\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7268\,
            I => \N__7264\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7267\,
            I => \N__7261\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7264\,
            I => \N__7256\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__7261\,
            I => \N__7256\
        );

    \I__1414\ : Span4Mux_v
    port map (
            O => \N__7256\,
            I => \N__7250\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7255\,
            I => \N__7247\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__7254\,
            I => \N__7243\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7253\,
            I => \N__7237\
        );

    \I__1410\ : Span4Mux_v
    port map (
            O => \N__7250\,
            I => \N__7232\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__7247\,
            I => \N__7232\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7246\,
            I => \N__7227\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7243\,
            I => \N__7227\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7242\,
            I => \N__7224\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7241\,
            I => \N__7221\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7240\,
            I => \N__7218\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7237\,
            I => \N__7207\
        );

    \I__1402\ : Sp12to4
    port map (
            O => \N__7232\,
            I => \N__7207\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7227\,
            I => \N__7207\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7224\,
            I => \N__7207\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7221\,
            I => \N__7207\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__7218\,
            I => \N__7204\
        );

    \I__1397\ : Span12Mux_h
    port map (
            O => \N__7207\,
            I => \N__7201\
        );

    \I__1396\ : Span12Mux_v
    port map (
            O => \N__7204\,
            I => \N__7198\
        );

    \I__1395\ : Span12Mux_v
    port map (
            O => \N__7201\,
            I => \N__7195\
        );

    \I__1394\ : Odrv12
    port map (
            O => \N__7198\,
            I => \RESETn_c\
        );

    \I__1393\ : Odrv12
    port map (
            O => \N__7195\,
            I => \RESETn_c\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7190\,
            I => \N__7187\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7187\,
            I => \N__7183\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__7186\,
            I => \N__7180\
        );

    \I__1389\ : Span4Mux_v
    port map (
            O => \N__7183\,
            I => \N__7177\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7180\,
            I => \N__7174\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__7177\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7174\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__7169\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7166\,
            I => \N__7162\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7165\,
            I => \N__7158\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__7162\,
            I => \N__7155\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7161\,
            I => \N__7151\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7158\,
            I => \N__7145\
        );

    \I__1379\ : Span4Mux_v
    port map (
            O => \N__7155\,
            I => \N__7145\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7154\,
            I => \N__7142\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7151\,
            I => \N__7139\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7150\,
            I => \N__7136\
        );

    \I__1375\ : Odrv4
    port map (
            O => \N__7145\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7142\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__7139\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7136\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1371\ : InMux
    port map (
            O => \N__7127\,
            I => \N__7124\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__7124\,
            I => \N__7120\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__7123\,
            I => \N__7117\
        );

    \I__1368\ : Span4Mux_v
    port map (
            O => \N__7120\,
            I => \N__7114\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7117\,
            I => \N__7111\
        );

    \I__1366\ : Odrv4
    port map (
            O => \N__7114\,
            I => \U111_CYCLE_SM.TA_DISZ0\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__7111\,
            I => \U111_CYCLE_SM.TA_DISZ0\
        );

    \I__1364\ : IoInMux
    port map (
            O => \N__7106\,
            I => \N__7103\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__7103\,
            I => \N__7100\
        );

    \I__1362\ : Span4Mux_s3_v
    port map (
            O => \N__7100\,
            I => \N__7097\
        );

    \I__1361\ : Span4Mux_h
    port map (
            O => \N__7097\,
            I => \N__7094\
        );

    \I__1360\ : Span4Mux_v
    port map (
            O => \N__7094\,
            I => \N__7091\
        );

    \I__1359\ : Span4Mux_v
    port map (
            O => \N__7091\,
            I => \N__7088\
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__7088\,
            I => \TAn_1_i\
        );

    \I__1357\ : InMux
    port map (
            O => \N__7085\,
            I => \N__7082\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7082\,
            I => \N__7079\
        );

    \I__1355\ : Span4Mux_v
    port map (
            O => \N__7079\,
            I => \N__7076\
        );

    \I__1354\ : Sp12to4
    port map (
            O => \N__7076\,
            I => \N__7073\
        );

    \I__1353\ : Span12Mux_h
    port map (
            O => \N__7073\,
            I => \N__7070\
        );

    \I__1352\ : Odrv12
    port map (
            O => \N__7070\,
            I => \D_LM_AMIGA_in_4\
        );

    \I__1351\ : IoInMux
    port map (
            O => \N__7067\,
            I => \N__7064\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__7064\,
            I => \N__7061\
        );

    \I__1349\ : IoSpan4Mux
    port map (
            O => \N__7061\,
            I => \N__7058\
        );

    \I__1348\ : Span4Mux_s2_h
    port map (
            O => \N__7058\,
            I => \N__7055\
        );

    \I__1347\ : Span4Mux_h
    port map (
            O => \N__7055\,
            I => \N__7052\
        );

    \I__1346\ : Sp12to4
    port map (
            O => \N__7052\,
            I => \N__7049\
        );

    \I__1345\ : Span12Mux_h
    port map (
            O => \N__7049\,
            I => \N__7046\
        );

    \I__1344\ : Odrv12
    port map (
            O => \N__7046\,
            I => \un2_D_LM_AMIGA_4\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7043\,
            I => \N__7040\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7040\,
            I => \N__7037\
        );

    \I__1341\ : Span4Mux_v
    port map (
            O => \N__7037\,
            I => \N__7034\
        );

    \I__1340\ : Odrv4
    port map (
            O => \N__7034\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7026\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7030\,
            I => \N__7023\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7029\,
            I => \N__7020\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7026\,
            I => \N__7017\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7023\,
            I => \N__7014\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7020\,
            I => \N__7011\
        );

    \I__1333\ : Span4Mux_v
    port map (
            O => \N__7017\,
            I => \N__7006\
        );

    \I__1332\ : Span4Mux_v
    port map (
            O => \N__7014\,
            I => \N__7006\
        );

    \I__1331\ : Span4Mux_v
    port map (
            O => \N__7011\,
            I => \N__7003\
        );

    \I__1330\ : Sp12to4
    port map (
            O => \N__7006\,
            I => \N__6998\
        );

    \I__1329\ : Sp12to4
    port map (
            O => \N__7003\,
            I => \N__6998\
        );

    \I__1328\ : Span12Mux_h
    port map (
            O => \N__6998\,
            I => \N__6995\
        );

    \I__1327\ : Span12Mux_v
    port map (
            O => \N__6995\,
            I => \N__6992\
        );

    \I__1326\ : Odrv12
    port map (
            O => \N__6992\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1325\ : IoInMux
    port map (
            O => \N__6989\,
            I => \N__6986\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6986\,
            I => \N__6983\
        );

    \I__1323\ : IoSpan4Mux
    port map (
            O => \N__6983\,
            I => \N__6980\
        );

    \I__1322\ : Sp12to4
    port map (
            O => \N__6980\,
            I => \N__6977\
        );

    \I__1321\ : Span12Mux_v
    port map (
            O => \N__6977\,
            I => \N__6974\
        );

    \I__1320\ : Span12Mux_h
    port map (
            O => \N__6974\,
            I => \N__6971\
        );

    \I__1319\ : Odrv12
    port map (
            O => \N__6971\,
            I => \un1_D_UU_AMIGA_5\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6968\,
            I => \N__6965\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6965\,
            I => \N__6960\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6964\,
            I => \N__6957\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6963\,
            I => \N__6954\
        );

    \I__1314\ : Span4Mux_v
    port map (
            O => \N__6960\,
            I => \N__6949\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6957\,
            I => \N__6949\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6954\,
            I => \N__6946\
        );

    \I__1311\ : Span4Mux_v
    port map (
            O => \N__6949\,
            I => \N__6943\
        );

    \I__1310\ : Sp12to4
    port map (
            O => \N__6946\,
            I => \N__6940\
        );

    \I__1309\ : Sp12to4
    port map (
            O => \N__6943\,
            I => \N__6937\
        );

    \I__1308\ : Span12Mux_v
    port map (
            O => \N__6940\,
            I => \N__6934\
        );

    \I__1307\ : Span12Mux_h
    port map (
            O => \N__6937\,
            I => \N__6931\
        );

    \I__1306\ : Odrv12
    port map (
            O => \N__6934\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__1305\ : Odrv12
    port map (
            O => \N__6931\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6926\,
            I => \N__6923\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6923\,
            I => \N__6920\
        );

    \I__1302\ : Odrv12
    port map (
            O => \N__6920\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\
        );

    \I__1301\ : IoInMux
    port map (
            O => \N__6917\,
            I => \N__6914\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6914\,
            I => \N__6911\
        );

    \I__1299\ : Span4Mux_s3_h
    port map (
            O => \N__6911\,
            I => \N__6908\
        );

    \I__1298\ : Span4Mux_h
    port map (
            O => \N__6908\,
            I => \N__6905\
        );

    \I__1297\ : Sp12to4
    port map (
            O => \N__6905\,
            I => \N__6902\
        );

    \I__1296\ : Span12Mux_s11_v
    port map (
            O => \N__6902\,
            I => \N__6899\
        );

    \I__1295\ : Odrv12
    port map (
            O => \N__6899\,
            I => \un1_D_UM_AMIGA_1\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6896\,
            I => \N__6893\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6893\,
            I => \N__6890\
        );

    \I__1292\ : Odrv12
    port map (
            O => \N__6890\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6887\,
            I => \N__6883\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6886\,
            I => \N__6880\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6883\,
            I => \N__6877\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6880\,
            I => \N__6874\
        );

    \I__1287\ : Span4Mux_v
    port map (
            O => \N__6877\,
            I => \N__6871\
        );

    \I__1286\ : Span4Mux_v
    port map (
            O => \N__6874\,
            I => \N__6868\
        );

    \I__1285\ : Sp12to4
    port map (
            O => \N__6871\,
            I => \N__6864\
        );

    \I__1284\ : Span4Mux_v
    port map (
            O => \N__6868\,
            I => \N__6861\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6867\,
            I => \N__6858\
        );

    \I__1282\ : Span12Mux_h
    port map (
            O => \N__6864\,
            I => \N__6855\
        );

    \I__1281\ : Sp12to4
    port map (
            O => \N__6861\,
            I => \N__6850\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__6858\,
            I => \N__6850\
        );

    \I__1279\ : Span12Mux_v
    port map (
            O => \N__6855\,
            I => \N__6847\
        );

    \I__1278\ : Span12Mux_h
    port map (
            O => \N__6850\,
            I => \N__6844\
        );

    \I__1277\ : Odrv12
    port map (
            O => \N__6847\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1276\ : Odrv12
    port map (
            O => \N__6844\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1275\ : IoInMux
    port map (
            O => \N__6839\,
            I => \N__6836\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__6836\,
            I => \N__6833\
        );

    \I__1273\ : Span4Mux_s3_v
    port map (
            O => \N__6833\,
            I => \N__6830\
        );

    \I__1272\ : Span4Mux_v
    port map (
            O => \N__6830\,
            I => \N__6827\
        );

    \I__1271\ : Sp12to4
    port map (
            O => \N__6827\,
            I => \N__6824\
        );

    \I__1270\ : Span12Mux_h
    port map (
            O => \N__6824\,
            I => \N__6821\
        );

    \I__1269\ : Odrv12
    port map (
            O => \N__6821\,
            I => \un1_D_UU_AMIGA_0\
        );

    \I__1268\ : IoInMux
    port map (
            O => \N__6818\,
            I => \N__6815\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__6815\,
            I => \N__6812\
        );

    \I__1266\ : Odrv12
    port map (
            O => \N__6812\,
            I => \LBENn_c_i_0\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6809\,
            I => \N__6806\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6806\,
            I => \N__6803\
        );

    \I__1263\ : Span4Mux_v
    port map (
            O => \N__6803\,
            I => \N__6800\
        );

    \I__1262\ : Sp12to4
    port map (
            O => \N__6800\,
            I => \N__6797\
        );

    \I__1261\ : Span12Mux_h
    port map (
            O => \N__6797\,
            I => \N__6794\
        );

    \I__1260\ : Odrv12
    port map (
            O => \N__6794\,
            I => \D_LL_AMIGA_in_7\
        );

    \I__1259\ : IoInMux
    port map (
            O => \N__6791\,
            I => \N__6788\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__6788\,
            I => \N__6785\
        );

    \I__1257\ : IoSpan4Mux
    port map (
            O => \N__6785\,
            I => \N__6782\
        );

    \I__1256\ : Span4Mux_s3_h
    port map (
            O => \N__6782\,
            I => \N__6779\
        );

    \I__1255\ : Sp12to4
    port map (
            O => \N__6779\,
            I => \N__6776\
        );

    \I__1254\ : Span12Mux_h
    port map (
            O => \N__6776\,
            I => \N__6773\
        );

    \I__1253\ : Odrv12
    port map (
            O => \N__6773\,
            I => \un2_D_LL_AMIGA_7\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6770\,
            I => \N__6767\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__6767\,
            I => \N__6761\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6766\,
            I => \N__6757\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6754\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6764\,
            I => \N__6751\
        );

    \I__1247\ : Span12Mux_s6_h
    port map (
            O => \N__6761\,
            I => \N__6748\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6760\,
            I => \N__6745\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6757\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6754\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__6751\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1242\ : Odrv12
    port map (
            O => \N__6748\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6745\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1240\ : CascadeMux
    port map (
            O => \N__6734\,
            I => \N__6731\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6728\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6728\,
            I => \N__6725\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__6725\,
            I => \U111_CYCLE_SM.N_119_0\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6722\,
            I => \N__6719\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6719\,
            I => \N__6716\
        );

    \I__1234\ : Odrv4
    port map (
            O => \N__6716\,
            I => \U111_CYCLE_SM.N_117_0\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6713\,
            I => \N__6702\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6712\,
            I => \N__6702\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6711\,
            I => \N__6702\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6710\,
            I => \N__6697\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6709\,
            I => \N__6697\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__6702\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6697\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__6692\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_cascade_\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6689\,
            I => \N__6686\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6686\,
            I => \N__6682\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6685\,
            I => \N__6679\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__6682\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__6679\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__6674\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1_cascade_\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6671\,
            I => \N__6668\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6668\,
            I => \N__6665\
        );

    \I__1217\ : Span4Mux_h
    port map (
            O => \N__6665\,
            I => \N__6659\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6664\,
            I => \N__6656\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6663\,
            I => \N__6653\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6662\,
            I => \N__6650\
        );

    \I__1213\ : Odrv4
    port map (
            O => \N__6659\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6656\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6653\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6650\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6641\,
            I => \N__6634\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6627\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6639\,
            I => \N__6627\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6638\,
            I => \N__6627\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6637\,
            I => \N__6624\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__6634\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6627\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__6624\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6617\,
            I => \N__6612\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6616\,
            I => \N__6609\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6615\,
            I => \N__6606\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6612\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6609\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__6606\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6599\,
            I => \N__6592\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6598\,
            I => \N__6589\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6597\,
            I => \N__6584\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6584\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6581\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__6592\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__6589\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6584\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__6581\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__6572\,
            I => \U111_CYCLE_SM.N_131_cascade_\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6569\,
            I => \N__6566\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6566\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0\
        );

    \I__1183\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6560\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6560\,
            I => \U111_CYCLE_SM.TS_EN6\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6557\,
            I => \N__6554\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6554\,
            I => \N__6550\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6553\,
            I => \N__6547\
        );

    \I__1178\ : Odrv4
    port map (
            O => \N__6550\,
            I => \U111_CYCLE_SM.N_144\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6547\,
            I => \U111_CYCLE_SM.N_144\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6542\,
            I => \N__6539\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6539\,
            I => \N__6536\
        );

    \I__1174\ : Span12Mux_s9_v
    port map (
            O => \N__6536\,
            I => \N__6533\
        );

    \I__1173\ : Odrv12
    port map (
            O => \N__6533\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6530\,
            I => \N__6527\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6527\,
            I => \N__6524\
        );

    \I__1170\ : Span4Mux_v
    port map (
            O => \N__6524\,
            I => \N__6519\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6523\,
            I => \N__6516\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6522\,
            I => \N__6513\
        );

    \I__1167\ : Span4Mux_v
    port map (
            O => \N__6519\,
            I => \N__6510\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6516\,
            I => \N__6507\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6513\,
            I => \N__6504\
        );

    \I__1164\ : Span4Mux_v
    port map (
            O => \N__6510\,
            I => \N__6501\
        );

    \I__1163\ : Span4Mux_v
    port map (
            O => \N__6507\,
            I => \N__6498\
        );

    \I__1162\ : Span12Mux_h
    port map (
            O => \N__6504\,
            I => \N__6495\
        );

    \I__1161\ : Sp12to4
    port map (
            O => \N__6501\,
            I => \N__6490\
        );

    \I__1160\ : Sp12to4
    port map (
            O => \N__6498\,
            I => \N__6490\
        );

    \I__1159\ : Span12Mux_v
    port map (
            O => \N__6495\,
            I => \N__6485\
        );

    \I__1158\ : Span12Mux_h
    port map (
            O => \N__6490\,
            I => \N__6485\
        );

    \I__1157\ : Odrv12
    port map (
            O => \N__6485\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__1156\ : IoInMux
    port map (
            O => \N__6482\,
            I => \N__6479\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6479\,
            I => \N__6476\
        );

    \I__1154\ : Span4Mux_s3_h
    port map (
            O => \N__6476\,
            I => \N__6473\
        );

    \I__1153\ : Span4Mux_h
    port map (
            O => \N__6473\,
            I => \N__6470\
        );

    \I__1152\ : Sp12to4
    port map (
            O => \N__6470\,
            I => \N__6467\
        );

    \I__1151\ : Span12Mux_s8_v
    port map (
            O => \N__6467\,
            I => \N__6464\
        );

    \I__1150\ : Odrv12
    port map (
            O => \N__6464\,
            I => \un1_D_UU_AMIGA_1\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6461\,
            I => \N__6458\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6458\,
            I => \N__6455\
        );

    \I__1147\ : Span12Mux_v
    port map (
            O => \N__6455\,
            I => \N__6452\
        );

    \I__1146\ : Span12Mux_h
    port map (
            O => \N__6452\,
            I => \N__6449\
        );

    \I__1145\ : Odrv12
    port map (
            O => \N__6449\,
            I => \D_UM_040_in_3\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6442\
        );

    \I__1143\ : IoInMux
    port map (
            O => \N__6445\,
            I => \N__6439\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__6442\,
            I => \N__6436\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__6439\,
            I => \N__6433\
        );

    \I__1140\ : Span4Mux_v
    port map (
            O => \N__6436\,
            I => \N__6430\
        );

    \I__1139\ : Span4Mux_s3_h
    port map (
            O => \N__6433\,
            I => \N__6427\
        );

    \I__1138\ : Sp12to4
    port map (
            O => \N__6430\,
            I => \N__6424\
        );

    \I__1137\ : Sp12to4
    port map (
            O => \N__6427\,
            I => \N__6421\
        );

    \I__1136\ : Span12Mux_h
    port map (
            O => \N__6424\,
            I => \N__6418\
        );

    \I__1135\ : Span12Mux_v
    port map (
            O => \N__6421\,
            I => \N__6415\
        );

    \I__1134\ : Span12Mux_v
    port map (
            O => \N__6418\,
            I => \N__6412\
        );

    \I__1133\ : Span12Mux_h
    port map (
            O => \N__6415\,
            I => \N__6409\
        );

    \I__1132\ : Span12Mux_v
    port map (
            O => \N__6412\,
            I => \N__6404\
        );

    \I__1131\ : Span12Mux_h
    port map (
            O => \N__6409\,
            I => \N__6404\
        );

    \I__1130\ : Odrv12
    port map (
            O => \N__6404\,
            I => \D_LL_040_in_3\
        );

    \I__1129\ : IoInMux
    port map (
            O => \N__6401\,
            I => \N__6398\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6398\,
            I => \N__6395\
        );

    \I__1127\ : IoSpan4Mux
    port map (
            O => \N__6395\,
            I => \N__6392\
        );

    \I__1126\ : Span4Mux_s2_h
    port map (
            O => \N__6392\,
            I => \N__6389\
        );

    \I__1125\ : Sp12to4
    port map (
            O => \N__6389\,
            I => \N__6386\
        );

    \I__1124\ : Odrv12
    port map (
            O => \N__6386\,
            I => \un1_D_UM_040_3\
        );

    \I__1123\ : IoInMux
    port map (
            O => \N__6383\,
            I => \N__6380\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6380\,
            I => \N__6377\
        );

    \I__1121\ : IoSpan4Mux
    port map (
            O => \N__6377\,
            I => \N__6374\
        );

    \I__1120\ : IoSpan4Mux
    port map (
            O => \N__6374\,
            I => \N__6370\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6373\,
            I => \N__6367\
        );

    \I__1118\ : Span4Mux_s2_h
    port map (
            O => \N__6370\,
            I => \N__6364\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__6367\,
            I => \N__6361\
        );

    \I__1116\ : Sp12to4
    port map (
            O => \N__6364\,
            I => \N__6358\
        );

    \I__1115\ : Span12Mux_s10_v
    port map (
            O => \N__6361\,
            I => \N__6355\
        );

    \I__1114\ : Span12Mux_h
    port map (
            O => \N__6358\,
            I => \N__6350\
        );

    \I__1113\ : Span12Mux_v
    port map (
            O => \N__6355\,
            I => \N__6350\
        );

    \I__1112\ : Span12Mux_h
    port map (
            O => \N__6350\,
            I => \N__6347\
        );

    \I__1111\ : Odrv12
    port map (
            O => \N__6347\,
            I => \D_LM_040_in_3\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6344\,
            I => \N__6341\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6341\,
            I => \N__6338\
        );

    \I__1108\ : Span4Mux_v
    port map (
            O => \N__6338\,
            I => \N__6335\
        );

    \I__1107\ : Span4Mux_h
    port map (
            O => \N__6335\,
            I => \N__6332\
        );

    \I__1106\ : Sp12to4
    port map (
            O => \N__6332\,
            I => \N__6329\
        );

    \I__1105\ : Span12Mux_h
    port map (
            O => \N__6329\,
            I => \N__6326\
        );

    \I__1104\ : Odrv12
    port map (
            O => \N__6326\,
            I => \D_UU_040_in_3\
        );

    \I__1103\ : IoInMux
    port map (
            O => \N__6323\,
            I => \N__6320\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6320\,
            I => \N__6317\
        );

    \I__1101\ : Span12Mux_s6_v
    port map (
            O => \N__6317\,
            I => \N__6314\
        );

    \I__1100\ : Odrv12
    port map (
            O => \N__6314\,
            I => \un1_D_UU_040_3\
        );

    \I__1099\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6308\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__6308\,
            I => \U111_CYCLE_SM.N_124_0\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__6305\,
            I => \U111_CYCLE_SM.N_132_cascade_\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__6302\,
            I => \N__6299\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6299\,
            I => \N__6295\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6292\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6295\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__6292\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__6287\,
            I => \N__6284\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6284\,
            I => \N__6281\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__6281\,
            I => \N__6278\
        );

    \I__1088\ : Span4Mux_v
    port map (
            O => \N__6278\,
            I => \N__6275\
        );

    \I__1087\ : Span4Mux_v
    port map (
            O => \N__6275\,
            I => \N__6271\
        );

    \I__1086\ : IoInMux
    port map (
            O => \N__6274\,
            I => \N__6268\
        );

    \I__1085\ : Sp12to4
    port map (
            O => \N__6271\,
            I => \N__6265\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__6268\,
            I => \N__6262\
        );

    \I__1083\ : Span12Mux_h
    port map (
            O => \N__6265\,
            I => \N__6259\
        );

    \I__1082\ : IoSpan4Mux
    port map (
            O => \N__6262\,
            I => \N__6256\
        );

    \I__1081\ : Odrv12
    port map (
            O => \N__6259\,
            I => \TBIn_c\
        );

    \I__1080\ : Odrv4
    port map (
            O => \N__6256\,
            I => \TBIn_c\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6251\,
            I => \N__6248\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6248\,
            I => \U111_CYCLE_SM.un7_CYCLE_STATE_0\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__6245\,
            I => \U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__6242\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6239\,
            I => \N__6229\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6238\,
            I => \N__6229\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6237\,
            I => \N__6229\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6236\,
            I => \N__6225\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__6229\,
            I => \N__6222\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6228\,
            I => \N__6219\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6225\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__6222\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__6219\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__6212\,
            I => \N__6209\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6209\,
            I => \N__6203\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6208\,
            I => \N__6198\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6207\,
            I => \N__6198\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6206\,
            I => \N__6195\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__6203\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6198\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6195\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6188\,
            I => \N__6185\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6185\,
            I => \N__6177\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6174\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6183\,
            I => \N__6171\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6182\,
            I => \N__6164\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6164\
        );

    \I__1052\ : InMux
    port map (
            O => \N__6180\,
            I => \N__6164\
        );

    \I__1051\ : Odrv4
    port map (
            O => \N__6177\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6174\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6171\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__6164\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6155\,
            I => \N__6149\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6154\,
            I => \N__6149\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__6149\,
            I => \N__6146\
        );

    \I__1044\ : Sp12to4
    port map (
            O => \N__6146\,
            I => \N__6143\
        );

    \I__1043\ : Span12Mux_v
    port map (
            O => \N__6143\,
            I => \N__6140\
        );

    \I__1042\ : Span12Mux_h
    port map (
            O => \N__6140\,
            I => \N__6137\
        );

    \I__1041\ : Odrv12
    port map (
            O => \N__6137\,
            I => \SIZ_c_1\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__6134\,
            I => \N__6130\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__6133\,
            I => \N__6127\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6130\,
            I => \N__6122\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6127\,
            I => \N__6122\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6122\,
            I => \N__6119\
        );

    \I__1035\ : Span12Mux_v
    port map (
            O => \N__6119\,
            I => \N__6116\
        );

    \I__1034\ : Span12Mux_h
    port map (
            O => \N__6116\,
            I => \N__6113\
        );

    \I__1033\ : Odrv12
    port map (
            O => \N__6113\,
            I => \SIZ_c_0\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__6110\,
            I => \N__6107\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6107\,
            I => \N__6104\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6104\,
            I => \N__6101\
        );

    \I__1029\ : Span4Mux_v
    port map (
            O => \N__6101\,
            I => \N__6098\
        );

    \I__1028\ : Span4Mux_h
    port map (
            O => \N__6098\,
            I => \N__6095\
        );

    \I__1027\ : Odrv4
    port map (
            O => \N__6095\,
            I => \U111_CYCLE_SM.FLIP_WORD_2\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6089\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__6089\,
            I => \N__6085\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6081\
        );

    \I__1023\ : Span4Mux_v
    port map (
            O => \N__6085\,
            I => \N__6078\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6084\,
            I => \N__6075\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__6081\,
            I => \N__6072\
        );

    \I__1020\ : Sp12to4
    port map (
            O => \N__6078\,
            I => \N__6067\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6075\,
            I => \N__6067\
        );

    \I__1018\ : Span4Mux_h
    port map (
            O => \N__6072\,
            I => \N__6064\
        );

    \I__1017\ : Span12Mux_h
    port map (
            O => \N__6067\,
            I => \N__6061\
        );

    \I__1016\ : Span4Mux_v
    port map (
            O => \N__6064\,
            I => \N__6058\
        );

    \I__1015\ : Span12Mux_v
    port map (
            O => \N__6061\,
            I => \N__6055\
        );

    \I__1014\ : Span4Mux_v
    port map (
            O => \N__6058\,
            I => \N__6052\
        );

    \I__1013\ : Odrv12
    port map (
            O => \N__6055\,
            I => \PORTSIZE_c\
        );

    \I__1012\ : Odrv4
    port map (
            O => \N__6052\,
            I => \PORTSIZE_c\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6047\,
            I => \N__6040\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6046\,
            I => \N__6040\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6045\,
            I => \N__6037\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6040\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6037\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__1006\ : InMux
    port map (
            O => \N__6032\,
            I => \N__6029\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__6029\,
            I => \U111_CYCLE_SM.PORT_MISMATCH_2\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6026\,
            I => \N__6020\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6025\,
            I => \N__6020\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6020\,
            I => \N__6017\
        );

    \I__1001\ : Span4Mux_h
    port map (
            O => \N__6017\,
            I => \N__6014\
        );

    \I__1000\ : Sp12to4
    port map (
            O => \N__6014\,
            I => \N__6011\
        );

    \I__999\ : Span12Mux_v
    port map (
            O => \N__6011\,
            I => \N__6007\
        );

    \I__998\ : InMux
    port map (
            O => \N__6010\,
            I => \N__6004\
        );

    \I__997\ : Odrv12
    port map (
            O => \N__6007\,
            I => \U111_CYCLE_SM.A2_ENZ0\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__6004\,
            I => \U111_CYCLE_SM.A2_ENZ0\
        );

    \I__995\ : InMux
    port map (
            O => \N__5999\,
            I => \N__5996\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5996\,
            I => \N__5993\
        );

    \I__993\ : Span4Mux_v
    port map (
            O => \N__5993\,
            I => \N__5990\
        );

    \I__992\ : Sp12to4
    port map (
            O => \N__5990\,
            I => \N__5987\
        );

    \I__991\ : Odrv12
    port map (
            O => \N__5987\,
            I => \D_LM_AMIGA_in_5\
        );

    \I__990\ : IoInMux
    port map (
            O => \N__5984\,
            I => \N__5981\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__5981\,
            I => \N__5978\
        );

    \I__988\ : IoSpan4Mux
    port map (
            O => \N__5978\,
            I => \N__5975\
        );

    \I__987\ : Sp12to4
    port map (
            O => \N__5975\,
            I => \N__5972\
        );

    \I__986\ : Span12Mux_s7_h
    port map (
            O => \N__5972\,
            I => \N__5969\
        );

    \I__985\ : Span12Mux_h
    port map (
            O => \N__5969\,
            I => \N__5966\
        );

    \I__984\ : Odrv12
    port map (
            O => \N__5966\,
            I => \un2_D_LM_AMIGA_5\
        );

    \I__983\ : IoInMux
    port map (
            O => \N__5963\,
            I => \N__5960\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5960\,
            I => \N__5956\
        );

    \I__981\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5953\
        );

    \I__980\ : IoSpan4Mux
    port map (
            O => \N__5956\,
            I => \N__5950\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__5953\,
            I => \N__5947\
        );

    \I__978\ : Span4Mux_s2_h
    port map (
            O => \N__5950\,
            I => \N__5944\
        );

    \I__977\ : Sp12to4
    port map (
            O => \N__5947\,
            I => \N__5941\
        );

    \I__976\ : Span4Mux_v
    port map (
            O => \N__5944\,
            I => \N__5938\
        );

    \I__975\ : Span12Mux_v
    port map (
            O => \N__5941\,
            I => \N__5935\
        );

    \I__974\ : Sp12to4
    port map (
            O => \N__5938\,
            I => \N__5932\
        );

    \I__973\ : Span12Mux_v
    port map (
            O => \N__5935\,
            I => \N__5929\
        );

    \I__972\ : Span12Mux_s9_h
    port map (
            O => \N__5932\,
            I => \N__5926\
        );

    \I__971\ : Span12Mux_h
    port map (
            O => \N__5929\,
            I => \N__5923\
        );

    \I__970\ : Span12Mux_h
    port map (
            O => \N__5926\,
            I => \N__5920\
        );

    \I__969\ : Odrv12
    port map (
            O => \N__5923\,
            I => \D_LM_040_in_0\
        );

    \I__968\ : Odrv12
    port map (
            O => \N__5920\,
            I => \D_LM_040_in_0\
        );

    \I__967\ : InMux
    port map (
            O => \N__5915\,
            I => \N__5912\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5912\,
            I => \N__5909\
        );

    \I__965\ : Span4Mux_v
    port map (
            O => \N__5909\,
            I => \N__5906\
        );

    \I__964\ : Span4Mux_h
    port map (
            O => \N__5906\,
            I => \N__5903\
        );

    \I__963\ : Sp12to4
    port map (
            O => \N__5903\,
            I => \N__5900\
        );

    \I__962\ : Span12Mux_h
    port map (
            O => \N__5900\,
            I => \N__5897\
        );

    \I__961\ : Odrv12
    port map (
            O => \N__5897\,
            I => \D_UU_040_in_0\
        );

    \I__960\ : IoInMux
    port map (
            O => \N__5894\,
            I => \N__5891\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__5891\,
            I => \N__5888\
        );

    \I__958\ : Span12Mux_s6_v
    port map (
            O => \N__5888\,
            I => \N__5885\
        );

    \I__957\ : Odrv12
    port map (
            O => \N__5885\,
            I => \un1_D_UU_040_0\
        );

    \I__956\ : InMux
    port map (
            O => \N__5882\,
            I => \N__5879\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5879\,
            I => \N__5876\
        );

    \I__954\ : Span4Mux_v
    port map (
            O => \N__5876\,
            I => \N__5873\
        );

    \I__953\ : Span4Mux_h
    port map (
            O => \N__5873\,
            I => \N__5870\
        );

    \I__952\ : Sp12to4
    port map (
            O => \N__5870\,
            I => \N__5867\
        );

    \I__951\ : Odrv12
    port map (
            O => \N__5867\,
            I => \D_LL_AMIGA_in_6\
        );

    \I__950\ : IoInMux
    port map (
            O => \N__5864\,
            I => \N__5861\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5861\,
            I => \N__5858\
        );

    \I__948\ : Span4Mux_s3_h
    port map (
            O => \N__5858\,
            I => \N__5855\
        );

    \I__947\ : Span4Mux_v
    port map (
            O => \N__5855\,
            I => \N__5852\
        );

    \I__946\ : Span4Mux_v
    port map (
            O => \N__5852\,
            I => \N__5849\
        );

    \I__945\ : Sp12to4
    port map (
            O => \N__5849\,
            I => \N__5846\
        );

    \I__944\ : Span12Mux_s10_h
    port map (
            O => \N__5846\,
            I => \N__5843\
        );

    \I__943\ : Odrv12
    port map (
            O => \N__5843\,
            I => \un2_D_LL_AMIGA_6\
        );

    \I__942\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5837\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5837\,
            I => \N__5834\
        );

    \I__940\ : Span4Mux_v
    port map (
            O => \N__5834\,
            I => \N__5831\
        );

    \I__939\ : Span4Mux_h
    port map (
            O => \N__5831\,
            I => \N__5828\
        );

    \I__938\ : Sp12to4
    port map (
            O => \N__5828\,
            I => \N__5825\
        );

    \I__937\ : Span12Mux_h
    port map (
            O => \N__5825\,
            I => \N__5822\
        );

    \I__936\ : Odrv12
    port map (
            O => \N__5822\,
            I => \D_UU_040_in_6\
        );

    \I__935\ : IoInMux
    port map (
            O => \N__5819\,
            I => \N__5816\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5816\,
            I => \N__5812\
        );

    \I__933\ : InMux
    port map (
            O => \N__5815\,
            I => \N__5809\
        );

    \I__932\ : Span4Mux_s2_h
    port map (
            O => \N__5812\,
            I => \N__5806\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5809\,
            I => \N__5803\
        );

    \I__930\ : Span4Mux_v
    port map (
            O => \N__5806\,
            I => \N__5800\
        );

    \I__929\ : Span4Mux_v
    port map (
            O => \N__5803\,
            I => \N__5797\
        );

    \I__928\ : Sp12to4
    port map (
            O => \N__5800\,
            I => \N__5794\
        );

    \I__927\ : Span4Mux_v
    port map (
            O => \N__5797\,
            I => \N__5791\
        );

    \I__926\ : Span12Mux_h
    port map (
            O => \N__5794\,
            I => \N__5786\
        );

    \I__925\ : Sp12to4
    port map (
            O => \N__5791\,
            I => \N__5786\
        );

    \I__924\ : Span12Mux_h
    port map (
            O => \N__5786\,
            I => \N__5783\
        );

    \I__923\ : Odrv12
    port map (
            O => \N__5783\,
            I => \D_LM_040_in_6\
        );

    \I__922\ : IoInMux
    port map (
            O => \N__5780\,
            I => \N__5777\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__5777\,
            I => \N__5774\
        );

    \I__920\ : Span4Mux_s3_v
    port map (
            O => \N__5774\,
            I => \N__5771\
        );

    \I__919\ : Span4Mux_h
    port map (
            O => \N__5771\,
            I => \N__5768\
        );

    \I__918\ : Span4Mux_h
    port map (
            O => \N__5768\,
            I => \N__5765\
        );

    \I__917\ : Odrv4
    port map (
            O => \N__5765\,
            I => \un1_D_UU_040_6\
        );

    \I__916\ : InMux
    port map (
            O => \N__5762\,
            I => \N__5759\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__5759\,
            I => \N__5756\
        );

    \I__914\ : Span4Mux_v
    port map (
            O => \N__5756\,
            I => \N__5753\
        );

    \I__913\ : Sp12to4
    port map (
            O => \N__5753\,
            I => \N__5750\
        );

    \I__912\ : Odrv12
    port map (
            O => \N__5750\,
            I => \D_LL_AMIGA_in_3\
        );

    \I__911\ : IoInMux
    port map (
            O => \N__5747\,
            I => \N__5744\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__5744\,
            I => \N__5741\
        );

    \I__909\ : Span12Mux_s7_h
    port map (
            O => \N__5741\,
            I => \N__5738\
        );

    \I__908\ : Span12Mux_h
    port map (
            O => \N__5738\,
            I => \N__5735\
        );

    \I__907\ : Odrv12
    port map (
            O => \N__5735\,
            I => \un2_D_LL_AMIGA_3\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__5732\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa_cascade_\
        );

    \I__905\ : InMux
    port map (
            O => \N__5729\,
            I => \N__5725\
        );

    \I__904\ : InMux
    port map (
            O => \N__5728\,
            I => \N__5722\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5725\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_0\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5722\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_0\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__5717\,
            I => \N__5714\
        );

    \I__900\ : InMux
    port map (
            O => \N__5714\,
            I => \N__5711\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__5711\,
            I => \U111_CYCLE_SM.TS_EN_6\
        );

    \I__898\ : IoInMux
    port map (
            O => \N__5708\,
            I => \N__5704\
        );

    \I__897\ : IoInMux
    port map (
            O => \N__5707\,
            I => \N__5701\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5704\,
            I => \N__5698\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__5701\,
            I => \N__5695\
        );

    \I__894\ : Span12Mux_s6_v
    port map (
            O => \N__5698\,
            I => \N__5690\
        );

    \I__893\ : Span12Mux_s6_v
    port map (
            O => \N__5695\,
            I => \N__5690\
        );

    \I__892\ : Odrv12
    port map (
            O => \N__5690\,
            I => \CONSTANT_ONE_NET\
        );

    \I__891\ : InMux
    port map (
            O => \N__5687\,
            I => \N__5684\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5684\,
            I => \N__5681\
        );

    \I__889\ : Span4Mux_v
    port map (
            O => \N__5681\,
            I => \N__5678\
        );

    \I__888\ : Sp12to4
    port map (
            O => \N__5678\,
            I => \N__5675\
        );

    \I__887\ : Span12Mux_h
    port map (
            O => \N__5675\,
            I => \N__5672\
        );

    \I__886\ : Odrv12
    port map (
            O => \N__5672\,
            I => \D_LL_AMIGA_in_2\
        );

    \I__885\ : IoInMux
    port map (
            O => \N__5669\,
            I => \N__5666\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5666\,
            I => \N__5663\
        );

    \I__883\ : Span4Mux_s2_h
    port map (
            O => \N__5663\,
            I => \N__5660\
        );

    \I__882\ : Sp12to4
    port map (
            O => \N__5660\,
            I => \N__5657\
        );

    \I__881\ : Span12Mux_s8_v
    port map (
            O => \N__5657\,
            I => \N__5654\
        );

    \I__880\ : Span12Mux_h
    port map (
            O => \N__5654\,
            I => \N__5651\
        );

    \I__879\ : Odrv12
    port map (
            O => \N__5651\,
            I => \un2_D_LL_AMIGA_2\
        );

    \I__878\ : InMux
    port map (
            O => \N__5648\,
            I => \N__5645\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5645\,
            I => \N__5642\
        );

    \I__876\ : Span4Mux_v
    port map (
            O => \N__5642\,
            I => \N__5639\
        );

    \I__875\ : Sp12to4
    port map (
            O => \N__5639\,
            I => \N__5636\
        );

    \I__874\ : Span12Mux_h
    port map (
            O => \N__5636\,
            I => \N__5633\
        );

    \I__873\ : Odrv12
    port map (
            O => \N__5633\,
            I => \D_LM_AMIGA_in_0\
        );

    \I__872\ : IoInMux
    port map (
            O => \N__5630\,
            I => \N__5627\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5627\,
            I => \N__5624\
        );

    \I__870\ : IoSpan4Mux
    port map (
            O => \N__5624\,
            I => \N__5621\
        );

    \I__869\ : Span4Mux_s3_h
    port map (
            O => \N__5621\,
            I => \N__5618\
        );

    \I__868\ : Sp12to4
    port map (
            O => \N__5618\,
            I => \N__5615\
        );

    \I__867\ : Span12Mux_s8_h
    port map (
            O => \N__5615\,
            I => \N__5612\
        );

    \I__866\ : Span12Mux_h
    port map (
            O => \N__5612\,
            I => \N__5609\
        );

    \I__865\ : Odrv12
    port map (
            O => \N__5609\,
            I => \un2_D_LM_AMIGA_0\
        );

    \I__864\ : IoInMux
    port map (
            O => \N__5606\,
            I => \N__5603\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5603\,
            I => \N__5600\
        );

    \I__862\ : Span12Mux_s5_v
    port map (
            O => \N__5600\,
            I => \N__5597\
        );

    \I__861\ : Odrv12
    port map (
            O => \N__5597\,
            I => \TSn_c\
        );

    \I__860\ : InMux
    port map (
            O => \N__5594\,
            I => \N__5590\
        );

    \I__859\ : InMux
    port map (
            O => \N__5593\,
            I => \N__5587\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5590\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__5587\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__856\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__854\ : Span4Mux_v
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__853\ : Sp12to4
    port map (
            O => \N__5573\,
            I => \N__5570\
        );

    \I__852\ : Span12Mux_h
    port map (
            O => \N__5570\,
            I => \N__5567\
        );

    \I__851\ : Span12Mux_v
    port map (
            O => \N__5567\,
            I => \N__5564\
        );

    \I__850\ : Odrv12
    port map (
            O => \N__5564\,
            I => \D_UM_040_in_1\
        );

    \I__849\ : IoInMux
    port map (
            O => \N__5561\,
            I => \N__5558\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__5558\,
            I => \N__5554\
        );

    \I__847\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5551\
        );

    \I__846\ : Span4Mux_s3_h
    port map (
            O => \N__5554\,
            I => \N__5548\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5551\,
            I => \N__5545\
        );

    \I__844\ : Sp12to4
    port map (
            O => \N__5548\,
            I => \N__5542\
        );

    \I__843\ : Span12Mux_v
    port map (
            O => \N__5545\,
            I => \N__5539\
        );

    \I__842\ : Span12Mux_v
    port map (
            O => \N__5542\,
            I => \N__5536\
        );

    \I__841\ : Span12Mux_v
    port map (
            O => \N__5539\,
            I => \N__5533\
        );

    \I__840\ : Span12Mux_h
    port map (
            O => \N__5536\,
            I => \N__5530\
        );

    \I__839\ : Span12Mux_h
    port map (
            O => \N__5533\,
            I => \N__5527\
        );

    \I__838\ : Span12Mux_h
    port map (
            O => \N__5530\,
            I => \N__5524\
        );

    \I__837\ : Odrv12
    port map (
            O => \N__5527\,
            I => \D_LL_040_in_1\
        );

    \I__836\ : Odrv12
    port map (
            O => \N__5524\,
            I => \D_LL_040_in_1\
        );

    \I__835\ : IoInMux
    port map (
            O => \N__5519\,
            I => \N__5516\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5516\,
            I => \N__5513\
        );

    \I__833\ : Span4Mux_s3_h
    port map (
            O => \N__5513\,
            I => \N__5510\
        );

    \I__832\ : Span4Mux_h
    port map (
            O => \N__5510\,
            I => \N__5507\
        );

    \I__831\ : Span4Mux_h
    port map (
            O => \N__5507\,
            I => \N__5504\
        );

    \I__830\ : Odrv4
    port map (
            O => \N__5504\,
            I => \un1_D_UM_040_1\
        );

    \I__829\ : InMux
    port map (
            O => \N__5501\,
            I => \N__5498\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5498\,
            I => \N__5495\
        );

    \I__827\ : Span4Mux_v
    port map (
            O => \N__5495\,
            I => \N__5492\
        );

    \I__826\ : Sp12to4
    port map (
            O => \N__5492\,
            I => \N__5489\
        );

    \I__825\ : Span12Mux_h
    port map (
            O => \N__5489\,
            I => \N__5486\
        );

    \I__824\ : Odrv12
    port map (
            O => \N__5486\,
            I => \D_LM_AMIGA_in_6\
        );

    \I__823\ : IoInMux
    port map (
            O => \N__5483\,
            I => \N__5480\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5480\,
            I => \N__5477\
        );

    \I__821\ : IoSpan4Mux
    port map (
            O => \N__5477\,
            I => \N__5474\
        );

    \I__820\ : Sp12to4
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__819\ : Span12Mux_s9_h
    port map (
            O => \N__5471\,
            I => \N__5468\
        );

    \I__818\ : Odrv12
    port map (
            O => \N__5468\,
            I => \un2_D_LM_AMIGA_6\
        );

    \I__817\ : IoInMux
    port map (
            O => \N__5465\,
            I => \N__5462\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5462\,
            I => \N__5459\
        );

    \I__815\ : Span4Mux_s3_h
    port map (
            O => \N__5459\,
            I => \N__5456\
        );

    \I__814\ : Span4Mux_h
    port map (
            O => \N__5456\,
            I => \N__5452\
        );

    \I__813\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5449\
        );

    \I__812\ : Span4Mux_h
    port map (
            O => \N__5452\,
            I => \N__5446\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5449\,
            I => \N__5443\
        );

    \I__810\ : Sp12to4
    port map (
            O => \N__5446\,
            I => \N__5438\
        );

    \I__809\ : Span12Mux_v
    port map (
            O => \N__5443\,
            I => \N__5438\
        );

    \I__808\ : Span12Mux_v
    port map (
            O => \N__5438\,
            I => \N__5435\
        );

    \I__807\ : Span12Mux_h
    port map (
            O => \N__5435\,
            I => \N__5432\
        );

    \I__806\ : Odrv12
    port map (
            O => \N__5432\,
            I => \D_LM_040_in_1\
        );

    \I__805\ : InMux
    port map (
            O => \N__5429\,
            I => \N__5426\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5426\,
            I => \N__5423\
        );

    \I__803\ : Span12Mux_v
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__802\ : Span12Mux_h
    port map (
            O => \N__5420\,
            I => \N__5417\
        );

    \I__801\ : Odrv12
    port map (
            O => \N__5417\,
            I => \D_UU_040_in_1\
        );

    \I__800\ : IoInMux
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__5411\,
            I => \N__5408\
        );

    \I__798\ : Span4Mux_s3_h
    port map (
            O => \N__5408\,
            I => \N__5405\
        );

    \I__797\ : Span4Mux_h
    port map (
            O => \N__5405\,
            I => \N__5402\
        );

    \I__796\ : Span4Mux_h
    port map (
            O => \N__5402\,
            I => \N__5399\
        );

    \I__795\ : Odrv4
    port map (
            O => \N__5399\,
            I => \un1_D_UU_040_1\
        );

    \I__794\ : IoInMux
    port map (
            O => \N__5396\,
            I => \N__5392\
        );

    \I__793\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5389\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5392\,
            I => \N__5386\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__5389\,
            I => \N__5383\
        );

    \I__790\ : IoSpan4Mux
    port map (
            O => \N__5386\,
            I => \N__5380\
        );

    \I__789\ : Span4Mux_v
    port map (
            O => \N__5383\,
            I => \N__5377\
        );

    \I__788\ : Span4Mux_s2_h
    port map (
            O => \N__5380\,
            I => \N__5374\
        );

    \I__787\ : Sp12to4
    port map (
            O => \N__5377\,
            I => \N__5371\
        );

    \I__786\ : Span4Mux_v
    port map (
            O => \N__5374\,
            I => \N__5368\
        );

    \I__785\ : Span12Mux_h
    port map (
            O => \N__5371\,
            I => \N__5365\
        );

    \I__784\ : Sp12to4
    port map (
            O => \N__5368\,
            I => \N__5362\
        );

    \I__783\ : Span12Mux_v
    port map (
            O => \N__5365\,
            I => \N__5359\
        );

    \I__782\ : Span12Mux_h
    port map (
            O => \N__5362\,
            I => \N__5356\
        );

    \I__781\ : Span12Mux_v
    port map (
            O => \N__5359\,
            I => \N__5353\
        );

    \I__780\ : Span12Mux_h
    port map (
            O => \N__5356\,
            I => \N__5350\
        );

    \I__779\ : Odrv12
    port map (
            O => \N__5353\,
            I => \D_LL_040_in_5\
        );

    \I__778\ : Odrv12
    port map (
            O => \N__5350\,
            I => \D_LL_040_in_5\
        );

    \I__777\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5342\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__5342\,
            I => \N__5339\
        );

    \I__775\ : Span4Mux_v
    port map (
            O => \N__5339\,
            I => \N__5336\
        );

    \I__774\ : Span4Mux_h
    port map (
            O => \N__5336\,
            I => \N__5333\
        );

    \I__773\ : Sp12to4
    port map (
            O => \N__5333\,
            I => \N__5330\
        );

    \I__772\ : Span12Mux_h
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__771\ : Odrv12
    port map (
            O => \N__5327\,
            I => \D_UM_040_in_5\
        );

    \I__770\ : IoInMux
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5321\,
            I => \N__5318\
        );

    \I__768\ : IoSpan4Mux
    port map (
            O => \N__5318\,
            I => \N__5315\
        );

    \I__767\ : Span4Mux_s2_v
    port map (
            O => \N__5315\,
            I => \N__5312\
        );

    \I__766\ : Span4Mux_h
    port map (
            O => \N__5312\,
            I => \N__5309\
        );

    \I__765\ : Span4Mux_v
    port map (
            O => \N__5309\,
            I => \N__5306\
        );

    \I__764\ : Odrv4
    port map (
            O => \N__5306\,
            I => \un1_D_UM_040_5\
        );

    \I__763\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5300\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__5300\,
            I => \WRITE_CYCLE_ACTIVE_rep13_i_ess\
        );

    \I__761\ : InMux
    port map (
            O => \N__5297\,
            I => \N__5294\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__5294\,
            I => \WRITE_CYCLE_ACTIVE_rep4_i_ess\
        );

    \I__759\ : IoInMux
    port map (
            O => \N__5291\,
            I => \N__5288\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5288\,
            I => \N__5285\
        );

    \I__757\ : IoSpan4Mux
    port map (
            O => \N__5285\,
            I => \N__5282\
        );

    \I__756\ : Span4Mux_s3_v
    port map (
            O => \N__5282\,
            I => \N__5279\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__5279\,
            I => \N_217_i\
        );

    \I__754\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5273\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5273\,
            I => \N__5270\
        );

    \I__752\ : Span4Mux_v
    port map (
            O => \N__5270\,
            I => \N__5267\
        );

    \I__751\ : Sp12to4
    port map (
            O => \N__5267\,
            I => \N__5264\
        );

    \I__750\ : Odrv12
    port map (
            O => \N__5264\,
            I => \D_LL_AMIGA_in_4\
        );

    \I__749\ : IoInMux
    port map (
            O => \N__5261\,
            I => \N__5258\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__747\ : Span4Mux_s2_h
    port map (
            O => \N__5255\,
            I => \N__5252\
        );

    \I__746\ : Sp12to4
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__745\ : Span12Mux_s8_v
    port map (
            O => \N__5249\,
            I => \N__5246\
        );

    \I__744\ : Span12Mux_h
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__743\ : Odrv12
    port map (
            O => \N__5243\,
            I => \un2_D_LL_AMIGA_4\
        );

    \I__742\ : IoInMux
    port map (
            O => \N__5240\,
            I => \N__5236\
        );

    \I__741\ : InMux
    port map (
            O => \N__5239\,
            I => \N__5233\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5236\,
            I => \N__5230\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5233\,
            I => \N__5227\
        );

    \I__738\ : IoSpan4Mux
    port map (
            O => \N__5230\,
            I => \N__5224\
        );

    \I__737\ : Span4Mux_v
    port map (
            O => \N__5227\,
            I => \N__5221\
        );

    \I__736\ : Span4Mux_s2_h
    port map (
            O => \N__5224\,
            I => \N__5218\
        );

    \I__735\ : Sp12to4
    port map (
            O => \N__5221\,
            I => \N__5215\
        );

    \I__734\ : Sp12to4
    port map (
            O => \N__5218\,
            I => \N__5212\
        );

    \I__733\ : Span12Mux_h
    port map (
            O => \N__5215\,
            I => \N__5209\
        );

    \I__732\ : Span12Mux_h
    port map (
            O => \N__5212\,
            I => \N__5206\
        );

    \I__731\ : Span12Mux_v
    port map (
            O => \N__5209\,
            I => \N__5203\
        );

    \I__730\ : Span12Mux_h
    port map (
            O => \N__5206\,
            I => \N__5200\
        );

    \I__729\ : Odrv12
    port map (
            O => \N__5203\,
            I => \D_LL_040_in_0\
        );

    \I__728\ : Odrv12
    port map (
            O => \N__5200\,
            I => \D_LL_040_in_0\
        );

    \I__727\ : InMux
    port map (
            O => \N__5195\,
            I => \N__5192\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5192\,
            I => \N__5189\
        );

    \I__725\ : Span12Mux_h
    port map (
            O => \N__5189\,
            I => \N__5186\
        );

    \I__724\ : Span12Mux_h
    port map (
            O => \N__5186\,
            I => \N__5183\
        );

    \I__723\ : Odrv12
    port map (
            O => \N__5183\,
            I => \D_UM_040_in_0\
        );

    \I__722\ : IoInMux
    port map (
            O => \N__5180\,
            I => \N__5177\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__5177\,
            I => \N__5174\
        );

    \I__720\ : IoSpan4Mux
    port map (
            O => \N__5174\,
            I => \N__5171\
        );

    \I__719\ : Span4Mux_s1_h
    port map (
            O => \N__5171\,
            I => \N__5168\
        );

    \I__718\ : Span4Mux_h
    port map (
            O => \N__5168\,
            I => \N__5165\
        );

    \I__717\ : Span4Mux_h
    port map (
            O => \N__5165\,
            I => \N__5162\
        );

    \I__716\ : Odrv4
    port map (
            O => \N__5162\,
            I => \un1_D_UM_040_0\
        );

    \I__715\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5156\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__5156\,
            I => \N__5153\
        );

    \I__713\ : Span12Mux_h
    port map (
            O => \N__5153\,
            I => \N__5150\
        );

    \I__712\ : Odrv12
    port map (
            O => \N__5150\,
            I => \D_LM_AMIGA_in_3\
        );

    \I__711\ : IoInMux
    port map (
            O => \N__5147\,
            I => \N__5144\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5144\,
            I => \N__5141\
        );

    \I__709\ : IoSpan4Mux
    port map (
            O => \N__5141\,
            I => \N__5138\
        );

    \I__708\ : Span4Mux_s0_h
    port map (
            O => \N__5138\,
            I => \N__5135\
        );

    \I__707\ : Sp12to4
    port map (
            O => \N__5135\,
            I => \N__5132\
        );

    \I__706\ : Span12Mux_s9_h
    port map (
            O => \N__5132\,
            I => \N__5129\
        );

    \I__705\ : Span12Mux_h
    port map (
            O => \N__5129\,
            I => \N__5126\
        );

    \I__704\ : Odrv12
    port map (
            O => \N__5126\,
            I => \un2_D_LM_AMIGA_3\
        );

    \I__703\ : IoInMux
    port map (
            O => \N__5123\,
            I => \N__5120\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5120\,
            I => \N__5117\
        );

    \I__701\ : IoSpan4Mux
    port map (
            O => \N__5117\,
            I => \N__5114\
        );

    \I__700\ : Span4Mux_s2_v
    port map (
            O => \N__5114\,
            I => \N__5111\
        );

    \I__699\ : Span4Mux_v
    port map (
            O => \N__5111\,
            I => \N__5108\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__5108\,
            I => \LBENn_c_i\
        );

    \I__697\ : InMux
    port map (
            O => \N__5105\,
            I => \N__5102\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5102\,
            I => \WRITE_CYCLE_ACTIVE_rep2_i_ess\
        );

    \I__695\ : IoInMux
    port map (
            O => \N__5099\,
            I => \N__5096\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__5096\,
            I => \N__5093\
        );

    \I__693\ : Span4Mux_s2_v
    port map (
            O => \N__5093\,
            I => \N__5090\
        );

    \I__692\ : Span4Mux_h
    port map (
            O => \N__5090\,
            I => \N__5087\
        );

    \I__691\ : Span4Mux_v
    port map (
            O => \N__5087\,
            I => \N__5084\
        );

    \I__690\ : Odrv4
    port map (
            O => \N__5084\,
            I => \N_215_i\
        );

    \I__689\ : InMux
    port map (
            O => \N__5081\,
            I => \N__5078\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__5078\,
            I => \N__5075\
        );

    \I__687\ : Span4Mux_v
    port map (
            O => \N__5075\,
            I => \N__5072\
        );

    \I__686\ : Sp12to4
    port map (
            O => \N__5072\,
            I => \N__5069\
        );

    \I__685\ : Span12Mux_h
    port map (
            O => \N__5069\,
            I => \N__5066\
        );

    \I__684\ : Odrv12
    port map (
            O => \N__5066\,
            I => \D_UM_040_in_6\
        );

    \I__683\ : IoInMux
    port map (
            O => \N__5063\,
            I => \N__5060\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5060\,
            I => \N__5057\
        );

    \I__681\ : IoSpan4Mux
    port map (
            O => \N__5057\,
            I => \N__5054\
        );

    \I__680\ : Span4Mux_s1_h
    port map (
            O => \N__5054\,
            I => \N__5050\
        );

    \I__679\ : InMux
    port map (
            O => \N__5053\,
            I => \N__5047\
        );

    \I__678\ : Span4Mux_h
    port map (
            O => \N__5050\,
            I => \N__5044\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5047\,
            I => \N__5041\
        );

    \I__676\ : Span4Mux_h
    port map (
            O => \N__5044\,
            I => \N__5036\
        );

    \I__675\ : Span4Mux_v
    port map (
            O => \N__5041\,
            I => \N__5036\
        );

    \I__674\ : Sp12to4
    port map (
            O => \N__5036\,
            I => \N__5033\
        );

    \I__673\ : Span12Mux_v
    port map (
            O => \N__5033\,
            I => \N__5030\
        );

    \I__672\ : Span12Mux_h
    port map (
            O => \N__5030\,
            I => \N__5027\
        );

    \I__671\ : Odrv12
    port map (
            O => \N__5027\,
            I => \D_LL_040_in_6\
        );

    \I__670\ : IoInMux
    port map (
            O => \N__5024\,
            I => \N__5021\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5021\,
            I => \N__5018\
        );

    \I__668\ : Span12Mux_s2_h
    port map (
            O => \N__5018\,
            I => \N__5015\
        );

    \I__667\ : Span12Mux_v
    port map (
            O => \N__5015\,
            I => \N__5012\
        );

    \I__666\ : Odrv12
    port map (
            O => \N__5012\,
            I => \un1_D_UM_040_6\
        );

    \I__665\ : InMux
    port map (
            O => \N__5009\,
            I => \N__5006\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__5006\,
            I => \N__5003\
        );

    \I__663\ : Odrv12
    port map (
            O => \N__5003\,
            I => \D_LM_AMIGA_in_2\
        );

    \I__662\ : IoInMux
    port map (
            O => \N__5000\,
            I => \N__4997\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4997\,
            I => \N__4994\
        );

    \I__660\ : Sp12to4
    port map (
            O => \N__4994\,
            I => \N__4991\
        );

    \I__659\ : Span12Mux_h
    port map (
            O => \N__4991\,
            I => \N__4988\
        );

    \I__658\ : Span12Mux_v
    port map (
            O => \N__4988\,
            I => \N__4985\
        );

    \I__657\ : Odrv12
    port map (
            O => \N__4985\,
            I => \un2_D_LM_AMIGA_2\
        );

    \I__656\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__4979\,
            I => \WRITE_CYCLE_ACTIVE_rep0_i_ess\
        );

    \I__654\ : IoInMux
    port map (
            O => \N__4976\,
            I => \N__4973\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4973\,
            I => \N__4970\
        );

    \I__652\ : Span4Mux_s3_v
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__651\ : Span4Mux_v
    port map (
            O => \N__4967\,
            I => \N__4964\
        );

    \I__650\ : Odrv4
    port map (
            O => \N__4964\,
            I => \N_213_i\
        );

    \I__649\ : IoInMux
    port map (
            O => \N__4961\,
            I => \N__4958\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4958\,
            I => \N__4955\
        );

    \I__647\ : Span4Mux_s3_v
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__646\ : Span4Mux_h
    port map (
            O => \N__4952\,
            I => \N__4949\
        );

    \I__645\ : Span4Mux_v
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__644\ : Odrv4
    port map (
            O => \N__4946\,
            I => \N_226_i\
        );

    \I__643\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4940\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__4940\,
            I => \N__4937\
        );

    \I__641\ : Odrv4
    port map (
            O => \N__4937\,
            I => \WRITE_CYCLE_ACTIVE_rep6_i_ess\
        );

    \I__640\ : InMux
    port map (
            O => \N__4934\,
            I => \N__4931\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4931\,
            I => \N__4928\
        );

    \I__638\ : Span12Mux_v
    port map (
            O => \N__4928\,
            I => \N__4925\
        );

    \I__637\ : Odrv12
    port map (
            O => \N__4925\,
            I => \D_LL_AMIGA_in_1\
        );

    \I__636\ : IoInMux
    port map (
            O => \N__4922\,
            I => \N__4919\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4919\,
            I => \N__4916\
        );

    \I__634\ : Span4Mux_s3_h
    port map (
            O => \N__4916\,
            I => \N__4913\
        );

    \I__633\ : Sp12to4
    port map (
            O => \N__4913\,
            I => \N__4910\
        );

    \I__632\ : Span12Mux_s8_v
    port map (
            O => \N__4910\,
            I => \N__4907\
        );

    \I__631\ : Span12Mux_h
    port map (
            O => \N__4907\,
            I => \N__4904\
        );

    \I__630\ : Odrv12
    port map (
            O => \N__4904\,
            I => \un2_D_LL_AMIGA_1\
        );

    \I__629\ : InMux
    port map (
            O => \N__4901\,
            I => \N__4898\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__4898\,
            I => \N__4895\
        );

    \I__627\ : Span4Mux_v
    port map (
            O => \N__4895\,
            I => \N__4892\
        );

    \I__626\ : Span4Mux_v
    port map (
            O => \N__4892\,
            I => \N__4888\
        );

    \I__625\ : InMux
    port map (
            O => \N__4891\,
            I => \N__4885\
        );

    \I__624\ : Sp12to4
    port map (
            O => \N__4888\,
            I => \N__4880\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__4885\,
            I => \N__4880\
        );

    \I__622\ : Span12Mux_h
    port map (
            O => \N__4880\,
            I => \N__4877\
        );

    \I__621\ : Odrv12
    port map (
            O => \N__4877\,
            I => \A_040_c_1\
        );

    \I__620\ : InMux
    port map (
            O => \N__4874\,
            I => \N__4871\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4871\,
            I => \N__4868\
        );

    \I__618\ : Odrv4
    port map (
            O => \N__4868\,
            I => \WRITE_CYCLE_ACTIVE_rep21_i_ess\
        );

    \I__617\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4862\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4862\,
            I => \N__4859\
        );

    \I__615\ : Span4Mux_v
    port map (
            O => \N__4859\,
            I => \N__4856\
        );

    \I__614\ : Odrv4
    port map (
            O => \N__4856\,
            I => \WRITE_CYCLE_ACTIVE_rep23_i_ess\
        );

    \I__613\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4850\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4850\,
            I => \WRITE_CYCLE_ACTIVE_rep7_i_ess\
        );

    \I__611\ : IoInMux
    port map (
            O => \N__4847\,
            I => \N__4844\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4844\,
            I => \N__4841\
        );

    \I__609\ : IoSpan4Mux
    port map (
            O => \N__4841\,
            I => \N__4838\
        );

    \I__608\ : Span4Mux_s2_v
    port map (
            O => \N__4838\,
            I => \N__4835\
        );

    \I__607\ : Span4Mux_v
    port map (
            O => \N__4835\,
            I => \N__4832\
        );

    \I__606\ : Odrv4
    port map (
            O => \N__4832\,
            I => \N_220_i\
        );

    \I__605\ : InMux
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4826\,
            I => \WRITE_CYCLE_ACTIVE_rep3_i_ess\
        );

    \I__603\ : IoInMux
    port map (
            O => \N__4823\,
            I => \N__4820\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4820\,
            I => \N__4817\
        );

    \I__601\ : IoSpan4Mux
    port map (
            O => \N__4817\,
            I => \N__4814\
        );

    \I__600\ : Span4Mux_s3_v
    port map (
            O => \N__4814\,
            I => \N__4811\
        );

    \I__599\ : Odrv4
    port map (
            O => \N__4811\,
            I => \N_219_i\
        );

    \I__598\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4805\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4805\,
            I => \N__4802\
        );

    \I__596\ : Span4Mux_v
    port map (
            O => \N__4802\,
            I => \N__4799\
        );

    \I__595\ : Sp12to4
    port map (
            O => \N__4799\,
            I => \N__4796\
        );

    \I__594\ : Odrv12
    port map (
            O => \N__4796\,
            I => \D_LL_AMIGA_in_0\
        );

    \I__593\ : IoInMux
    port map (
            O => \N__4793\,
            I => \N__4790\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4790\,
            I => \N__4787\
        );

    \I__591\ : Span12Mux_s11_h
    port map (
            O => \N__4787\,
            I => \N__4784\
        );

    \I__590\ : Span12Mux_h
    port map (
            O => \N__4784\,
            I => \N__4781\
        );

    \I__589\ : Odrv12
    port map (
            O => \N__4781\,
            I => \un2_D_LL_AMIGA_0\
        );

    \I__588\ : InMux
    port map (
            O => \N__4778\,
            I => \N__4775\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4775\,
            I => \N__4772\
        );

    \I__586\ : Odrv12
    port map (
            O => \N__4772\,
            I => \D_LM_AMIGA_in_1\
        );

    \I__585\ : IoInMux
    port map (
            O => \N__4769\,
            I => \N__4766\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__583\ : Span4Mux_s3_h
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__582\ : Span4Mux_h
    port map (
            O => \N__4760\,
            I => \N__4757\
        );

    \I__581\ : Sp12to4
    port map (
            O => \N__4757\,
            I => \N__4754\
        );

    \I__580\ : Span12Mux_v
    port map (
            O => \N__4754\,
            I => \N__4751\
        );

    \I__579\ : Span12Mux_h
    port map (
            O => \N__4751\,
            I => \N__4748\
        );

    \I__578\ : Odrv12
    port map (
            O => \N__4748\,
            I => \un2_D_LM_AMIGA_1\
        );

    \I__577\ : InMux
    port map (
            O => \N__4745\,
            I => \N__4742\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__4742\,
            I => \N__4739\
        );

    \I__575\ : Span12Mux_h
    port map (
            O => \N__4739\,
            I => \N__4736\
        );

    \I__574\ : Span12Mux_h
    port map (
            O => \N__4736\,
            I => \N__4733\
        );

    \I__573\ : Odrv12
    port map (
            O => \N__4733\,
            I => \D_UM_040_in_2\
        );

    \I__572\ : IoInMux
    port map (
            O => \N__4730\,
            I => \N__4726\
        );

    \I__571\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4723\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4726\,
            I => \N__4720\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__4723\,
            I => \N__4717\
        );

    \I__568\ : IoSpan4Mux
    port map (
            O => \N__4720\,
            I => \N__4714\
        );

    \I__567\ : Span4Mux_v
    port map (
            O => \N__4717\,
            I => \N__4711\
        );

    \I__566\ : Span4Mux_s2_h
    port map (
            O => \N__4714\,
            I => \N__4708\
        );

    \I__565\ : Sp12to4
    port map (
            O => \N__4711\,
            I => \N__4705\
        );

    \I__564\ : Sp12to4
    port map (
            O => \N__4708\,
            I => \N__4702\
        );

    \I__563\ : Span12Mux_v
    port map (
            O => \N__4705\,
            I => \N__4699\
        );

    \I__562\ : Span12Mux_h
    port map (
            O => \N__4702\,
            I => \N__4696\
        );

    \I__561\ : Span12Mux_h
    port map (
            O => \N__4699\,
            I => \N__4693\
        );

    \I__560\ : Span12Mux_h
    port map (
            O => \N__4696\,
            I => \N__4690\
        );

    \I__559\ : Odrv12
    port map (
            O => \N__4693\,
            I => \D_LL_040_in_2\
        );

    \I__558\ : Odrv12
    port map (
            O => \N__4690\,
            I => \D_LL_040_in_2\
        );

    \I__557\ : IoInMux
    port map (
            O => \N__4685\,
            I => \N__4682\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4682\,
            I => \N__4679\
        );

    \I__555\ : Span4Mux_s3_h
    port map (
            O => \N__4679\,
            I => \N__4676\
        );

    \I__554\ : Span4Mux_h
    port map (
            O => \N__4676\,
            I => \N__4673\
        );

    \I__553\ : Span4Mux_v
    port map (
            O => \N__4673\,
            I => \N__4670\
        );

    \I__552\ : Odrv4
    port map (
            O => \N__4670\,
            I => \un1_D_UM_040_2\
        );

    \I__551\ : IoInMux
    port map (
            O => \N__4667\,
            I => \N__4664\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4664\,
            I => \N__4661\
        );

    \I__549\ : Span4Mux_s3_v
    port map (
            O => \N__4661\,
            I => \N__4658\
        );

    \I__548\ : Span4Mux_h
    port map (
            O => \N__4658\,
            I => \N__4655\
        );

    \I__547\ : Odrv4
    port map (
            O => \N__4655\,
            I => \N_216_i\
        );

    \I__546\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__4649\,
            I => \N__4646\
        );

    \I__544\ : Odrv12
    port map (
            O => \N__4646\,
            I => \WRITE_CYCLE_ACTIVE_rep5_i_ess\
        );

    \I__543\ : IoInMux
    port map (
            O => \N__4643\,
            I => \N__4640\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4640\,
            I => \N__4637\
        );

    \I__541\ : Span4Mux_s3_h
    port map (
            O => \N__4637\,
            I => \N__4634\
        );

    \I__540\ : Span4Mux_v
    port map (
            O => \N__4634\,
            I => \N__4631\
        );

    \I__539\ : Odrv4
    port map (
            O => \N__4631\,
            I => \N_218_i\
        );

    \I__538\ : InMux
    port map (
            O => \N__4628\,
            I => \N__4625\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__536\ : Span4Mux_h
    port map (
            O => \N__4622\,
            I => \N__4619\
        );

    \I__535\ : Span4Mux_v
    port map (
            O => \N__4619\,
            I => \N__4616\
        );

    \I__534\ : Odrv4
    port map (
            O => \N__4616\,
            I => \A_040_c_0\
        );

    \I__533\ : IoInMux
    port map (
            O => \N__4613\,
            I => \N__4610\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__531\ : Span4Mux_s2_v
    port map (
            O => \N__4607\,
            I => \N__4604\
        );

    \I__530\ : Span4Mux_v
    port map (
            O => \N__4604\,
            I => \N__4601\
        );

    \I__529\ : Odrv4
    port map (
            O => \N__4601\,
            I => \A_AMIGA_c_0\
        );

    \I__528\ : IoInMux
    port map (
            O => \N__4598\,
            I => \N__4595\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4595\,
            I => \N__4592\
        );

    \I__526\ : Odrv12
    port map (
            O => \N__4592\,
            I => \U111_CYCLE_SM_A_AMIGA_0_i_1\
        );

    \I__525\ : InMux
    port map (
            O => \N__4589\,
            I => \N__4586\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4586\,
            I => \WRITE_CYCLE_ACTIVE_rep28_i_ess\
        );

    \I__523\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4580\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4580\,
            I => \N__4577\
        );

    \I__521\ : Span4Mux_v
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__520\ : Odrv4
    port map (
            O => \N__4574\,
            I => \WRITE_CYCLE_ACTIVE_rep27_i_ess\
        );

    \I__519\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4568\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4568\,
            I => \WRITE_CYCLE_ACTIVE_rep19_i_ess\
        );

    \I__517\ : IoInMux
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4562\,
            I => \N__4559\
        );

    \I__515\ : Odrv12
    port map (
            O => \N__4559\,
            I => \N_231_i\
        );

    \I__514\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4553\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4553\,
            I => \WRITE_CYCLE_ACTIVE_rep18_i_ess\
        );

    \I__512\ : IoInMux
    port map (
            O => \N__4550\,
            I => \N__4547\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4547\,
            I => \N__4544\
        );

    \I__510\ : Odrv12
    port map (
            O => \N__4544\,
            I => \N_232_i\
        );

    \I__509\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4538\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4538\,
            I => \WRITE_CYCLE_ACTIVE_rep8_i_ess\
        );

    \I__507\ : InMux
    port map (
            O => \N__4535\,
            I => \N__4532\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4532\,
            I => \WRITE_CYCLE_ACTIVE_rep20_i_ess\
        );

    \I__505\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4526\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__4526\,
            I => \WRITE_CYCLE_ACTIVE_rep11_i_ess\
        );

    \I__503\ : InMux
    port map (
            O => \N__4523\,
            I => \N__4520\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4520\,
            I => \WRITE_CYCLE_ACTIVE_rep22_i_ess\
        );

    \I__501\ : InMux
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4514\,
            I => \WRITE_CYCLE_ACTIVE_rep14_i_ess\
        );

    \I__499\ : InMux
    port map (
            O => \N__4511\,
            I => \N__4508\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4508\,
            I => \WRITE_CYCLE_ACTIVE_rep1_i_ess\
        );

    \I__497\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4502\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__4502\,
            I => \WRITE_CYCLE_ACTIVE_rep12_i_ess\
        );

    \I__495\ : IoInMux
    port map (
            O => \N__4499\,
            I => \N__4496\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4496\,
            I => \N__4493\
        );

    \I__493\ : IoSpan4Mux
    port map (
            O => \N__4493\,
            I => \N__4490\
        );

    \I__492\ : Span4Mux_s2_h
    port map (
            O => \N__4490\,
            I => \N__4487\
        );

    \I__491\ : Odrv4
    port map (
            O => \N__4487\,
            I => \N_214_i\
        );

    \I__490\ : IoInMux
    port map (
            O => \N__4484\,
            I => \N__4481\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4481\,
            I => \N__4478\
        );

    \I__488\ : IoSpan4Mux
    port map (
            O => \N__4478\,
            I => \N__4475\
        );

    \I__487\ : Span4Mux_s3_h
    port map (
            O => \N__4475\,
            I => \N__4472\
        );

    \I__486\ : Odrv4
    port map (
            O => \N__4472\,
            I => \N_228_i\
        );

    \I__485\ : IoInMux
    port map (
            O => \N__4469\,
            I => \N__4466\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4466\,
            I => \N__4463\
        );

    \I__483\ : IoSpan4Mux
    port map (
            O => \N__4463\,
            I => \N__4460\
        );

    \I__482\ : Span4Mux_s2_h
    port map (
            O => \N__4460\,
            I => \N__4457\
        );

    \I__481\ : Odrv4
    port map (
            O => \N__4457\,
            I => \N_225_i\
        );

    \I__480\ : InMux
    port map (
            O => \N__4454\,
            I => \N__4451\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4451\,
            I => \WRITE_CYCLE_ACTIVE_rep15_i_ess\
        );

    \I__478\ : IoInMux
    port map (
            O => \N__4448\,
            I => \N__4445\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4445\,
            I => \N__4442\
        );

    \I__476\ : IoSpan4Mux
    port map (
            O => \N__4442\,
            I => \N__4439\
        );

    \I__475\ : Span4Mux_s1_h
    port map (
            O => \N__4439\,
            I => \N__4436\
        );

    \I__474\ : Span4Mux_h
    port map (
            O => \N__4436\,
            I => \N__4433\
        );

    \I__473\ : Odrv4
    port map (
            O => \N__4433\,
            I => \N_241_i\
        );

    \I__472\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4427\,
            I => \WRITE_CYCLE_ACTIVE_rep25_i_ess\
        );

    \I__470\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4421\,
            I => \WRITE_CYCLE_ACTIVE_rep30_i_ess\
        );

    \I__468\ : InMux
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4415\,
            I => \WRITE_CYCLE_ACTIVE_i_ess\
        );

    \I__466\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4409\,
            I => \WRITE_CYCLE_ACTIVE_rep16_i_ess\
        );

    \I__464\ : IoInMux
    port map (
            O => \N__4406\,
            I => \N__4403\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4403\,
            I => \N__4400\
        );

    \I__462\ : Span12Mux_s4_h
    port map (
            O => \N__4400\,
            I => \N__4397\
        );

    \I__461\ : Odrv12
    port map (
            O => \N__4397\,
            I => \N_223_i\
        );

    \I__460\ : IoInMux
    port map (
            O => \N__4394\,
            I => \N__4391\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__4391\,
            I => \N__4388\
        );

    \I__458\ : IoSpan4Mux
    port map (
            O => \N__4388\,
            I => \N__4385\
        );

    \I__457\ : Span4Mux_s3_h
    port map (
            O => \N__4385\,
            I => \N__4382\
        );

    \I__456\ : Odrv4
    port map (
            O => \N__4382\,
            I => \N_233_i\
        );

    \I__455\ : InMux
    port map (
            O => \N__4379\,
            I => \N__4376\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__4376\,
            I => \WRITE_CYCLE_ACTIVE_rep10_i_ess\
        );

    \I__453\ : IoInMux
    port map (
            O => \N__4373\,
            I => \N__4370\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4370\,
            I => \N__4367\
        );

    \I__451\ : Span12Mux_s4_h
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__450\ : Odrv12
    port map (
            O => \N__4364\,
            I => \N_234_i\
        );

    \I__449\ : InMux
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4358\,
            I => \WRITE_CYCLE_ACTIVE_rep9_i_ess\
        );

    \I__447\ : IoInMux
    port map (
            O => \N__4355\,
            I => \N__4352\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__4352\,
            I => \N__4349\
        );

    \I__445\ : IoSpan4Mux
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__444\ : Span4Mux_s3_h
    port map (
            O => \N__4346\,
            I => \N__4343\
        );

    \I__443\ : Odrv4
    port map (
            O => \N__4343\,
            I => \N_222_i\
        );

    \I__442\ : IoInMux
    port map (
            O => \N__4340\,
            I => \N__4337\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__4337\,
            I => \N__4334\
        );

    \I__440\ : IoSpan4Mux
    port map (
            O => \N__4334\,
            I => \N__4331\
        );

    \I__439\ : Span4Mux_s3_h
    port map (
            O => \N__4331\,
            I => \N__4328\
        );

    \I__438\ : Odrv4
    port map (
            O => \N__4328\,
            I => \N_236_i\
        );

    \I__437\ : IoInMux
    port map (
            O => \N__4325\,
            I => \N__4322\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__435\ : Span4Mux_s0_h
    port map (
            O => \N__4319\,
            I => \N__4316\
        );

    \I__434\ : Span4Mux_h
    port map (
            O => \N__4316\,
            I => \N__4313\
        );

    \I__433\ : Odrv4
    port map (
            O => \N__4313\,
            I => \N_235_i\
        );

    \I__432\ : IoInMux
    port map (
            O => \N__4310\,
            I => \N__4307\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__4307\,
            I => \N__4304\
        );

    \I__430\ : Span4Mux_s3_h
    port map (
            O => \N__4304\,
            I => \N__4301\
        );

    \I__429\ : Span4Mux_v
    port map (
            O => \N__4301\,
            I => \N__4298\
        );

    \I__428\ : Odrv4
    port map (
            O => \N__4298\,
            I => \N_224_i\
        );

    \I__427\ : IoInMux
    port map (
            O => \N__4295\,
            I => \N__4292\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__425\ : Span12Mux_s4_h
    port map (
            O => \N__4289\,
            I => \N__4286\
        );

    \I__424\ : Odrv12
    port map (
            O => \N__4286\,
            I => \N_227_i\
        );

    \I__423\ : IoInMux
    port map (
            O => \N__4283\,
            I => \N__4280\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4280\,
            I => \N__4277\
        );

    \I__421\ : Span4Mux_s0_h
    port map (
            O => \N__4277\,
            I => \N__4274\
        );

    \I__420\ : Span4Mux_h
    port map (
            O => \N__4274\,
            I => \N__4271\
        );

    \I__419\ : Odrv4
    port map (
            O => \N__4271\,
            I => \N_243_i\
        );

    \I__418\ : IoInMux
    port map (
            O => \N__4268\,
            I => \N__4265\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__4265\,
            I => \N__4262\
        );

    \I__416\ : Span12Mux_s4_h
    port map (
            O => \N__4262\,
            I => \N__4259\
        );

    \I__415\ : Odrv12
    port map (
            O => \N__4259\,
            I => \N_229_i\
        );

    \I__414\ : IoInMux
    port map (
            O => \N__4256\,
            I => \N__4253\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__412\ : Span4Mux_s0_h
    port map (
            O => \N__4250\,
            I => \N__4247\
        );

    \I__411\ : Span4Mux_h
    port map (
            O => \N__4247\,
            I => \N__4244\
        );

    \I__410\ : Odrv4
    port map (
            O => \N__4244\,
            I => \N_244_i\
        );

    \I__409\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4238\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__4238\,
            I => \N__4235\
        );

    \I__407\ : Odrv4
    port map (
            O => \N__4235\,
            I => \WRITE_CYCLE_ACTIVE_rep29_i_ess\
        );

    \I__406\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4229\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__4229\,
            I => \WRITE_CYCLE_ACTIVE_rep17_i_ess\
        );

    \I__404\ : IoInMux
    port map (
            O => \N__4226\,
            I => \N__4223\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__4223\,
            I => \N__4220\
        );

    \I__402\ : IoSpan4Mux
    port map (
            O => \N__4220\,
            I => \N__4217\
        );

    \I__401\ : Span4Mux_s3_h
    port map (
            O => \N__4217\,
            I => \N__4214\
        );

    \I__400\ : Odrv4
    port map (
            O => \N__4214\,
            I => \N_230_i\
        );

    \I__399\ : IoInMux
    port map (
            O => \N__4211\,
            I => \N__4208\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__4208\,
            I => \N__4205\
        );

    \I__397\ : Odrv12
    port map (
            O => \N__4205\,
            I => \RESETn_c_i\
        );

    \I__396\ : IoInMux
    port map (
            O => \N__4202\,
            I => \N__4199\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4199\,
            I => \N__4196\
        );

    \I__394\ : IoSpan4Mux
    port map (
            O => \N__4196\,
            I => \N__4193\
        );

    \I__393\ : Span4Mux_s1_h
    port map (
            O => \N__4193\,
            I => \N__4190\
        );

    \I__392\ : Odrv4
    port map (
            O => \N__4190\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_0\
        );

    \I__391\ : IoInMux
    port map (
            O => \N__4187\,
            I => \N__4184\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__4184\,
            I => \N__4181\
        );

    \I__389\ : Odrv12
    port map (
            O => \N__4181\,
            I => \N_221_i\
        );

    \I__388\ : IoInMux
    port map (
            O => \N__4178\,
            I => \N__4175\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__4175\,
            I => \N__4172\
        );

    \I__386\ : Span4Mux_s0_v
    port map (
            O => \N__4172\,
            I => \N__4169\
        );

    \I__385\ : Sp12to4
    port map (
            O => \N__4169\,
            I => \N__4166\
        );

    \I__384\ : Span12Mux_h
    port map (
            O => \N__4166\,
            I => \N__4163\
        );

    \I__383\ : Span12Mux_v
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__382\ : Span12Mux_v
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__381\ : Odrv12
    port map (
            O => \N__4157\,
            I => \TAn_in\
        );

    \I__380\ : IoInMux
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__4151\,
            I => \N__4148\
        );

    \I__378\ : IoSpan4Mux
    port map (
            O => \N__4148\,
            I => \N__4145\
        );

    \I__377\ : Span4Mux_s3_h
    port map (
            O => \N__4145\,
            I => \N__4142\
        );

    \I__376\ : Odrv4
    port map (
            O => \N__4142\,
            I => \N_240_i\
        );

    \I__375\ : IoInMux
    port map (
            O => \N__4139\,
            I => \N__4136\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__4136\,
            I => \N__4133\
        );

    \I__373\ : Span4Mux_s3_h
    port map (
            O => \N__4133\,
            I => \N__4130\
        );

    \I__372\ : Span4Mux_v
    port map (
            O => \N__4130\,
            I => \N__4127\
        );

    \I__371\ : Odrv4
    port map (
            O => \N__4127\,
            I => \N_237_i\
        );

    \I__370\ : IoInMux
    port map (
            O => \N__4124\,
            I => \N__4121\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__4121\,
            I => \N__4118\
        );

    \I__368\ : IoSpan4Mux
    port map (
            O => \N__4118\,
            I => \N__4115\
        );

    \I__367\ : Span4Mux_s2_h
    port map (
            O => \N__4115\,
            I => \N__4112\
        );

    \I__366\ : Odrv4
    port map (
            O => \N__4112\,
            I => \N_239_i\
        );

    \I__365\ : InMux
    port map (
            O => \N__4109\,
            I => \N__4106\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__4106\,
            I => \WRITE_CYCLE_ACTIVE_rep26_i_ess\
        );

    \I__363\ : IoInMux
    port map (
            O => \N__4103\,
            I => \N__4100\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__361\ : Span4Mux_s3_h
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__360\ : Span4Mux_v
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__359\ : Odrv4
    port map (
            O => \N__4091\,
            I => \N_238_i\
        );

    \I__358\ : InMux
    port map (
            O => \N__4088\,
            I => \N__4085\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__356\ : Odrv4
    port map (
            O => \N__4082\,
            I => \WRITE_CYCLE_ACTIVE_rep24_i_ess\
        );

    \I__355\ : IoInMux
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__353\ : Span4Mux_s0_h
    port map (
            O => \N__4073\,
            I => \N__4070\
        );

    \I__352\ : Span4Mux_h
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__351\ : Odrv4
    port map (
            O => \N__4067\,
            I => \N_242_i\
        );

    \I__350\ : IoInMux
    port map (
            O => \N__4064\,
            I => \N__4061\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__348\ : IoSpan4Mux
    port map (
            O => \N__4058\,
            I => \N__4055\
        );

    \I__347\ : Span4Mux_s3_h
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__346\ : Sp12to4
    port map (
            O => \N__4052\,
            I => \N__4049\
        );

    \I__345\ : Span12Mux_s8_h
    port map (
            O => \N__4049\,
            I => \N__4046\
        );

    \I__344\ : Span12Mux_v
    port map (
            O => \N__4046\,
            I => \N__4043\
        );

    \I__343\ : Span12Mux_v
    port map (
            O => \N__4043\,
            I => \N__4040\
        );

    \I__342\ : Span12Mux_h
    port map (
            O => \N__4040\,
            I => \N__4037\
        );

    \I__341\ : Odrv12
    port map (
            O => \N__4037\,
            I => \TCIn_c\
        );

    \INVU111_CYCLE_SM.TSnC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TSnC_net\,
            I => \N__12817\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4211\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4202\,
            GLOBALBUFFEROUTPUT => \U111_CYCLE_SM.CYCLE_STATE_0_g_0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_3_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4583\,
            lcout => \N_240_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_0_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4088\,
            lcout => \N_237_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_2_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4109\,
            lcout => \N_239_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__10382\,
            in1 => \N__11764\,
            in2 => \N__12216\,
            in3 => \N__10703\,
            lcout => \WRITE_CYCLE_ACTIVE_rep26_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12843\,
            ce => \N__12626\,
            sr => \N__12473\
        );

    \D_LL_AMIGA_iobuf_RNO_1_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4430\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_238_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__11077\,
            in1 => \N__12167\,
            in2 => \N__11630\,
            in3 => \N__10586\,
            lcout => \WRITE_CYCLE_ACTIVE_rep24_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12837\,
            ce => \N__12620\,
            sr => \N__12469\
        );

    \D_LL_AMIGA_iobuf_RNO_5_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4241\,
            lcout => \N_242_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4424\,
            lcout => \N_243_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_0_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4412\,
            lcout => \N_229_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_7_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4418\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_244_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__10573\,
            in1 => \N__12116\,
            in2 => \N__11759\,
            in3 => \N__11023\,
            lcout => \WRITE_CYCLE_ACTIVE_rep17_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12831\,
            ce => \N__12614\,
            sr => \N__12462\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__11024\,
            in1 => \N__12117\,
            in2 => \N__10585\,
            in3 => \N__11748\,
            lcout => \WRITE_CYCLE_ACTIVE_rep29_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12831\,
            ce => \N__12614\,
            sr => \N__12462\
        );

    \D_LM_AMIGA_iobuf_RNO_1_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4232\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_230_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7241\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__12515\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6770\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_0_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4541\,
            lcout => \N_221_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_2_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4379\,
            lcout => \N_223_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_4_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4535\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_233_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__11109\,
            in1 => \N__12022\,
            in2 => \N__11716\,
            in3 => \N__10535\,
            lcout => \WRITE_CYCLE_ACTIVE_rep10_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12820\,
            ce => \N__12615\,
            sr => \N__12466\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__12023\,
            in1 => \N__11688\,
            in2 => \N__10572\,
            in3 => \N__11113\,
            lcout => \WRITE_CYCLE_ACTIVE_rep9_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12820\,
            ce => \N__12615\,
            sr => \N__12466\
        );

    \D_LM_AMIGA_iobuf_RNO_5_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4874\,
            lcout => \N_234_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_1_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4361\,
            lcout => \N_222_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_7_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4865\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_236_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_6_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4523\,
            lcout => \N_235_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_3_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4529\,
            lcout => \N_224_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_6_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4517\,
            lcout => \N_227_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_1_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4511\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_214_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_7_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4454\,
            lcout => \N_228_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_4_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4505\,
            lcout => \N_225_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__10571\,
            in1 => \N__12166\,
            in2 => \N__11703\,
            in3 => \N__11168\,
            lcout => \WRITE_CYCLE_ACTIVE_rep15_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12798\,
            ce => \N__12630\,
            sr => \N__12487\
        );

    \D_LL_AMIGA_iobuf_RNO_4_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4589\,
            lcout => \N_241_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__10883\,
            in1 => \N__12243\,
            in2 => \N__11765\,
            in3 => \N__10584\,
            lcout => \WRITE_CYCLE_ACTIVE_rep25_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12838\,
            ce => \N__12627\,
            sr => \N__12474\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__10884\,
            in1 => \N__12089\,
            in2 => \N__11760\,
            in3 => \N__10582\,
            lcout => \WRITE_CYCLE_ACTIVE_rep30_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12834\,
            ce => \N__12621\,
            sr => \N__12470\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__12206\,
            in1 => \N__11744\,
            in2 => \N__10992\,
            in3 => \N__10581\,
            lcout => \WRITE_CYCLE_ACTIVE_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12832\,
            ce => \N__12619\,
            sr => \N__12467\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__10993\,
            in1 => \N__12205\,
            in2 => \N__11758\,
            in3 => \N__10554\,
            lcout => \WRITE_CYCLE_ACTIVE_rep16_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12827\,
            ce => \N__12617\,
            sr => \N__12463\
        );

    \D_LM_AMIGA_iobuf_RNO_3_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4571\,
            lcout => \N_232_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__11079\,
            in1 => \N__12204\,
            in2 => \N__11740\,
            in3 => \N__10504\,
            lcout => \WRITE_CYCLE_ACTIVE_rep8_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12822\,
            ce => \N__12613\,
            sr => \N__12464\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__12202\,
            in1 => \N__10503\,
            in2 => \N__11137\,
            in3 => \N__11588\,
            lcout => \WRITE_CYCLE_ACTIVE_rep20_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12821\,
            ce => \N__12616\,
            sr => \N__12468\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__12227\,
            in1 => \N__10485\,
            in2 => \N__11167\,
            in3 => \N__11684\,
            lcout => \WRITE_CYCLE_ACTIVE_rep11_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12815\,
            ce => \N__12622\,
            sr => \N__12475\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11632\,
            in1 => \N__12230\,
            in2 => \N__10549\,
            in3 => \N__11150\,
            lcout => \WRITE_CYCLE_ACTIVE_rep5_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12810\,
            ce => \N__12624\,
            sr => \N__12477\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11631\,
            in1 => \N__12229\,
            in2 => \N__10548\,
            in3 => \N__11149\,
            lcout => \WRITE_CYCLE_ACTIVE_rep22_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12810\,
            ce => \N__12624\,
            sr => \N__12477\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__10493\,
            in1 => \N__12252\,
            in2 => \N__11166\,
            in3 => \N__11649\,
            lcout => \WRITE_CYCLE_ACTIVE_rep14_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12805\,
            ce => \N__12628\,
            sr => \N__12482\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11650\,
            in1 => \N__10494\,
            in2 => \N__12260\,
            in3 => \N__11142\,
            lcout => \WRITE_CYCLE_ACTIVE_rep1_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12805\,
            ce => \N__12628\,
            sr => \N__12482\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__11144\,
            in1 => \N__12257\,
            in2 => \N__11705\,
            in3 => \N__10498\,
            lcout => \WRITE_CYCLE_ACTIVE_rep12_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12799\,
            ce => \N__12631\,
            sr => \N__12488\
        );

    \D_UU_AMIGA_iobuf_RNO_3_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4829\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_216_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_5_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4652\,
            lcout => \N_218_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__4628\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6025\,
            lcout => \A_AMIGA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__6026\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4891\,
            lcout => \U111_CYCLE_SM_A_AMIGA_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_3_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__10381\,
            in1 => \N__12244\,
            in2 => \N__11654\,
            in3 => \N__10693\,
            lcout => \WRITE_CYCLE_ACTIVE_rep28_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12839\,
            ce => \N__12634\,
            sr => \N__12484\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_3_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__12242\,
            in1 => \N__11589\,
            in2 => \N__11076\,
            in3 => \N__10583\,
            lcout => \WRITE_CYCLE_ACTIVE_rep27_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12836\,
            ce => \N__12632\,
            sr => \N__12478\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__10569\,
            in1 => \N__12203\,
            in2 => \N__11584\,
            in3 => \N__10994\,
            lcout => \WRITE_CYCLE_ACTIVE_rep19_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12823\,
            ce => \N__12612\,
            sr => \N__12465\
        );

    \D_LM_AMIGA_iobuf_RNO_2_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4556\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_231_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__10502\,
            in1 => \N__12171\,
            in2 => \N__11587\,
            in3 => \N__11078\,
            lcout => \WRITE_CYCLE_ACTIVE_rep18_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12819\,
            ce => \N__12618\,
            sr => \N__12471\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11506\,
            in1 => \N__12217\,
            in2 => \N__10372\,
            in3 => \N__11083\,
            lcout => \WRITE_CYCLE_ACTIVE_rep21_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12816\,
            ce => \N__12623\,
            sr => \N__12476\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__12226\,
            in1 => \N__11505\,
            in2 => \N__10568\,
            in3 => \N__11138\,
            lcout => \WRITE_CYCLE_ACTIVE_rep23_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12811\,
            ce => \N__12625\,
            sr => \N__12479\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__10486\,
            in1 => \N__12228\,
            in2 => \N__11453\,
            in3 => \N__11148\,
            lcout => \WRITE_CYCLE_ACTIVE_rep7_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12806\,
            ce => \N__12629\,
            sr => \N__12483\
        );

    \D_UU_AMIGA_iobuf_RNO_7_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4853\,
            lcout => \N_220_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11601\,
            in1 => \N__12256\,
            in2 => \N__10550\,
            in3 => \N__11143\,
            lcout => \WRITE_CYCLE_ACTIVE_rep3_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12793\,
            ce => \N__12633\,
            sr => \N__12490\
        );

    \D_UU_AMIGA_iobuf_RNO_6_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4943\,
            lcout => \N_219_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8827\,
            in1 => \N__4808\,
            in2 => \_gnd_net_\,
            in3 => \N__8975\,
            lcout => \un2_D_LL_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8735\,
            in1 => \N__6530\,
            in2 => \_gnd_net_\,
            in3 => \N__4778\,
            lcout => \un2_D_LM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__4745\,
            in1 => \N__8741\,
            in2 => \_gnd_net_\,
            in3 => \N__4729\,
            lcout => \un1_D_UM_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5081\,
            in1 => \N__5053\,
            in2 => \_gnd_net_\,
            in3 => \N__8792\,
            lcout => \un1_D_UM_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8791\,
            in1 => \N__7698\,
            in2 => \_gnd_net_\,
            in3 => \N__5009\,
            lcout => \un2_D_LM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__10461\,
            in1 => \N__12251\,
            in2 => \N__11182\,
            in3 => \N__11560\,
            lcout => \WRITE_CYCLE_ACTIVE_rep0_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12790\,
            ce => \N__12635\,
            sr => \N__12491\
        );

    \D_UU_AMIGA_iobuf_RNO_0_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4982\,
            lcout => \N_213_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_5_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5303\,
            lcout => \N_226_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__12073\,
            in1 => \N__11558\,
            in2 => \N__11183\,
            in3 => \N__10528\,
            lcout => \WRITE_CYCLE_ACTIVE_rep4_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12784\,
            ce => \N__12638\,
            sr => \N__12493\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11559\,
            in1 => \N__12074\,
            in2 => \N__10570\,
            in3 => \N__11181\,
            lcout => \WRITE_CYCLE_ACTIVE_rep6_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12784\,
            ce => \N__12638\,
            sr => \N__12493\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6963\,
            in1 => \N__4934\,
            in2 => \_gnd_net_\,
            in3 => \N__8828\,
            lcout => \un2_D_LL_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6088\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4901\,
            lcout => \U111_CYCLE_SM.FLIP_WORD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__11161\,
            in1 => \N__12259\,
            in2 => \N__11655\,
            in3 => \N__10527\,
            lcout => \WRITE_CYCLE_ACTIVE_rep13_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12783\,
            ce => \N__12637\,
            sr => \N__12492\
        );

    \D_UU_AMIGA_iobuf_RNO_4_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5297\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_217_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5276\,
            in1 => \N__8465\,
            in2 => \_gnd_net_\,
            in3 => \N__8823\,
            lcout => \un2_D_LL_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5239\,
            in1 => \N__5195\,
            in2 => \_gnd_net_\,
            in3 => \N__8710\,
            lcout => \un1_D_UM_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8645\,
            in1 => \N__8006\,
            in2 => \_gnd_net_\,
            in3 => \N__5159\,
            lcout => \un2_D_LM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11522\,
            in1 => \N__12258\,
            in2 => \N__10454\,
            in3 => \N__11157\,
            lcout => \WRITE_CYCLE_ACTIVE_rep2_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12782\,
            ce => \N__12639\,
            sr => \N__12494\
        );

    \BUFENn_obuf_RNO_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11174\,
            lcout => \LBENn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_2_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5105\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_215_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9392\,
            in1 => \N__5687\,
            in2 => \_gnd_net_\,
            in3 => \N__8768\,
            lcout => \un2_D_LL_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8769\,
            in1 => \N__6887\,
            in2 => \_gnd_net_\,
            in3 => \N__5648\,
            lcout => \un2_D_LM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TSn_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7240\,
            in2 => \_gnd_net_\,
            in3 => \N__5593\,
            lcout => \TSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TSnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011111111"
        )
    port map (
            in0 => \N__6722\,
            in1 => \N__5594\,
            in2 => \N__5717\,
            in3 => \N__5729\,
            lcout => \U111_CYCLE_SM.TS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12812\,
            ce => 'H',
            sr => \N__12472\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5582\,
            in1 => \N__5557\,
            in2 => \_gnd_net_\,
            in3 => \N__8745\,
            lcout => \un1_D_UM_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8746\,
            in1 => \N__7920\,
            in2 => \_gnd_net_\,
            in3 => \N__5501\,
            lcout => \un2_D_LM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5455\,
            in1 => \N__5429\,
            in2 => \_gnd_net_\,
            in3 => \N__8747\,
            lcout => \un1_D_UU_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8797\,
            in1 => \N__5395\,
            in2 => \_gnd_net_\,
            in3 => \N__5345\,
            lcout => \un1_D_UM_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8798\,
            in1 => \N__5840\,
            in2 => \_gnd_net_\,
            in3 => \N__5815\,
            lcout => \un1_D_UU_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8734\,
            in1 => \N__5762\,
            in2 => \_gnd_net_\,
            in3 => \N__7540\,
            lcout => \un2_D_LL_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LATCH_EN_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__6689\,
            in1 => \N__5728\,
            in2 => \N__9025\,
            in3 => \N__6766\,
            lcout => \U111_CYCLE_SM.LATCH_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12813\,
            ce => 'H',
            sr => \N__12480\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIDUAQ_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__12094\,
            in1 => \N__11704\,
            in2 => \N__11133\,
            in3 => \N__6760\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\,
            ltout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIC4111_3_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__6181\,
            in1 => \_gnd_net_\,
            in2 => \N__5732\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.un1_CYCLE_STATE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_4_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7242\,
            in2 => \_gnd_net_\,
            in3 => \N__6182\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6180\,
            in1 => \N__6598\,
            in2 => \N__7186\,
            in3 => \N__6228\,
            lcout => \U111_CYCLE_SM.TS_EN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__6639\,
            in1 => \N__6154\,
            in2 => \N__6133\,
            in3 => \N__6599\,
            lcout => \U111_CYCLE_SM.BURSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12800\,
            ce => 'H',
            sr => \N__12481\
        );

    \U111_CYCLE_SM.BURST_COUNT_1_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__6671\,
            in1 => \N__6638\,
            in2 => \N__6302\,
            in3 => \N__6617\,
            lcout => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12800\,
            ce => 'H',
            sr => \N__12481\
        );

    \U111_CYCLE_SM.LW_TRANS_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__6640\,
            in1 => \N__6155\,
            in2 => \N__6134\,
            in3 => \N__6046\,
            lcout => \U111_CYCLE_SM.LW_TRANSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12800\,
            ce => 'H',
            sr => \N__12481\
        );

    \U111_CYCLE_SM.TA_DIS_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__6184\,
            in1 => \N__6237\,
            in2 => \N__7123\,
            in3 => \N__6032\,
            lcout => \U111_CYCLE_SM.TA_DISZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12800\,
            ce => 'H',
            sr => \N__12481\
        );

    \U111_CYCLE_SM.FLIP_WORD_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__8596\,
            in1 => \N__6183\,
            in2 => \N__6110\,
            in3 => \N__6238\,
            lcout => \U111_CYCLE_SM.FLIP_WORDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12800\,
            ce => 'H',
            sr => \N__12481\
        );

    \U111_CYCLE_SM.PORT_MISMATCH_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__6047\,
            in1 => \N__6239\,
            in2 => \N__6212\,
            in3 => \N__6084\,
            lcout => \U111_CYCLE_SM.PORT_MISMATCHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12800\,
            ce => 'H',
            sr => \N__12481\
        );

    \U111_CYCLE_SM.TA_DIS_RNO_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6092\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6045\,
            lcout => \U111_CYCLE_SM.PORT_MISMATCH_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__6188\,
            in1 => \N__6010\,
            in2 => \_gnd_net_\,
            in3 => \N__6553\,
            lcout => \U111_CYCLE_SM.A2_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12795\,
            ce => 'H',
            sr => \N__12485\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7029\,
            in1 => \N__5999\,
            in2 => \_gnd_net_\,
            in3 => \N__8666\,
            lcout => \un2_D_LM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5959\,
            in1 => \N__5915\,
            in2 => \_gnd_net_\,
            in3 => \N__8796\,
            lcout => \un1_D_UU_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8807\,
            in1 => \N__9332\,
            in2 => \_gnd_net_\,
            in3 => \N__5882\,
            lcout => \un2_D_LL_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6522\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12808\,
            ce => \N__7868\,
            sr => \N__7796\
        );

    \U111_CYCLE_SM.CYCLE_STATE_1_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__6641\,
            in1 => \N__6557\,
            in2 => \N__7254\,
            in3 => \N__6597\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12801\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7166\,
            in2 => \_gnd_net_\,
            in3 => \N__6711\,
            lcout => \U111_CYCLE_SM.N_124_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__6712\,
            in1 => \N__6206\,
            in2 => \N__7414\,
            in3 => \N__6251\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_132_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_0_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111111111"
        )
    port map (
            in0 => \N__7329\,
            in1 => \N__6311\,
            in2 => \N__6305\,
            in3 => \N__6569\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12801\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__6298\,
            in1 => \N__6615\,
            in2 => \N__6287\,
            in3 => \N__6596\,
            lcout => \U111_CYCLE_SM.un7_CYCLE_STATE_0\,
            ltout => \U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010111"
        )
    port map (
            in0 => \N__7330\,
            in1 => \N__7405\,
            in2 => \N__6245\,
            in3 => \N__6207\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_2_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__6713\,
            in1 => \N__7255\,
            in2 => \N__6242\,
            in3 => \N__6236\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12801\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_3_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6663\,
            in1 => \N__7246\,
            in2 => \_gnd_net_\,
            in3 => \N__6208\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12801\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_COUNT_0_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6637\,
            in1 => \N__6664\,
            in2 => \_gnd_net_\,
            in3 => \N__6616\,
            lcout => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12796\,
            ce => 'H',
            sr => \N__12486\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__7410\,
            in1 => \N__7150\,
            in2 => \_gnd_net_\,
            in3 => \N__6595\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_131_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001100"
        )
    port map (
            in0 => \N__6563\,
            in1 => \N__7267\,
            in2 => \N__6572\,
            in3 => \N__6765\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_4_0_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__11037\,
            in1 => \N__12013\,
            in2 => \_gnd_net_\,
            in3 => \N__11605\,
            lcout => \U111_CYCLE_SM.TS_EN6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__7409\,
            in1 => \N__7332\,
            in2 => \_gnd_net_\,
            in3 => \N__7154\,
            lcout => \U111_CYCLE_SM.N_144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6542\,
            in1 => \N__6523\,
            in2 => \_gnd_net_\,
            in3 => \N__9096\,
            lcout => \un1_D_UU_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6461\,
            in1 => \N__6446\,
            in2 => \_gnd_net_\,
            in3 => \N__8781\,
            lcout => \un1_D_UM_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6373\,
            in1 => \N__6344\,
            in2 => \_gnd_net_\,
            in3 => \N__8815\,
            lcout => \un1_D_UU_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LBENn_c_sbtinv_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10686\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \LBENn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8808\,
            in1 => \N__8318\,
            in2 => \_gnd_net_\,
            in3 => \N__6809\,
            lcout => \un2_D_LL_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_2_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7368\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7311\,
            lcout => \U111_CYCLE_SM.N_119_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__10567\,
            in1 => \N__12093\,
            in2 => \N__11585\,
            in3 => \N__10876\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12802\,
            ce => \N__12636\,
            sr => \N__12489\
        );

    \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__6710\,
            in1 => \N__6764\,
            in2 => \N__6734\,
            in3 => \N__7161\,
            lcout => \U111_CYCLE_SM.N_117_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__7386\,
            in1 => \N__7331\,
            in2 => \_gnd_net_\,
            in3 => \N__6709\,
            lcout => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa\,
            ltout => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3B1_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110101"
        )
    port map (
            in0 => \N__7253\,
            in1 => \_gnd_net_\,
            in2 => \N__6692\,
            in3 => \N__6685\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1\,
            ltout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNI9Q9V1_2_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6674\,
            in3 => \N__6662\,
            lcout => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7031\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12792\,
            ce => \N__7858\,
            sr => \N__7794\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6968\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12792\,
            ce => \N__7858\,
            sr => \N__7794\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6886\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12792\,
            ce => \N__7858\,
            sr => \N__7794\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7387\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7333\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_5_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__7268\,
            in1 => \N__7190\,
            in2 => \N__7169\,
            in3 => \N__7165\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11038\,
            in2 => \_gnd_net_\,
            in3 => \N__7127\,
            lcout => \TAn_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7085\,
            in1 => \N__7600\,
            in2 => \_gnd_net_\,
            in3 => \N__8721\,
            lcout => \un2_D_LM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9105\,
            in1 => \N__7043\,
            in2 => \_gnd_net_\,
            in3 => \N__7030\,
            lcout => \un1_D_UU_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6964\,
            in1 => \N__6926\,
            in2 => \_gnd_net_\,
            in3 => \N__9104\,
            lcout => \un1_D_UM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6896\,
            in1 => \N__6867\,
            in2 => \_gnd_net_\,
            in3 => \N__9107\,
            lcout => \un1_D_UU_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7457\,
            in1 => \N__8261\,
            in2 => \_gnd_net_\,
            in3 => \N__8756\,
            lcout => \un2_D_LL_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8967\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12794\,
            ce => \N__7865\,
            sr => \N__7797\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8311\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12791\,
            ce => \N__7867\,
            sr => \N__7795\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7928\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12791\,
            ce => \N__7867\,
            sr => \N__7795\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9384\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12791\,
            ce => \N__7867\,
            sr => \N__7795\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8005\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12787\,
            ce => \N__7866\,
            sr => \N__7798\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8464\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12787\,
            ce => \N__7866\,
            sr => \N__7798\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9321\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12787\,
            ce => \N__7866\,
            sr => \N__7798\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8375\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12787\,
            ce => \N__7866\,
            sr => \N__7798\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7541\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12787\,
            ce => \N__7866\,
            sr => \N__7798\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7599\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12787\,
            ce => \N__7866\,
            sr => \N__7798\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8256\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12787\,
            ce => \N__7866\,
            sr => \N__7798\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7700\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12785\,
            ce => \N__7857\,
            sr => \N__7805\
        );

    \GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7763\,
            lcout => \GB_BUFFER_CLK80_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9085\,
            in1 => \N__7709\,
            in2 => \_gnd_net_\,
            in3 => \N__7699\,
            lcout => \un1_D_UU_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8371\,
            in1 => \N__7640\,
            in2 => \_gnd_net_\,
            in3 => \N__9089\,
            lcout => \un1_D_UU_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__7610\,
            in1 => \_gnd_net_\,
            in2 => \N__9106\,
            in3 => \N__7601\,
            lcout => \un1_D_UU_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7536\,
            in1 => \N__7490\,
            in2 => \_gnd_net_\,
            in3 => \N__9090\,
            lcout => \un1_D_UM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9091\,
            in1 => \N__8474\,
            in2 => \_gnd_net_\,
            in3 => \N__8457\,
            lcout => \un1_D_UM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8393\,
            in1 => \N__8370\,
            in2 => \_gnd_net_\,
            in3 => \N__8757\,
            lcout => \un2_D_LM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9095\,
            in1 => \N__8327\,
            in2 => \_gnd_net_\,
            in3 => \N__8310\,
            lcout => \un1_D_UM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8260\,
            in1 => \N__8213\,
            in2 => \_gnd_net_\,
            in3 => \N__9108\,
            lcout => \un1_D_UM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8177\,
            in1 => \N__8159\,
            in2 => \_gnd_net_\,
            in3 => \N__8799\,
            lcout => \un1_D_UU_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8800\,
            in1 => \N__8096\,
            in2 => \_gnd_net_\,
            in3 => \N__8068\,
            lcout => \un1_D_UU_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7992\,
            in1 => \N__7961\,
            in2 => \_gnd_net_\,
            in3 => \N__9109\,
            lcout => \un1_D_UU_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7927\,
            in1 => \N__7898\,
            in2 => \_gnd_net_\,
            in3 => \N__9110\,
            lcout => \un1_D_UU_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9398\,
            in1 => \N__9391\,
            in2 => \_gnd_net_\,
            in3 => \N__9051\,
            lcout => \un1_D_UM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9338\,
            in1 => \N__9328\,
            in2 => \_gnd_net_\,
            in3 => \N__9052\,
            lcout => \un1_D_UM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9268\,
            in1 => \N__9224\,
            in2 => \_gnd_net_\,
            in3 => \N__8816\,
            lcout => \un1_D_UM_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8821\,
            in1 => \N__9182\,
            in2 => \_gnd_net_\,
            in3 => \N__9154\,
            lcout => \un1_D_UU_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9026\,
            in1 => \N__8984\,
            in2 => \_gnd_net_\,
            in3 => \N__8971\,
            lcout => \un1_D_UM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8915\,
            in1 => \N__8890\,
            in2 => \_gnd_net_\,
            in3 => \N__8817\,
            lcout => \un1_D_UM_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8822\,
            in1 => \N__8555\,
            in2 => \_gnd_net_\,
            in3 => \N__8527\,
            lcout => \un1_D_UU_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__12090\,
            in1 => \N__11126\,
            in2 => \N__10446\,
            in3 => \N__11507\,
            lcout => \READ_CYCLE_ACTIVE_rep4_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12786\,
            ce => \N__12643\,
            sr => \N__12500\
        );

    \D_UU_040_iobuf_RNO_4_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9509\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_185_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__12049\,
            in1 => \N__11513\,
            in2 => \N__10445\,
            in3 => \N__11162\,
            lcout => \READ_CYCLE_ACTIVE_rep2_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12789\,
            ce => \N__12645\,
            sr => \N__12501\
        );

    \D_UU_040_iobuf_RNO_2_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9488\,
            lcout => \N_183_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__11053\,
            in1 => \N__11937\,
            in2 => \N__10350\,
            in3 => \N__11342\,
            lcout => \READ_CYCLE_ACTIVE_rep0_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12809\,
            ce => \N__12646\,
            sr => \N__12502\
        );

    \D_UU_040_iobuf_RNO_0_LC_22_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9467\,
            lcout => \N_181_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_22_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11514\,
            in1 => \N__11938\,
            in2 => \N__10351\,
            in3 => \N__11054\,
            lcout => \READ_CYCLE_ACTIVE_rep7_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12797\,
            ce => \N__12649\,
            sr => \N__12507\
        );

    \D_UU_040_iobuf_RNO_7_LC_22_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9443\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_188_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_4_LC_23_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9404\,
            lcout => \N_209_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_23_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__12092\,
            in1 => \N__11710\,
            in2 => \N__10820\,
            in3 => \N__10444\,
            lcout => \READ_CYCLE_ACTIVE_rep28_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12842\,
            ce => \N__12653\,
            sr => \N__12505\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_23_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__12091\,
            in1 => \N__10450\,
            in2 => \N__11064\,
            in3 => \N__11709\,
            lcout => \READ_CYCLE_ACTIVE_rep26_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12840\,
            ce => \N__12650\,
            sr => \N__12503\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_23_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__10449\,
            in1 => \N__12043\,
            in2 => \N__11708\,
            in3 => \N__10961\,
            lcout => \READ_CYCLE_ACTIVE_rep18_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12835\,
            ce => \N__12647\,
            sr => \N__12498\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_23_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__12042\,
            in1 => \N__10448\,
            in2 => \N__11065\,
            in3 => \N__11667\,
            lcout => \READ_CYCLE_ACTIVE_rep17_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12835\,
            ce => \N__12647\,
            sr => \N__12498\
        );

    \GB_BUFFER_CLK40_THRU_LUT4_0_LC_23_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12848\,
            lcout => \GB_BUFFER_CLK40_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_23_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11971\,
            in1 => \N__11608\,
            in2 => \N__10447\,
            in3 => \N__11066\,
            lcout => \READ_CYCLE_ACTIVE_rep21_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12825\,
            ce => \N__12641\,
            sr => \N__12495\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_23_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__10238\,
            in1 => \N__12051\,
            in2 => \N__11131\,
            in3 => \N__11596\,
            lcout => \READ_CYCLE_ACTIVE_rep5_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12803\,
            ce => \N__12652\,
            sr => \N__12509\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__10239\,
            in1 => \N__12052\,
            in2 => \N__11132\,
            in3 => \N__11597\,
            lcout => \READ_CYCLE_ACTIVE_rep6_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12803\,
            ce => \N__12652\,
            sr => \N__12509\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_23_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__10237\,
            in1 => \N__12050\,
            in2 => \N__11130\,
            in3 => \N__11595\,
            lcout => \READ_CYCLE_ACTIVE_rep15_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12803\,
            ce => \N__12652\,
            sr => \N__12509\
        );

    \D_UU_040_iobuf_RNO_5_LC_23_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9551\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_186_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_040_iobuf_RNO_6_LC_23_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9530\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_187_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_4_LC_23_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10028\,
            lcout => \N_193_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_5_LC_23_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12266\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_194_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_0_LC_24_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9644\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_205_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_1_LC_24_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9650\,
            lcout => \N_206_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_3_LC_24_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9638\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_208_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_24_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__10442\,
            in1 => \N__12047\,
            in2 => \N__11739\,
            in3 => \N__10824\,
            lcout => \READ_CYCLE_ACTIVE_rep25_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12844\,
            ce => \N__12655\,
            sr => \N__12508\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_24_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__12046\,
            in1 => \N__11711\,
            in2 => \N__10953\,
            in3 => \N__10441\,
            lcout => \READ_CYCLE_ACTIVE_rep24_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12844\,
            ce => \N__12655\,
            sr => \N__12508\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_24_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__12048\,
            in1 => \N__11715\,
            in2 => \N__10954\,
            in3 => \N__10443\,
            lcout => \READ_CYCLE_ACTIVE_rep27_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12844\,
            ce => \N__12655\,
            sr => \N__12508\
        );

    \D_LL_040_iobuf_RNO_6_LC_24_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9824\,
            lcout => \N_211_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_2_LC_24_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9845\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_207_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_24_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__10338\,
            in1 => \N__12044\,
            in2 => \N__11554\,
            in3 => \N__10839\,
            lcout => \READ_CYCLE_ACTIVE_rep30_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12841\,
            ce => \N__12651\,
            sr => \N__12504\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_24_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__12045\,
            in1 => \N__11457\,
            in2 => \N__10965\,
            in3 => \N__10339\,
            lcout => \READ_CYCLE_ACTIVE_rep31_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12841\,
            ce => \N__12651\,
            sr => \N__12504\
        );

    \D_LM_040_iobuf_RNO_1_LC_24_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9818\,
            lcout => \N_198_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_2_LC_24_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9797\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_199_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_7_LC_24_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9779\,
            lcout => \N_212_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_0_LC_24_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9935\,
            lcout => \N_197_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_3_LC_24_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9731\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_200_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_24_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11973\,
            in1 => \N__11662\,
            in2 => \N__10966\,
            in3 => \N__10249\,
            lcout => \READ_CYCLE_ACTIVE_rep19_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12833\,
            ce => \N__12644\,
            sr => \N__12497\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_24_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__10248\,
            in1 => \N__11972\,
            in2 => \N__11706\,
            in3 => \N__10843\,
            lcout => \READ_CYCLE_ACTIVE_rep16_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12833\,
            ce => \N__12644\,
            sr => \N__12497\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_24_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__10250\,
            in1 => \N__11974\,
            in2 => \N__11707\,
            in3 => \N__10847\,
            lcout => \READ_CYCLE_ACTIVE_rep20_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12833\,
            ce => \N__12644\,
            sr => \N__12497\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_24_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11975\,
            in1 => \N__11666\,
            in2 => \N__10967\,
            in3 => \N__10251\,
            lcout => \READ_CYCLE_ACTIVE_rep8_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12833\,
            ce => \N__12644\,
            sr => \N__12497\
        );

    \D_LM_040_iobuf_RNO_4_LC_24_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9929\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_201_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_0_LC_24_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9911\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_189_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_5_LC_24_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9896\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_202_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_5_LC_24_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10022\,
            lcout => \N_210_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_2_LC_24_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9851\,
            lcout => \N_191_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_24_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11606\,
            in1 => \N__11903\,
            in2 => \N__10336\,
            in3 => \N__10851\,
            lcout => \READ_CYCLE_ACTIVE_rep10_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12826\,
            ce => \N__12640\,
            sr => \N__12496\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_24_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11607\,
            in1 => \N__11904\,
            in2 => \N__10337\,
            in3 => \N__10852\,
            lcout => \READ_CYCLE_ACTIVE_rep29_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12826\,
            ce => \N__12640\,
            sr => \N__12496\
        );

    \D_UM_040_iobuf_RNO_6_LC_24_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10004\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_195_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_24_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__10854\,
            in1 => \N__11901\,
            in2 => \N__10241\,
            in3 => \N__11489\,
            lcout => \READ_CYCLE_ACTIVE_rep22_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12824\,
            ce => \N__12642\,
            sr => \N__12499\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_24_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__11902\,
            in1 => \N__10170\,
            in2 => \N__11586\,
            in3 => \N__10855\,
            lcout => \READ_CYCLE_ACTIVE_rep23_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12824\,
            ce => \N__12642\,
            sr => \N__12499\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_24_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__10853\,
            in1 => \N__11900\,
            in2 => \N__10240\,
            in3 => \N__11488\,
            lcout => \READ_CYCLE_ACTIVE_rep14_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12824\,
            ce => \N__12642\,
            sr => \N__12499\
        );

    \D_LM_040_iobuf_RNO_6_LC_24_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9998\,
            lcout => \N_203_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_7_LC_24_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9980\,
            lcout => \N_204_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_24_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11925\,
            in1 => \N__11538\,
            in2 => \N__10232\,
            in3 => \N__10968\,
            lcout => \READ_CYCLE_ACTIVE_rep9_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12818\,
            ce => \N__12648\,
            sr => \N__12506\
        );

    \D_UM_040_iobuf_RNO_1_LC_24_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9956\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_190_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_24_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11926\,
            in1 => \N__11535\,
            in2 => \N__10233\,
            in3 => \N__10969\,
            lcout => \READ_CYCLE_ACTIVE_rep11_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12814\,
            ce => \N__12654\,
            sr => \N__12510\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_24_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11536\,
            in1 => \N__11927\,
            in2 => \N__11067\,
            in3 => \N__10148\,
            lcout => \READ_CYCLE_ACTIVE_rep1_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12814\,
            ce => \N__12654\,
            sr => \N__12510\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_24_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11928\,
            in1 => \N__11537\,
            in2 => \N__10234\,
            in3 => \N__10973\,
            lcout => \READ_CYCLE_ACTIVE_rep3_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12814\,
            ce => \N__12654\,
            sr => \N__12510\
        );

    \D_UM_040_iobuf_RNO_3_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12350\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_192_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_040_iobuf_RNO_3_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12329\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_184_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_7_LC_24_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12305\,
            lcout => \N_196_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_040_iobuf_RNO_1_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12284\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_182_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_24_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11994\,
            in1 => \N__11594\,
            in2 => \N__11069\,
            in3 => \N__10236\,
            lcout => \READ_CYCLE_ACTIVE_rep13_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12804\,
            ce => \N__12656\,
            sr => \N__12511\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_24_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11993\,
            in1 => \N__11593\,
            in2 => \N__11068\,
            in3 => \N__10235\,
            lcout => \READ_CYCLE_ACTIVE_rep12_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12804\,
            ce => \N__12656\,
            sr => \N__12511\
        );
end \INTERFACE\;
